
module router ( clk, reset, currx, curry, flitin_0, flitin_1, flitout_0, 
        flitout_1, creditin_0, creditin_1, creditout_0, creditout_1, seu );
  input [2:0] currx;
  input [2:0] curry;
  input [11:0] flitin_0;
  input [11:0] flitin_1;
  output [11:0] flitout_0;
  output [11:0] flitout_1;
  input clk, reset, creditin_0, creditin_1, seu;
  output creditout_0, creditout_1;
  wire   nomorebufs_0, debitout_0, tailout_0, nomorebufs_1, debitout_1,
         tailout_1, net1, c0nm_n2, c0nm_n1, c0nm__logic0_, c0nm_b0m_n1,
         c0nm_b0m_n9, c0nm_b0m_dqenablereg, c0nm_b0m_wdata_2_,
         c0nm_b0m_wdata_3_, c0nm_b0m_wdata_4_, c0nm_b0m_wdata_5_,
         c0nm_b0m_wdata_6_, c0nm_b0m_wdata_7_, c0nm_b0m_wdata_8_,
         c0nm_b0m_wdata_9_, c0nm_b0m_wdata_10_, c0nm_b0m_wdata_11_,
         c0nm_b0m_headflit_8_, c0nm_b0m_headflit_9_, c0nm_b0m_headflit_10_,
         c0nm_b0m_headflit_11_, c0nm_b0m__logic0_, c0nm_b0m_v0m_n276,
         c0nm_b0m_v0m_n275, c0nm_b0m_v0m_n274, c0nm_b0m_v0m_n273,
         c0nm_b0m_v0m_n272, c0nm_b0m_v0m_n271, c0nm_b0m_v0m_n270,
         c0nm_b0m_v0m_n269, c0nm_b0m_v0m_n268, c0nm_b0m_v0m_n267,
         c0nm_b0m_v0m_n266, c0nm_b0m_v0m_n265, c0nm_b0m_v0m_n264,
         c0nm_b0m_v0m_n263, c0nm_b0m_v0m_n262, c0nm_b0m_v0m_n195,
         c0nm_b0m_v0m_n194, c0nm_b0m_v0m_n193, c0nm_b0m_v0m_n192,
         c0nm_b0m_v0m_n191, c0nm_b0m_v0m_n190, c0nm_b0m_v0m_n189,
         c0nm_b0m_v0m_n188, c0nm_b0m_v0m_n187, c0nm_b0m_v0m_n186,
         c0nm_b0m_v0m_n185, c0nm_b0m_v0m_n184, c0nm_b0m_v0m_n183,
         c0nm_b0m_v0m_n182, c0nm_b0m_v0m_n181, c0nm_b0m_v0m_n180,
         c0nm_b0m_v0m_n179, c0nm_b0m_v0m_n178, c0nm_b0m_v0m_n177,
         c0nm_b0m_v0m_n176, c0nm_b0m_v0m_n175, c0nm_b0m_v0m_n174,
         c0nm_b0m_v0m_n173, c0nm_b0m_v0m_n172, c0nm_b0m_v0m_n171,
         c0nm_b0m_v0m_n170, c0nm_b0m_v0m_n169, c0nm_b0m_v0m_n168,
         c0nm_b0m_v0m_n167, c0nm_b0m_v0m_n166, c0nm_b0m_v0m_n165,
         c0nm_b0m_v0m_n164, c0nm_b0m_v0m_n163, c0nm_b0m_v0m_n162,
         c0nm_b0m_v0m_n161, c0nm_b0m_v0m_n160, c0nm_b0m_v0m_n159,
         c0nm_b0m_v0m_n158, c0nm_b0m_v0m_n157, c0nm_b0m_v0m_n156,
         c0nm_b0m_v0m_n155, c0nm_b0m_v0m_n154, c0nm_b0m_v0m_n153,
         c0nm_b0m_v0m_n152, c0nm_b0m_v0m_n151, c0nm_b0m_v0m_n150,
         c0nm_b0m_v0m_n149, c0nm_b0m_v0m_n148, c0nm_b0m_v0m_n147,
         c0nm_b0m_v0m_n146, c0nm_b0m_v0m_n145, c0nm_b0m_v0m_n144,
         c0nm_b0m_v0m_n143, c0nm_b0m_v0m_n142, c0nm_b0m_v0m_n141,
         c0nm_b0m_v0m_n140, c0nm_b0m_v0m_n139, c0nm_b0m_v0m_n138,
         c0nm_b0m_v0m_n137, c0nm_b0m_v0m_n136, c0nm_b0m_v0m_n135,
         c0nm_b0m_v0m_n134, c0nm_b0m_v0m_n133, c0nm_b0m_v0m_n132,
         c0nm_b0m_v0m_n131, c0nm_b0m_v0m_n130, c0nm_b0m_v0m_n129,
         c0nm_b0m_v0m_n128, c0nm_b0m_v0m_n127, c0nm_b0m_v0m_n126,
         c0nm_b0m_v0m_n125, c0nm_b0m_v0m_n124, c0nm_b0m_v0m_n123,
         c0nm_b0m_v0m_n122, c0nm_b0m_v0m_n121, c0nm_b0m_v0m_n120,
         c0nm_b0m_v0m_n119, c0nm_b0m_v0m_n118, c0nm_b0m_v0m_n117,
         c0nm_b0m_v0m_n116, c0nm_b0m_v0m_n115, c0nm_b0m_v0m_n114,
         c0nm_b0m_v0m_n113, c0nm_b0m_v0m_n112, c0nm_b0m_v0m_n111,
         c0nm_b0m_v0m_n110, c0nm_b0m_v0m_n109, c0nm_b0m_v0m_n108,
         c0nm_b0m_v0m_n107, c0nm_b0m_v0m_n106, c0nm_b0m_v0m_n105,
         c0nm_b0m_v0m_n104, c0nm_b0m_v0m_n103, c0nm_b0m_v0m_n102,
         c0nm_b0m_v0m_n101, c0nm_b0m_v0m_n100, c0nm_b0m_v0m_n99,
         c0nm_b0m_v0m_n98, c0nm_b0m_v0m_n97, c0nm_b0m_v0m_n96,
         c0nm_b0m_v0m_n95, c0nm_b0m_v0m_n94, c0nm_b0m_v0m_n93,
         c0nm_b0m_v0m_n92, c0nm_b0m_v0m_n91, c0nm_b0m_v0m_n90,
         c0nm_b0m_v0m_n89, c0nm_b0m_v0m_n88, c0nm_b0m_v0m_n87,
         c0nm_b0m_v0m_n86, c0nm_b0m_v0m_n85, c0nm_b0m_v0m_n84,
         c0nm_b0m_v0m_n83, c0nm_b0m_v0m_n82, c0nm_b0m_v0m_n81,
         c0nm_b0m_v0m_n80, c0nm_b0m_v0m_n79, c0nm_b0m_v0m_n78,
         c0nm_b0m_v0m_n77, c0nm_b0m_v0m_n76, c0nm_b0m_v0m_n75,
         c0nm_b0m_v0m_n74, c0nm_b0m_v0m_n73, c0nm_b0m_v0m_n72,
         c0nm_b0m_v0m_n71, c0nm_b0m_v0m_n70, c0nm_b0m_v0m_n69,
         c0nm_b0m_v0m_n68, c0nm_b0m_v0m_n67, c0nm_b0m_v0m_n66,
         c0nm_b0m_v0m_n65, c0nm_b0m_v0m_n64, c0nm_b0m_v0m_n63,
         c0nm_b0m_v0m_n62, c0nm_b0m_v0m_n49, c0nm_b0m_v0m_n48,
         c0nm_b0m_v0m_n47, c0nm_b0m_v0m_n46, c0nm_b0m_v0m_n45,
         c0nm_b0m_v0m_n44, c0nm_b0m_v0m_n43, c0nm_b0m_v0m_n42,
         c0nm_b0m_v0m_n41, c0nm_b0m_v0m_n40, c0nm_b0m_v0m_n39,
         c0nm_b0m_v0m_n38, c0nm_b0m_v0m_n37, c0nm_b0m_v0m_n36,
         c0nm_b0m_v0m_n35, c0nm_b0m_v0m_n34, c0nm_b0m_v0m_n33,
         c0nm_b0m_v0m_n32, c0nm_b0m_v0m_n31, c0nm_b0m_v0m_n30,
         c0nm_b0m_v0m_n29, c0nm_b0m_v0m_n28, c0nm_b0m_v0m_n27,
         c0nm_b0m_v0m_n26, c0nm_b0m_v0m_n25, c0nm_b0m_v0m_n24,
         c0nm_b0m_v0m_n23, c0nm_b0m_v0m_n22, c0nm_b0m_v0m_n21,
         c0nm_b0m_v0m_n20, c0nm_b0m_v0m_n19, c0nm_b0m_v0m_n18,
         c0nm_b0m_v0m_n17, c0nm_b0m_v0m_n16, c0nm_b0m_v0m_n15,
         c0nm_b0m_v0m_n14, c0nm_b0m_v0m_n13, c0nm_b0m_v0m_n12,
         c0nm_b0m_v0m_n11, c0nm_b0m_v0m_n10, c0nm_b0m_v0m_n8, c0nm_b0m_v0m_n7,
         c0nm_b0m_v0m_n6, c0nm_b0m_v0m_n5, c0nm_b0m_v0m_n4, c0nm_b0m_v0m_n3,
         c0nm_b0m_v0m_n2, c0nm_b0m_v0m_n1, c0nm_b0m_v0m_n261,
         c0nm_b0m_v0m_n260, c0nm_b0m_v0m_n259, c0nm_b0m_v0m_n258,
         c0nm_b0m_v0m_n257, c0nm_b0m_v0m_n256, c0nm_b0m_v0m_n255,
         c0nm_b0m_v0m_n254, c0nm_b0m_v0m_n253, c0nm_b0m_v0m_n252,
         c0nm_b0m_v0m_n251, c0nm_b0m_v0m_n250, c0nm_b0m_v0m_n249,
         c0nm_b0m_v0m_n248, c0nm_b0m_v0m_n247, c0nm_b0m_v0m_n246,
         c0nm_b0m_v0m_n245, c0nm_b0m_v0m_n244, c0nm_b0m_v0m_n243,
         c0nm_b0m_v0m_n242, c0nm_b0m_v0m_n241, c0nm_b0m_v0m_n240,
         c0nm_b0m_v0m_n239, c0nm_b0m_v0m_n238, c0nm_b0m_v0m_n237,
         c0nm_b0m_v0m_n236, c0nm_b0m_v0m_n235, c0nm_b0m_v0m_n234,
         c0nm_b0m_v0m_n233, c0nm_b0m_v0m_n232, c0nm_b0m_v0m_n231,
         c0nm_b0m_v0m_n230, c0nm_b0m_v0m_n229, c0nm_b0m_v0m_n228,
         c0nm_b0m_v0m_n227, c0nm_b0m_v0m_n226, c0nm_b0m_v0m_n225,
         c0nm_b0m_v0m_n224, c0nm_b0m_v0m_n223, c0nm_b0m_v0m_n222,
         c0nm_b0m_v0m_n221, c0nm_b0m_v0m_n220, c0nm_b0m_v0m_n219,
         c0nm_b0m_v0m_n218, c0nm_b0m_v0m_n217, c0nm_b0m_v0m_n216,
         c0nm_b0m_v0m_n215, c0nm_b0m_v0m_n214, c0nm_b0m_v0m_n213,
         c0nm_b0m_v0m_n212, c0nm_b0m_v0m_n211, c0nm_b0m_v0m_n210,
         c0nm_b0m_v0m_n209, c0nm_b0m_v0m_n208, c0nm_b0m_v0m_n207,
         c0nm_b0m_v0m_n206, c0nm_b0m_v0m_n205, c0nm_b0m_v0m_n204,
         c0nm_b0m_v0m_n203, c0nm_b0m_v0m_n202, c0nm_b0m_v0m_n201,
         c0nm_b0m_v0m_n200, c0nm_b0m_v0m_n199, c0nm_b0m_v0m_n198,
         c0nm_b0m_v0m_n197, c0nm_b0m_v0m_n196, c0nm_b0m_v0m_n61,
         c0nm_b0m_v0m_n60, c0nm_b0m_v0m_n59, c0nm_b0m_v0m_n58,
         c0nm_b0m_v0m_n57, c0nm_b0m_v0m_n56, c0nm_b0m_v0m_n55,
         c0nm_b0m_v0m_n54, c0nm_b0m_v0m_n53, c0nm_b0m_v0m_n52,
         c0nm_b0m_v0m_n51, c0nm_b0m_v0m_n50, c0nm_b0m_v0m_n9,
         c0nm_b0m_v0m_n1710, c0nm_b0m_v0m_tail_0_, c0nm_b0m_v0m_tail_1_,
         c0nm_b0m_v0m_buffers3_0_, c0nm_b0m_v0m_buffers3_1_,
         c0nm_b0m_v0m_buffers3_2_, c0nm_b0m_v0m_buffers3_3_,
         c0nm_b0m_v0m_buffers3_4_, c0nm_b0m_v0m_buffers3_5_,
         c0nm_b0m_v0m_buffers3_6_, c0nm_b0m_v0m_buffers3_7_,
         c0nm_b0m_v0m_buffers3_8_, c0nm_b0m_v0m_buffers3_9_,
         c0nm_b0m_v0m_buffers3_10_, c0nm_b0m_v0m_buffers3_11_,
         c0nm_b0m_v0m_buffers2_0_, c0nm_b0m_v0m_buffers2_1_,
         c0nm_b0m_v0m_buffers2_2_, c0nm_b0m_v0m_buffers2_3_,
         c0nm_b0m_v0m_buffers2_4_, c0nm_b0m_v0m_buffers2_5_,
         c0nm_b0m_v0m_buffers2_6_, c0nm_b0m_v0m_buffers2_7_,
         c0nm_b0m_v0m_buffers2_8_, c0nm_b0m_v0m_buffers2_9_,
         c0nm_b0m_v0m_buffers2_10_, c0nm_b0m_v0m_buffers2_11_,
         c0nm_b0m_v0m_buffers0_0_, c0nm_b0m_v0m_buffers0_1_,
         c0nm_b0m_v0m_buffers0_2_, c0nm_b0m_v0m_buffers0_3_,
         c0nm_b0m_v0m_buffers0_4_, c0nm_b0m_v0m_buffers0_5_,
         c0nm_b0m_v0m_buffers0_6_, c0nm_b0m_v0m_buffers0_7_,
         c0nm_b0m_v0m_buffers0_8_, c0nm_b0m_v0m_buffers0_9_,
         c0nm_b0m_v0m_buffers0_10_, c0nm_b0m_v0m_buffers0_11_,
         c0nm_b0m_v0m_head_0_, c0nm_b0m_v0m_head_1_, c0nm_b0m_v0m_head_2_,
         c0nm_r0m_n16, c0nm_r0m_n15, c0nm_r0m_n14, c0nm_r0m_n13, c0nm_r0m_n12,
         c0nm_r0m_n11, c0nm_r0m_n10, c0nm_r0m_n9, c0nm_r0m_n8, c0nm_r0m_n7,
         c0nm_r0m_n6, c0nm_r0m_n5, c0nm_r0m_n4, c0nm_r0m_n3, c0nm_r0m_n2,
         c0nm_r0m_n1, c0nm_r0m_n110, c0nm_r0m_n100, c0nm_v0m_n29, c0nm_v0m_n28,
         c0nm_v0m_n27, c0nm_v0m_n26, c0nm_v0m_n25, c0nm_v0m_n24, c0nm_v0m_n23,
         c0nm_v0m_n22, c0nm_v0m_n21, c0nm_v0m_n20, c0nm_v0m_n19, c0nm_v0m_n18,
         c0nm_v0m_n17, c0nm_v0m_n16, c0nm_v0m_n15, c0nm_v0m_n14, c0nm_v0m_n13,
         c0nm_v0m_n12, c0nm_v0m_n11, c0nm_v0m_n10, c0nm_v0m_n9, c0nm_v0m_n8,
         c0nm_v0m_n7, c0nm_v0m_n6, c0nm_v0m_n5, c0nm_v0m_n4, c0nm_v0m_n3,
         c0nm_v0m_n2, c0nm_v0m_n1, c0nm_v0m_n31, c0nm_v0m_n30, c0nm_v0m_n64,
         c0nm_v0m_n63, c0nm_v0m_n62, c0nm_v0m_n61, c0nm_v0m_n58, c0nm_v0m_n57,
         c0nm_v0m_full, c0nm_v0m_state_queuelen_0_, c0nm_v0m_state_queuelen_1_,
         c0nm_v0m_state_queuelen_2_, c0nm_v0m_state_status_0_,
         c0nm_v0m_state_status_1_, c0sm_n4, c0sm_n3, c0sm__logic0_,
         c0sm_b0m_n2, c0sm_b0m_n9, c0sm_b0m_dqenablereg, c0sm_b0m_wdata_2_,
         c0sm_b0m_wdata_3_, c0sm_b0m_wdata_4_, c0sm_b0m_wdata_5_,
         c0sm_b0m_wdata_6_, c0sm_b0m_wdata_7_, c0sm_b0m_wdata_8_,
         c0sm_b0m_wdata_9_, c0sm_b0m_wdata_10_, c0sm_b0m_wdata_11_,
         c0sm_b0m_headflit_8_, c0sm_b0m_headflit_9_, c0sm_b0m_headflit_10_,
         c0sm_b0m_headflit_11_, c0sm_b0m__logic0_, c0sm_b0m_v0m_n355,
         c0sm_b0m_v0m_n354, c0sm_b0m_v0m_n353, c0sm_b0m_v0m_n352,
         c0sm_b0m_v0m_n351, c0sm_b0m_v0m_n350, c0sm_b0m_v0m_n349,
         c0sm_b0m_v0m_n348, c0sm_b0m_v0m_n347, c0sm_b0m_v0m_n346,
         c0sm_b0m_v0m_n345, c0sm_b0m_v0m_n344, c0sm_b0m_v0m_n343,
         c0sm_b0m_v0m_n342, c0sm_b0m_v0m_n341, c0sm_b0m_v0m_n340,
         c0sm_b0m_v0m_n339, c0sm_b0m_v0m_n338, c0sm_b0m_v0m_n337,
         c0sm_b0m_v0m_n336, c0sm_b0m_v0m_n335, c0sm_b0m_v0m_n334,
         c0sm_b0m_v0m_n333, c0sm_b0m_v0m_n332, c0sm_b0m_v0m_n331,
         c0sm_b0m_v0m_n330, c0sm_b0m_v0m_n329, c0sm_b0m_v0m_n328,
         c0sm_b0m_v0m_n327, c0sm_b0m_v0m_n326, c0sm_b0m_v0m_n325,
         c0sm_b0m_v0m_n324, c0sm_b0m_v0m_n323, c0sm_b0m_v0m_n322,
         c0sm_b0m_v0m_n321, c0sm_b0m_v0m_n320, c0sm_b0m_v0m_n319,
         c0sm_b0m_v0m_n318, c0sm_b0m_v0m_n317, c0sm_b0m_v0m_n316,
         c0sm_b0m_v0m_n315, c0sm_b0m_v0m_n314, c0sm_b0m_v0m_n313,
         c0sm_b0m_v0m_n312, c0sm_b0m_v0m_n311, c0sm_b0m_v0m_n310,
         c0sm_b0m_v0m_n309, c0sm_b0m_v0m_n308, c0sm_b0m_v0m_n307,
         c0sm_b0m_v0m_n306, c0sm_b0m_v0m_n305, c0sm_b0m_v0m_n304,
         c0sm_b0m_v0m_n303, c0sm_b0m_v0m_n302, c0sm_b0m_v0m_n301,
         c0sm_b0m_v0m_n300, c0sm_b0m_v0m_n299, c0sm_b0m_v0m_n298,
         c0sm_b0m_v0m_n297, c0sm_b0m_v0m_n296, c0sm_b0m_v0m_n295,
         c0sm_b0m_v0m_n294, c0sm_b0m_v0m_n293, c0sm_b0m_v0m_n292,
         c0sm_b0m_v0m_n291, c0sm_b0m_v0m_n290, c0sm_b0m_v0m_n289,
         c0sm_b0m_v0m_n288, c0sm_b0m_v0m_n287, c0sm_b0m_v0m_n286,
         c0sm_b0m_v0m_n285, c0sm_b0m_v0m_n284, c0sm_b0m_v0m_n283,
         c0sm_b0m_v0m_n282, c0sm_b0m_v0m_n281, c0sm_b0m_v0m_n280,
         c0sm_b0m_v0m_n279, c0sm_b0m_v0m_n278, c0sm_b0m_v0m_n277,
         c0sm_b0m_v0m_n276, c0sm_b0m_v0m_n275, c0sm_b0m_v0m_n274,
         c0sm_b0m_v0m_n273, c0sm_b0m_v0m_n272, c0sm_b0m_v0m_n271,
         c0sm_b0m_v0m_n270, c0sm_b0m_v0m_n269, c0sm_b0m_v0m_n268,
         c0sm_b0m_v0m_n267, c0sm_b0m_v0m_n266, c0sm_b0m_v0m_n265,
         c0sm_b0m_v0m_n264, c0sm_b0m_v0m_n263, c0sm_b0m_v0m_n262,
         c0sm_b0m_v0m_n195, c0sm_b0m_v0m_n194, c0sm_b0m_v0m_n193,
         c0sm_b0m_v0m_n192, c0sm_b0m_v0m_n191, c0sm_b0m_v0m_n190,
         c0sm_b0m_v0m_n189, c0sm_b0m_v0m_n188, c0sm_b0m_v0m_n187,
         c0sm_b0m_v0m_n186, c0sm_b0m_v0m_n185, c0sm_b0m_v0m_n184,
         c0sm_b0m_v0m_n183, c0sm_b0m_v0m_n182, c0sm_b0m_v0m_n181,
         c0sm_b0m_v0m_n180, c0sm_b0m_v0m_n179, c0sm_b0m_v0m_n178,
         c0sm_b0m_v0m_n177, c0sm_b0m_v0m_n176, c0sm_b0m_v0m_n175,
         c0sm_b0m_v0m_n174, c0sm_b0m_v0m_n173, c0sm_b0m_v0m_n172,
         c0sm_b0m_v0m_n171, c0sm_b0m_v0m_n170, c0sm_b0m_v0m_n169,
         c0sm_b0m_v0m_n168, c0sm_b0m_v0m_n167, c0sm_b0m_v0m_n166,
         c0sm_b0m_v0m_n165, c0sm_b0m_v0m_n164, c0sm_b0m_v0m_n163,
         c0sm_b0m_v0m_n162, c0sm_b0m_v0m_n161, c0sm_b0m_v0m_n160,
         c0sm_b0m_v0m_n159, c0sm_b0m_v0m_n158, c0sm_b0m_v0m_n157,
         c0sm_b0m_v0m_n156, c0sm_b0m_v0m_n155, c0sm_b0m_v0m_n154,
         c0sm_b0m_v0m_n153, c0sm_b0m_v0m_n152, c0sm_b0m_v0m_n151,
         c0sm_b0m_v0m_n150, c0sm_b0m_v0m_n149, c0sm_b0m_v0m_n148,
         c0sm_b0m_v0m_n147, c0sm_b0m_v0m_n146, c0sm_b0m_v0m_n145,
         c0sm_b0m_v0m_n144, c0sm_b0m_v0m_n143, c0sm_b0m_v0m_n142,
         c0sm_b0m_v0m_n141, c0sm_b0m_v0m_n140, c0sm_b0m_v0m_n139,
         c0sm_b0m_v0m_n138, c0sm_b0m_v0m_n137, c0sm_b0m_v0m_n136,
         c0sm_b0m_v0m_n135, c0sm_b0m_v0m_n134, c0sm_b0m_v0m_n133,
         c0sm_b0m_v0m_n132, c0sm_b0m_v0m_n131, c0sm_b0m_v0m_n130,
         c0sm_b0m_v0m_n129, c0sm_b0m_v0m_n128, c0sm_b0m_v0m_n127,
         c0sm_b0m_v0m_n126, c0sm_b0m_v0m_n125, c0sm_b0m_v0m_n124,
         c0sm_b0m_v0m_n123, c0sm_b0m_v0m_n122, c0sm_b0m_v0m_n121,
         c0sm_b0m_v0m_n120, c0sm_b0m_v0m_n119, c0sm_b0m_v0m_n118,
         c0sm_b0m_v0m_n117, c0sm_b0m_v0m_n116, c0sm_b0m_v0m_n115,
         c0sm_b0m_v0m_n114, c0sm_b0m_v0m_n113, c0sm_b0m_v0m_n112,
         c0sm_b0m_v0m_n111, c0sm_b0m_v0m_n110, c0sm_b0m_v0m_n109,
         c0sm_b0m_v0m_n108, c0sm_b0m_v0m_n107, c0sm_b0m_v0m_n106,
         c0sm_b0m_v0m_n105, c0sm_b0m_v0m_n104, c0sm_b0m_v0m_n103,
         c0sm_b0m_v0m_n102, c0sm_b0m_v0m_n101, c0sm_b0m_v0m_n100,
         c0sm_b0m_v0m_n99, c0sm_b0m_v0m_n98, c0sm_b0m_v0m_n97,
         c0sm_b0m_v0m_n96, c0sm_b0m_v0m_n95, c0sm_b0m_v0m_n94,
         c0sm_b0m_v0m_n93, c0sm_b0m_v0m_n92, c0sm_b0m_v0m_n91,
         c0sm_b0m_v0m_n90, c0sm_b0m_v0m_n89, c0sm_b0m_v0m_n88,
         c0sm_b0m_v0m_n87, c0sm_b0m_v0m_n86, c0sm_b0m_v0m_n85,
         c0sm_b0m_v0m_n84, c0sm_b0m_v0m_n83, c0sm_b0m_v0m_n82,
         c0sm_b0m_v0m_n81, c0sm_b0m_v0m_n80, c0sm_b0m_v0m_n79,
         c0sm_b0m_v0m_n78, c0sm_b0m_v0m_n77, c0sm_b0m_v0m_n76,
         c0sm_b0m_v0m_n75, c0sm_b0m_v0m_n74, c0sm_b0m_v0m_n73,
         c0sm_b0m_v0m_n72, c0sm_b0m_v0m_n71, c0sm_b0m_v0m_n70,
         c0sm_b0m_v0m_n69, c0sm_b0m_v0m_n68, c0sm_b0m_v0m_n67,
         c0sm_b0m_v0m_n66, c0sm_b0m_v0m_n65, c0sm_b0m_v0m_n64,
         c0sm_b0m_v0m_n63, c0sm_b0m_v0m_n62, c0sm_b0m_v0m_n49,
         c0sm_b0m_v0m_n48, c0sm_b0m_v0m_n47, c0sm_b0m_v0m_n46,
         c0sm_b0m_v0m_n45, c0sm_b0m_v0m_n44, c0sm_b0m_v0m_n43,
         c0sm_b0m_v0m_n42, c0sm_b0m_v0m_n41, c0sm_b0m_v0m_n40,
         c0sm_b0m_v0m_n39, c0sm_b0m_v0m_n38, c0sm_b0m_v0m_n37,
         c0sm_b0m_v0m_n36, c0sm_b0m_v0m_n35, c0sm_b0m_v0m_n34,
         c0sm_b0m_v0m_n33, c0sm_b0m_v0m_n32, c0sm_b0m_v0m_n31,
         c0sm_b0m_v0m_n30, c0sm_b0m_v0m_n29, c0sm_b0m_v0m_n28,
         c0sm_b0m_v0m_n27, c0sm_b0m_v0m_n26, c0sm_b0m_v0m_n25,
         c0sm_b0m_v0m_n24, c0sm_b0m_v0m_n23, c0sm_b0m_v0m_n22,
         c0sm_b0m_v0m_n21, c0sm_b0m_v0m_n20, c0sm_b0m_v0m_n19,
         c0sm_b0m_v0m_n18, c0sm_b0m_v0m_n17, c0sm_b0m_v0m_n16,
         c0sm_b0m_v0m_n15, c0sm_b0m_v0m_n14, c0sm_b0m_v0m_n13,
         c0sm_b0m_v0m_n12, c0sm_b0m_v0m_n11, c0sm_b0m_v0m_n10, c0sm_b0m_v0m_n8,
         c0sm_b0m_v0m_n7, c0sm_b0m_v0m_n6, c0sm_b0m_v0m_n5, c0sm_b0m_v0m_n4,
         c0sm_b0m_v0m_n3, c0sm_b0m_v0m_n2, c0sm_b0m_v0m_n1, c0sm_b0m_v0m_n1710,
         c0sm_b0m_v0m_tail_0_, c0sm_b0m_v0m_tail_1_, c0sm_b0m_v0m_buffers3_0_,
         c0sm_b0m_v0m_buffers3_1_, c0sm_b0m_v0m_buffers3_2_,
         c0sm_b0m_v0m_buffers3_3_, c0sm_b0m_v0m_buffers3_4_,
         c0sm_b0m_v0m_buffers3_5_, c0sm_b0m_v0m_buffers3_6_,
         c0sm_b0m_v0m_buffers3_7_, c0sm_b0m_v0m_buffers3_8_,
         c0sm_b0m_v0m_buffers3_9_, c0sm_b0m_v0m_buffers3_10_,
         c0sm_b0m_v0m_buffers3_11_, c0sm_b0m_v0m_buffers2_0_,
         c0sm_b0m_v0m_buffers2_1_, c0sm_b0m_v0m_buffers2_2_,
         c0sm_b0m_v0m_buffers2_3_, c0sm_b0m_v0m_buffers2_4_,
         c0sm_b0m_v0m_buffers2_5_, c0sm_b0m_v0m_buffers2_6_,
         c0sm_b0m_v0m_buffers2_7_, c0sm_b0m_v0m_buffers2_8_,
         c0sm_b0m_v0m_buffers2_9_, c0sm_b0m_v0m_buffers2_10_,
         c0sm_b0m_v0m_buffers2_11_, c0sm_b0m_v0m_buffers0_0_,
         c0sm_b0m_v0m_buffers0_1_, c0sm_b0m_v0m_buffers0_2_,
         c0sm_b0m_v0m_buffers0_3_, c0sm_b0m_v0m_buffers0_4_,
         c0sm_b0m_v0m_buffers0_5_, c0sm_b0m_v0m_buffers0_6_,
         c0sm_b0m_v0m_buffers0_7_, c0sm_b0m_v0m_buffers0_8_,
         c0sm_b0m_v0m_buffers0_9_, c0sm_b0m_v0m_buffers0_10_,
         c0sm_b0m_v0m_buffers0_11_, c0sm_b0m_v0m_head_0_, c0sm_b0m_v0m_head_1_,
         c0sm_b0m_v0m_head_2_, c0sm_r0m_n16, c0sm_r0m_n15, c0sm_r0m_n14,
         c0sm_r0m_n13, c0sm_r0m_n12, c0sm_r0m_n11, c0sm_r0m_n10, c0sm_r0m_n9,
         c0sm_r0m_n8, c0sm_r0m_n7, c0sm_r0m_n6, c0sm_r0m_n5, c0sm_r0m_n4,
         c0sm_r0m_n3, c0sm_r0m_n2, c0sm_r0m_n1, c0sm_r0m_n110, c0sm_r0m_n100,
         c0sm_v0m_n33, c0sm_v0m_n32, c0sm_v0m_n29, c0sm_v0m_n28, c0sm_v0m_n27,
         c0sm_v0m_n26, c0sm_v0m_n25, c0sm_v0m_n24, c0sm_v0m_n23, c0sm_v0m_n22,
         c0sm_v0m_n21, c0sm_v0m_n20, c0sm_v0m_n19, c0sm_v0m_n18, c0sm_v0m_n17,
         c0sm_v0m_n16, c0sm_v0m_n15, c0sm_v0m_n14, c0sm_v0m_n13, c0sm_v0m_n12,
         c0sm_v0m_n11, c0sm_v0m_n10, c0sm_v0m_n9, c0sm_v0m_n8, c0sm_v0m_n7,
         c0sm_v0m_n6, c0sm_v0m_n5, c0sm_v0m_n4, c0sm_v0m_n3, c0sm_v0m_n2,
         c0sm_v0m_n1, c0sm_v0m_n64, c0sm_v0m_n63, c0sm_v0m_n62, c0sm_v0m_n61,
         c0sm_v0m_n58, c0sm_v0m_n57, c0sm_v0m_full, c0sm_v0m_state_queuelen_0_,
         c0sm_v0m_state_queuelen_1_, c0sm_v0m_state_queuelen_2_,
         c0sm_v0m_state_status_0_, c0sm_v0m_state_status_1_, s0m_n26, s0m_n21,
         s0m_n20, s0m_n19, s0m_n18, s0m_n17, s0m_n16, s0m_n15, s0m_n14,
         s0m_n13, s0m_n12, s0m_n11, s0m_n10, s0m_n9, s0m_n8, s0m_n7, s0m_n6,
         s0m_n5, s0m_n4, s0m_n3, s0m_n2, s0m_n1, s0m_n25, s0m_n24, s0m_n23,
         s0m_n22, s0m_no_bufs0, s0m_no_bufs1, s0m_tail_outvc1, s0m_tail_outvc0,
         s0m_debit_outvc1, s0m_state_invc1_0_, s0m_state_invc1_1_,
         s0m_debit_outvc0, s0m_state_invc0_0_, s0m_state_invc0_1_, s0m_elig_0_,
         s0m_elig_1_, s0m_outb1_0_, s0m_outb1_1_, s0m_outb0_0_, s0m_outb0_1_,
         s0m__logic0_, s0m_m0m_n3, s0m_m0m_n2, s0m_m0m_n1, s0m_m0m_n10,
         s0m_m0m_row1_0_, s0m_m1m_n3, s0m_m1m_n2, s0m_m1m_n1, s0m_m1m_n10,
         s0m_m1m_row1_0_, s0m_o0nm_n25, s0m_o0nm_n24, s0m_o0nm_n23,
         s0m_o0nm_n22, s0m_o0nm_n21, s0m_o0nm_n20, s0m_o0nm_n19, s0m_o0nm_n18,
         s0m_o0nm_n17, s0m_o0nm_n16, s0m_o0nm_n15, s0m_o0nm_n14, s0m_o0nm_n13,
         s0m_o0nm_n12, s0m_o0nm_n11, s0m_o0nm_n10, s0m_o0nm_n9, s0m_o0nm_n8,
         s0m_o0nm_n7, s0m_o0nm_n6, s0m_o0nm_n5, s0m_o0nm_n4, s0m_o0nm_n3,
         s0m_o0nm_n2, s0m_o0nm_n1, s0m_o0nm_n31, s0m_o0nm_n30, s0m_o0nm_n42,
         s0m_o0nm_n41, s0m_o0nm_n38, s0m_o0nm_n37, s0m_o0nm_n36, s0m_o0nm_n35,
         s0m_o0nm_state_assigned, s0m_o0nm_state_credits_0_,
         s0m_o0nm_state_credits_1_, s0m_o0nm_state_credits_2_, s0m_o0sm_n27,
         s0m_o0sm_n26, s0m_o0sm_n25, s0m_o0sm_n24, s0m_o0sm_n23, s0m_o0sm_n22,
         s0m_o0sm_n21, s0m_o0sm_n20, s0m_o0sm_n19, s0m_o0sm_n18, s0m_o0sm_n17,
         s0m_o0sm_n16, s0m_o0sm_n15, s0m_o0sm_n14, s0m_o0sm_n13, s0m_o0sm_n12,
         s0m_o0sm_n11, s0m_o0sm_n10, s0m_o0sm_n9, s0m_o0sm_n8, s0m_o0sm_n7,
         s0m_o0sm_n6, s0m_o0sm_n5, s0m_o0sm_n4, s0m_o0sm_n3, s0m_o0sm_n2,
         s0m_o0sm_n1, s0m_o0sm_n42, s0m_o0sm_n41, s0m_o0sm_n38, s0m_o0sm_n37,
         s0m_o0sm_n36, s0m_o0sm_n35, s0m_o0sm_state_assigned,
         s0m_o0sm_state_credits_0_, s0m_o0sm_state_credits_1_,
         s0m_o0sm_state_credits_2_, x0m_n6, x0m_n5, x0m_n4, x0m_n3,
         x0m_colsel1reg_0_, x0m_colsel1reg_1_, x0m_colsel0reg_0_,
         x0m_colsel0reg_1_, x0m__logic0_, x0m__logic1_, x0m_bx0m_m0m_int01,
         x0m_bx0m_m1m_int01, x0m_bx1m_m0m_int01, x0m_bx1m_m1m_int01,
         x0m_bx2m_m0m_int01, x0m_bx2m_m1m_int01, x0m_bx3m_m0m_int01,
         x0m_bx3m_m1m_int01, x0m_bx4m_m0m_int01, x0m_bx4m_m1m_int01,
         x0m_bx5m_m0m_int01, x0m_bx5m_m1m_int01, x0m_bx6m_m0m_int01,
         x0m_bx6m_m1m_int01, x0m_bx7m_m0m_int01, x0m_bx7m_m1m_int01,
         x0m_bx8m_m0m_int01, x0m_bx8m_m1m_int01, x0m_bx9m_m0m_int01,
         x0m_bx9m_m1m_int01, x0m_bx10m_m0m_int01, x0m_bx10m_m1m_int01,
         x0m_bx11m_m0m_int01, x0m_bx11m_m1m_int01;
  wire   [1:0] swalloc_req_0;
  wire   [1:0] swalloc_resp_0;
  wire   [11:0] flitout_switch_0;
  wire   [1:0] swalloc_req_1;
  wire   [1:0] swalloc_resp_1;
  wire   [11:0] flitout_switch_1;
  wire   [1:0] colsel0;
  wire   [1:0] colsel1;
  wire   [1:0] c0nm_routewire;
  wire   [7:0] c0nm_headflit;
  wire   [11:0] c0nm_b0m_rdata;
  wire   [1:0] c0sm_routewire;
  wire   [7:0] c0sm_headflit;
  wire   [11:0] c0sm_b0m_rdata;
  wire   [1:0] s0m_request0;
  wire   [1:0] s0m_request1;

  TIELO_X1M_A12TR u1 ( .Y(net1) );
  NOR2B_X0P5M_A12TR c0nm_u5 ( .AN(debitout_0), .B(reset), .Y(creditout_0) );
  NOR2B_X0P5M_A12TR c0nm_u4 ( .AN(c0nm_headflit[1]), .B(c0nm_headflit[0]), .Y(
        c0nm_n1) );
  NAND2_X0P5A_A12TR c0nm_u3 ( .A(flitin_0[1]), .B(flitin_0[0]), .Y(c0nm_n2) );
  TIELO_X1M_A12TR c0nm_u2 ( .Y(c0nm__logic0_) );
  NOR2B_X0P5M_A12TR c0nm_b0m_u27 ( .AN(debitout_0), .B(reset), .Y(c0nm_b0m_n9)
         );
  NAND2B_X0P5M_A12TR c0nm_b0m_u26 ( .AN(c0nm_b0m_rdata[0]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[0]) );
  AND2_X0P5M_A12TR c0nm_b0m_u25 ( .A(c0nm_b0m_rdata[10]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[10]) );
  AND2_X0P5M_A12TR c0nm_b0m_u24 ( .A(c0nm_b0m_rdata[11]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[11]) );
  NAND2B_X0P5M_A12TR c0nm_b0m_u23 ( .AN(c0nm_b0m_rdata[1]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[1]) );
  AND2_X0P5M_A12TR c0nm_b0m_u22 ( .A(c0nm_b0m_rdata[2]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[2]) );
  AND2_X0P5M_A12TR c0nm_b0m_u21 ( .A(c0nm_b0m_rdata[3]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[3]) );
  AND2_X0P5M_A12TR c0nm_b0m_u20 ( .A(c0nm_b0m_rdata[4]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[4]) );
  AND2_X0P5M_A12TR c0nm_b0m_u19 ( .A(c0nm_b0m_rdata[5]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[5]) );
  AND2_X0P5M_A12TR c0nm_b0m_u18 ( .A(c0nm_b0m_rdata[6]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[6]) );
  AND2_X0P5M_A12TR c0nm_b0m_u17 ( .A(c0nm_b0m_rdata[7]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[7]) );
  AND2_X0P5M_A12TR c0nm_b0m_u16 ( .A(c0nm_b0m_rdata[8]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[8]) );
  AND2_X0P5M_A12TR c0nm_b0m_u15 ( .A(c0nm_b0m_rdata[9]), .B(
        c0nm_b0m_dqenablereg), .Y(flitout_switch_0[9]) );
  NAND2_X0P5A_A12TR c0nm_b0m_u14 ( .A(flitin_0[1]), .B(flitin_0[0]), .Y(
        c0nm_b0m_n1) );
  AND2_X0P5M_A12TR c0nm_b0m_u13 ( .A(flitin_0[10]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_10_) );
  AND2_X0P5M_A12TR c0nm_b0m_u12 ( .A(flitin_0[11]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_11_) );
  AND2_X0P5M_A12TR c0nm_b0m_u11 ( .A(flitin_0[2]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_2_) );
  AND2_X0P5M_A12TR c0nm_b0m_u10 ( .A(flitin_0[3]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_3_) );
  AND2_X0P5M_A12TR c0nm_b0m_u9 ( .A(flitin_0[4]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_4_) );
  AND2_X0P5M_A12TR c0nm_b0m_u8 ( .A(flitin_0[5]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_5_) );
  AND2_X0P5M_A12TR c0nm_b0m_u7 ( .A(flitin_0[6]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_6_) );
  AND2_X0P5M_A12TR c0nm_b0m_u6 ( .A(flitin_0[7]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_7_) );
  AND2_X0P5M_A12TR c0nm_b0m_u5 ( .A(flitin_0[8]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_8_) );
  AND2_X0P5M_A12TR c0nm_b0m_u4 ( .A(flitin_0[9]), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_wdata_9_) );
  TIELO_X1M_A12TR c0nm_b0m_u3 ( .Y(c0nm_b0m__logic0_) );
  DFFQ_X1M_A12TR c0nm_b0m_dqenablereg_reg ( .D(c0nm_b0m_n9), .CK(clk), .Q(
        c0nm_b0m_dqenablereg) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u278 ( .A(c0nm_b0m_v0m_head_0_), .Y(
        c0nm_b0m_v0m_n16) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u277 ( .A(c0nm_b0m_v0m_head_2_), .Y(
        c0nm_b0m_v0m_n15) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u276 ( .A(c0nm_b0m_v0m_n16), .B(
        c0nm_b0m_v0m_n15), .C(c0nm_b0m_v0m_head_1_), .Y(c0nm_b0m_v0m_n187) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u275 ( .A(c0nm_b0m_v0m_buffers2_0_), .Y(
        c0nm_b0m_v0m_n105) );
  AOI21_X0P5M_A12TR c0nm_b0m_v0m_u274 ( .A0(c0nm_b0m_v0m_head_0_), .A1(
        c0nm_b0m_v0m_head_1_), .B0(c0nm_b0m_v0m_head_2_), .Y(c0nm_b0m_v0m_n73)
         );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u273 ( .A(c0nm_b0m_v0m_buffers3_0_), .Y(
        c0nm_b0m_v0m_n23) );
  NOR3_X0P5A_A12TR c0nm_b0m_v0m_u272 ( .A(c0nm_b0m_v0m_head_1_), .B(
        c0nm_b0m_v0m_head_2_), .C(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n193)
         );
  NOR3_X0P5A_A12TR c0nm_b0m_v0m_u271 ( .A(c0nm_b0m_v0m_head_1_), .B(
        c0nm_b0m_v0m_head_2_), .C(c0nm_b0m_v0m_n16), .Y(c0nm_b0m_v0m_n192) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u270 ( .A(c0nm_b0m_v0m_n61), .Y(
        c0nm_b0m_v0m_n114) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u269 ( .A0(c0nm_b0m_v0m_buffers0_0_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n114), 
        .Y(c0nm_b0m_v0m_n276) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u268 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n105), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n23), .C0(
        c0nm_b0m_v0m_n276), .Y(c0nm_headflit[0]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u267 ( .A(c0nm_b0m_v0m_buffers2_1_), .Y(
        c0nm_b0m_v0m_n122) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u266 ( .A(c0nm_b0m_v0m_buffers3_1_), .Y(
        c0nm_b0m_v0m_n29) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u265 ( .A(c0nm_b0m_v0m_n60), .Y(
        c0nm_b0m_v0m_n125) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u264 ( .A0(c0nm_b0m_v0m_buffers0_1_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n125), 
        .Y(c0nm_b0m_v0m_n275) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u263 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n122), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n29), .C0(
        c0nm_b0m_v0m_n275), .Y(c0nm_headflit[1]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u262 ( .A(c0nm_headflit[1]), .Y(
        c0nm_b0m_v0m_n264) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u261 ( .A(reset), .Y(c0nm_b0m_v0m_n4) );
  AND4_X0P5M_A12TR c0nm_b0m_v0m_u260 ( .A(debitout_0), .B(c0nm_headflit[0]), 
        .C(c0nm_b0m_v0m_n264), .D(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n1710) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u259 ( .A(c0nm_b0m_v0m_buffers2_10_), .Y(
        c0nm_b0m_v0m_n180) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u258 ( .A(c0nm_b0m_v0m_buffers3_10_), .Y(
        c0nm_b0m_v0m_n71) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u257 ( .A(c0nm_b0m_v0m_n51), .Y(
        c0nm_b0m_v0m_n183) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u256 ( .A0(c0nm_b0m_v0m_buffers0_10_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n183), 
        .Y(c0nm_b0m_v0m_n274) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u255 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n180), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n71), .C0(
        c0nm_b0m_v0m_n274), .Y(c0nm_b0m_headflit_10_) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u254 ( .A(c0nm_b0m_v0m_buffers2_11_), .Y(
        c0nm_b0m_v0m_n186) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u253 ( .A(c0nm_b0m_v0m_buffers3_11_), .Y(
        c0nm_b0m_v0m_n21) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u252 ( .A(c0nm_b0m_v0m_n50), .Y(
        c0nm_b0m_v0m_n190) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u251 ( .A0(c0nm_b0m_v0m_n193), .A1(
        c0nm_b0m_v0m_buffers0_11_), .B0(c0nm_b0m_v0m_n192), .B1(
        c0nm_b0m_v0m_n190), .Y(c0nm_b0m_v0m_n273) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u250 ( .A0(c0nm_b0m_v0m_n186), .A1(
        c0nm_b0m_v0m_n187), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n21), .C0(
        c0nm_b0m_v0m_n273), .Y(c0nm_b0m_headflit_11_) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u249 ( .A(c0nm_b0m_v0m_buffers2_2_), .Y(
        c0nm_b0m_v0m_n131) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u248 ( .A(c0nm_b0m_v0m_buffers3_2_), .Y(
        c0nm_b0m_v0m_n35) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u247 ( .A(c0nm_b0m_v0m_n59), .Y(
        c0nm_b0m_v0m_n134) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u246 ( .A0(c0nm_b0m_v0m_buffers0_2_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n134), 
        .Y(c0nm_b0m_v0m_n272) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u245 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n131), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n35), .C0(
        c0nm_b0m_v0m_n272), .Y(c0nm_headflit[2]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u244 ( .A(c0nm_b0m_v0m_buffers2_3_), .Y(
        c0nm_b0m_v0m_n138) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u243 ( .A(c0nm_b0m_v0m_buffers3_3_), .Y(
        c0nm_b0m_v0m_n38) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u242 ( .A(c0nm_b0m_v0m_n58), .Y(
        c0nm_b0m_v0m_n141) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u241 ( .A0(c0nm_b0m_v0m_buffers0_3_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n141), 
        .Y(c0nm_b0m_v0m_n271) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u240 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n138), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n38), .C0(
        c0nm_b0m_v0m_n271), .Y(c0nm_headflit[3]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u239 ( .A(c0nm_b0m_v0m_buffers2_4_), .Y(
        c0nm_b0m_v0m_n144) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u238 ( .A(c0nm_b0m_v0m_buffers3_4_), .Y(
        c0nm_b0m_v0m_n41) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u237 ( .A(c0nm_b0m_v0m_n57), .Y(
        c0nm_b0m_v0m_n147) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u236 ( .A0(c0nm_b0m_v0m_buffers0_4_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n147), 
        .Y(c0nm_b0m_v0m_n270) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u235 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n144), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n41), .C0(
        c0nm_b0m_v0m_n270), .Y(c0nm_headflit[4]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u234 ( .A(c0nm_b0m_v0m_buffers2_5_), .Y(
        c0nm_b0m_v0m_n150) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u233 ( .A(c0nm_b0m_v0m_buffers3_5_), .Y(
        c0nm_b0m_v0m_n44) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u232 ( .A(c0nm_b0m_v0m_n56), .Y(
        c0nm_b0m_v0m_n153) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u231 ( .A0(c0nm_b0m_v0m_buffers0_5_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n153), 
        .Y(c0nm_b0m_v0m_n269) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u230 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n150), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n44), .C0(
        c0nm_b0m_v0m_n269), .Y(c0nm_headflit[5]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u229 ( .A(c0nm_b0m_v0m_buffers2_6_), .Y(
        c0nm_b0m_v0m_n156) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u228 ( .A(c0nm_b0m_v0m_buffers3_6_), .Y(
        c0nm_b0m_v0m_n47) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u227 ( .A(c0nm_b0m_v0m_n55), .Y(
        c0nm_b0m_v0m_n159) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u226 ( .A0(c0nm_b0m_v0m_buffers0_6_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n159), 
        .Y(c0nm_b0m_v0m_n268) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u225 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n156), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n47), .C0(
        c0nm_b0m_v0m_n268), .Y(c0nm_headflit[6]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u224 ( .A(c0nm_b0m_v0m_buffers2_7_), .Y(
        c0nm_b0m_v0m_n162) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u223 ( .A(c0nm_b0m_v0m_buffers3_7_), .Y(
        c0nm_b0m_v0m_n62) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u222 ( .A(c0nm_b0m_v0m_n54), .Y(
        c0nm_b0m_v0m_n165) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u221 ( .A0(c0nm_b0m_v0m_buffers0_7_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n165), 
        .Y(c0nm_b0m_v0m_n267) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u220 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n162), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n62), .C0(
        c0nm_b0m_v0m_n267), .Y(c0nm_headflit[7]) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u219 ( .A(c0nm_b0m_v0m_buffers2_8_), .Y(
        c0nm_b0m_v0m_n168) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u218 ( .A(c0nm_b0m_v0m_buffers3_8_), .Y(
        c0nm_b0m_v0m_n65) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u217 ( .A(c0nm_b0m_v0m_n53), .Y(
        c0nm_b0m_v0m_n171) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u216 ( .A0(c0nm_b0m_v0m_buffers0_8_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n171), 
        .Y(c0nm_b0m_v0m_n266) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u215 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n168), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n65), .C0(
        c0nm_b0m_v0m_n266), .Y(c0nm_b0m_headflit_8_) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u214 ( .A(c0nm_b0m_v0m_buffers2_9_), .Y(
        c0nm_b0m_v0m_n174) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u213 ( .A(c0nm_b0m_v0m_buffers3_9_), .Y(
        c0nm_b0m_v0m_n68) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u212 ( .A(c0nm_b0m_v0m_n52), .Y(
        c0nm_b0m_v0m_n177) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u211 ( .A0(c0nm_b0m_v0m_buffers0_9_), .A1(
        c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n177), 
        .Y(c0nm_b0m_v0m_n265) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u210 ( .A0(c0nm_b0m_v0m_n187), .A1(
        c0nm_b0m_v0m_n174), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n68), .C0(
        c0nm_b0m_v0m_n265), .Y(c0nm_b0m_headflit_9_) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u209 ( .A(debitout_0), .B(reset), .Y(
        c0nm_b0m_v0m_n11) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u208 ( .A(c0nm_b0m_v0m_n11), .B(reset), .Y(
        c0nm_b0m_v0m_n10) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u207 ( .A0(c0nm_b0m_rdata[11]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_11_), 
        .Y(c0nm_b0m_v0m_n196) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u206 ( .A0(c0nm_b0m_rdata[10]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_10_), 
        .Y(c0nm_b0m_v0m_n197) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u205 ( .A0(c0nm_b0m_rdata[9]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_9_), 
        .Y(c0nm_b0m_v0m_n198) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u204 ( .A0(c0nm_b0m_rdata[8]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_8_), 
        .Y(c0nm_b0m_v0m_n199) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u203 ( .A0(c0nm_b0m_rdata[7]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[7]), .Y(
        c0nm_b0m_v0m_n200) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u202 ( .A0(c0nm_b0m_rdata[6]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[6]), .Y(
        c0nm_b0m_v0m_n201) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u201 ( .A0(c0nm_b0m_rdata[5]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[5]), .Y(
        c0nm_b0m_v0m_n202) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u200 ( .A0(c0nm_b0m_rdata[4]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[4]), .Y(
        c0nm_b0m_v0m_n203) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u199 ( .A0(c0nm_b0m_rdata[3]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[3]), .Y(
        c0nm_b0m_v0m_n204) );
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u198 ( .A0(c0nm_b0m_rdata[2]), .A1(
        c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[2]), .Y(
        c0nm_b0m_v0m_n205) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u197 ( .A(c0nm_b0m_v0m_n264), .B(
        c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n263) );
  MXT2_X0P5M_A12TR c0nm_b0m_v0m_u196 ( .A(c0nm_b0m_v0m_n263), .B(
        c0nm_b0m_rdata[1]), .S0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n206) );
  NAND2B_X0P5M_A12TR c0nm_b0m_v0m_u195 ( .AN(c0nm_headflit[0]), .B(
        c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n262) );
  MXT2_X0P5M_A12TR c0nm_b0m_v0m_u194 ( .A(c0nm_b0m_v0m_n262), .B(
        c0nm_b0m_rdata[0]), .S0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n207) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u193 ( .A(c0nm_b0m_v0m_tail_1_), .Y(
        c0nm_b0m_v0m_n7) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u192 ( .A(c0nm_b0m_v0m_tail_0_), .B(
        c0nm_b0m_v0m_n7), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n93) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u191 ( .A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_n1), 
        .Y(c0nm_b0m_v0m_n119) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u190 ( .A(c0nm_b0m_v0m_n119), .Y(
        c0nm_b0m_v0m_n135) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u189 ( .A(c0nm_b0m_v0m_tail_0_), .Y(
        c0nm_b0m_v0m_n3) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u188 ( .A(c0nm_b0m_v0m_tail_1_), .B(
        c0nm_b0m_v0m_n3), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n94) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u187 ( .A(c0nm_b0m_v0m_n94), .B(c0nm_b0m_n1), 
        .Y(c0nm_b0m_v0m_n121) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u186 ( .A(c0nm_b0m_v0m_n3), .B(
        c0nm_b0m_v0m_n7), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n95) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u185 ( .A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_n1), 
        .Y(c0nm_b0m_v0m_n120) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u184 ( .A0(c0nm_b0m_v0m_buffers2_11_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_11_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n194) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u183 ( .A(c0nm_b0m_v0m_n95), .B(
        c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n93), .Y(c0nm_b0m_v0m_n28) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u182 ( .A(c0nm_b0m_v0m_n28), .B(c0nm_b0m_n1), 
        .Y(c0nm_b0m_v0m_n128) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u181 ( .A0(c0nm_b0m_v0m_buffers3_11_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_n1), .B1(c0nm_b0m_wdata_11_), .Y(
        c0nm_b0m_v0m_n195) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u180 ( .A0(c0nm_b0m_v0m_n50), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n194), .C0(c0nm_b0m_v0m_n195), 
        .Y(c0nm_b0m_v0m_n19) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u179 ( .A(c0nm_b0m_v0m_n94), .Y(
        c0nm_b0m_v0m_n108) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u178 ( .A(c0nm_b0m_v0m_n108), .B(
        c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n129) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u177 ( .A(c0nm_b0m_v0m_n193), .Y(
        c0nm_b0m_v0m_n96) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u176 ( .A(c0nm_b0m_v0m_n192), .Y(
        c0nm_b0m_v0m_n104) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u175 ( .A(debitout_0), .Y(c0nm_b0m_v0m_n191) );
  NAND4_X0P5A_A12TR c0nm_b0m_v0m_u174 ( .A(c0nm_b0m_v0m_n96), .B(
        c0nm_b0m_v0m_n104), .C(c0nm_b0m_v0m_n187), .D(c0nm_b0m_v0m_n191), .Y(
        c0nm_b0m_v0m_n111) );
  OR2_X0P5M_A12TR c0nm_b0m_v0m_u173 ( .A(c0nm_b0m_v0m_n187), .B(debitout_0), 
        .Y(c0nm_b0m_v0m_n110) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u172 ( .A(c0nm_b0m_v0m_n96), .B(debitout_0), 
        .Y(c0nm_b0m_v0m_n115) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u171 ( .A(c0nm_b0m_v0m_n104), .B(debitout_0), 
        .Y(c0nm_b0m_v0m_n113) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u170 ( .A0(c0nm_b0m_v0m_n115), .A1(
        c0nm_b0m_v0m_buffers0_11_), .B0(c0nm_b0m_v0m_n113), .B1(
        c0nm_b0m_v0m_n190), .Y(c0nm_b0m_v0m_n189) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u169 ( .A0(c0nm_b0m_v0m_n21), .A1(
        c0nm_b0m_v0m_n111), .B0(c0nm_b0m_v0m_n186), .B1(c0nm_b0m_v0m_n110), 
        .C0(c0nm_b0m_v0m_n189), .Y(c0nm_b0m_v0m_n188) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u168 ( .A(c0nm_b0m_v0m_n188), .Y(
        c0nm_b0m_v0m_n17) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u167 ( .A(c0nm_b0m_v0m_n187), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n94), .Y(c0nm_b0m_v0m_n107) );
  OAI21_X0P5M_A12TR c0nm_b0m_v0m_u166 ( .A0(c0nm_b0m_v0m_n3), .A1(
        c0nm_b0m_v0m_n7), .B0(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n26) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u165 ( .A(c0nm_b0m_v0m_n26), .Y(
        c0nm_b0m_v0m_n72) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u164 ( .A(c0nm_b0m_v0m_n93), .B(
        c0nm_b0m_v0m_n95), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n109) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u163 ( .A(c0nm_b0m_v0m_n107), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n109), .Y(c0nm_b0m_v0m_n130) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u162 ( .A0(c0nm_b0m_v0m_n19), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n186), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n208)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u161 ( .A0(c0nm_b0m_v0m_buffers2_10_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_10_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n184) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u160 ( .A0(c0nm_b0m_v0m_buffers3_10_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_10_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n185) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u159 ( .A0(c0nm_b0m_v0m_n51), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n184), .C0(c0nm_b0m_v0m_n185), 
        .Y(c0nm_b0m_v0m_n70) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u158 ( .A0(c0nm_b0m_v0m_buffers0_10_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n183), 
        .Y(c0nm_b0m_v0m_n182) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u157 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n71), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n180), 
        .C0(c0nm_b0m_v0m_n182), .Y(c0nm_b0m_v0m_n181) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u156 ( .A(c0nm_b0m_v0m_n181), .Y(
        c0nm_b0m_v0m_n69) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u155 ( .A0(c0nm_b0m_v0m_n70), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n180), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n209)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u154 ( .A0(c0nm_b0m_v0m_buffers2_9_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_9_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n178) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u153 ( .A0(c0nm_b0m_v0m_buffers3_9_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_9_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n179) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u152 ( .A0(c0nm_b0m_v0m_n52), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n178), .C0(c0nm_b0m_v0m_n179), 
        .Y(c0nm_b0m_v0m_n67) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u151 ( .A0(c0nm_b0m_v0m_buffers0_9_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n177), 
        .Y(c0nm_b0m_v0m_n176) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u150 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n68), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n174), 
        .C0(c0nm_b0m_v0m_n176), .Y(c0nm_b0m_v0m_n175) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u149 ( .A(c0nm_b0m_v0m_n175), .Y(
        c0nm_b0m_v0m_n66) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u148 ( .A0(c0nm_b0m_v0m_n67), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n174), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n210)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u147 ( .A0(c0nm_b0m_v0m_buffers2_8_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_8_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n172) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u146 ( .A0(c0nm_b0m_v0m_buffers3_8_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_8_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n173) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u145 ( .A0(c0nm_b0m_v0m_n53), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n172), .C0(c0nm_b0m_v0m_n173), 
        .Y(c0nm_b0m_v0m_n64) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u144 ( .A0(c0nm_b0m_v0m_buffers0_8_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n171), 
        .Y(c0nm_b0m_v0m_n170) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u143 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n65), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n168), 
        .C0(c0nm_b0m_v0m_n170), .Y(c0nm_b0m_v0m_n169) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u142 ( .A(c0nm_b0m_v0m_n169), .Y(
        c0nm_b0m_v0m_n63) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u141 ( .A0(c0nm_b0m_v0m_n64), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n168), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n211)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u140 ( .A0(c0nm_b0m_v0m_buffers2_7_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_7_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n166) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u139 ( .A0(c0nm_b0m_v0m_buffers3_7_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_7_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n167) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u138 ( .A0(c0nm_b0m_v0m_n54), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n166), .C0(c0nm_b0m_v0m_n167), 
        .Y(c0nm_b0m_v0m_n49) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u137 ( .A0(c0nm_b0m_v0m_buffers0_7_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n165), 
        .Y(c0nm_b0m_v0m_n164) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u136 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n62), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n162), 
        .C0(c0nm_b0m_v0m_n164), .Y(c0nm_b0m_v0m_n163) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u135 ( .A(c0nm_b0m_v0m_n163), .Y(
        c0nm_b0m_v0m_n48) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u134 ( .A0(c0nm_b0m_v0m_n49), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n162), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n212)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u133 ( .A0(c0nm_b0m_v0m_buffers2_6_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_6_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n160) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u132 ( .A0(c0nm_b0m_v0m_buffers3_6_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_6_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n161) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u131 ( .A0(c0nm_b0m_v0m_n55), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n160), .C0(c0nm_b0m_v0m_n161), 
        .Y(c0nm_b0m_v0m_n46) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u130 ( .A0(c0nm_b0m_v0m_buffers0_6_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n159), 
        .Y(c0nm_b0m_v0m_n158) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u129 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n47), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n156), 
        .C0(c0nm_b0m_v0m_n158), .Y(c0nm_b0m_v0m_n157) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u128 ( .A(c0nm_b0m_v0m_n157), .Y(
        c0nm_b0m_v0m_n45) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u127 ( .A0(c0nm_b0m_v0m_n46), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n156), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n213)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u126 ( .A0(c0nm_b0m_v0m_buffers2_5_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_5_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n154) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u125 ( .A0(c0nm_b0m_v0m_buffers3_5_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_5_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n155) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u124 ( .A0(c0nm_b0m_v0m_n56), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n154), .C0(c0nm_b0m_v0m_n155), 
        .Y(c0nm_b0m_v0m_n43) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u123 ( .A0(c0nm_b0m_v0m_buffers0_5_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n153), 
        .Y(c0nm_b0m_v0m_n152) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u122 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n44), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n150), 
        .C0(c0nm_b0m_v0m_n152), .Y(c0nm_b0m_v0m_n151) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u121 ( .A(c0nm_b0m_v0m_n151), .Y(
        c0nm_b0m_v0m_n42) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u120 ( .A0(c0nm_b0m_v0m_n43), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n150), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n214)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u119 ( .A0(c0nm_b0m_v0m_buffers2_4_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_4_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n148) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u118 ( .A0(c0nm_b0m_v0m_buffers3_4_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_4_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n149) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u117 ( .A0(c0nm_b0m_v0m_n57), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n148), .C0(c0nm_b0m_v0m_n149), 
        .Y(c0nm_b0m_v0m_n40) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u116 ( .A0(c0nm_b0m_v0m_buffers0_4_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n147), 
        .Y(c0nm_b0m_v0m_n146) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u115 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n41), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n144), 
        .C0(c0nm_b0m_v0m_n146), .Y(c0nm_b0m_v0m_n145) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u114 ( .A(c0nm_b0m_v0m_n145), .Y(
        c0nm_b0m_v0m_n39) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u113 ( .A0(c0nm_b0m_v0m_n40), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n144), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n215)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u112 ( .A0(c0nm_b0m_v0m_buffers2_3_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_3_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n142) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u111 ( .A0(c0nm_b0m_v0m_buffers3_3_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_3_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n143) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u110 ( .A0(c0nm_b0m_v0m_n58), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n142), .C0(c0nm_b0m_v0m_n143), 
        .Y(c0nm_b0m_v0m_n37) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u109 ( .A0(c0nm_b0m_v0m_buffers0_3_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n141), 
        .Y(c0nm_b0m_v0m_n140) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u108 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n38), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n138), 
        .C0(c0nm_b0m_v0m_n140), .Y(c0nm_b0m_v0m_n139) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u107 ( .A(c0nm_b0m_v0m_n139), .Y(
        c0nm_b0m_v0m_n36) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u106 ( .A0(c0nm_b0m_v0m_n37), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n138), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n216)
         );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u105 ( .A0(c0nm_b0m_v0m_buffers2_2_), .A1(
        c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_2_), .B1(
        c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n136) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u104 ( .A0(c0nm_b0m_v0m_buffers3_2_), .A1(
        c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_2_), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n137) );
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u103 ( .A0(c0nm_b0m_v0m_n59), .A1(
        c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n136), .C0(c0nm_b0m_v0m_n137), 
        .Y(c0nm_b0m_v0m_n34) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u102 ( .A0(c0nm_b0m_v0m_buffers0_2_), .A1(
        c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n134), 
        .Y(c0nm_b0m_v0m_n133) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u101 ( .A0(c0nm_b0m_v0m_n111), .A1(
        c0nm_b0m_v0m_n35), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n131), 
        .C0(c0nm_b0m_v0m_n133), .Y(c0nm_b0m_v0m_n132) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u100 ( .A(c0nm_b0m_v0m_n132), .Y(
        c0nm_b0m_v0m_n33) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u99 ( .A0(c0nm_b0m_v0m_n34), .A1(
        c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n130), 
        .C0(c0nm_b0m_v0m_n131), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n217)
         );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u98 ( .A(c0nm_b0m_v0m_n128), .Y(
        c0nm_b0m_v0m_n116) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u97 ( .A0(c0nm_b0m_v0m_buffers0_1_), .A1(
        c0nm_b0m_v0m_n120), .B0(c0nm_b0m_v0m_buffers2_1_), .B1(
        c0nm_b0m_v0m_n121), .Y(c0nm_b0m_v0m_n126) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u96 ( .A0(c0nm_b0m_v0m_n119), .A1(
        c0nm_b0m_v0m_n125), .B0(flitin_0[1]), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n127) );
  OAI211_X0P5M_A12TR c0nm_b0m_v0m_u95 ( .A0(c0nm_b0m_v0m_n116), .A1(
        c0nm_b0m_v0m_n29), .B0(c0nm_b0m_v0m_n126), .C0(c0nm_b0m_v0m_n127), .Y(
        c0nm_b0m_v0m_n31) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u94 ( .A0(c0nm_b0m_v0m_n113), .A1(
        c0nm_b0m_v0m_n125), .B0(c0nm_b0m_v0m_buffers0_1_), .B1(
        c0nm_b0m_v0m_n115), .C0(debitout_0), .Y(c0nm_b0m_v0m_n124) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u93 ( .A0(c0nm_b0m_v0m_n110), .A1(
        c0nm_b0m_v0m_n122), .B0(c0nm_b0m_v0m_n111), .B1(c0nm_b0m_v0m_n29), 
        .C0(c0nm_b0m_v0m_n124), .Y(c0nm_b0m_v0m_n32) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u92 ( .A0(c0nm_b0m_v0m_n108), .A1(
        c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n109), .B1(c0nm_b0m_v0m_n32), .C0(
        reset), .Y(c0nm_b0m_v0m_n123) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u91 ( .A(c0nm_b0m_v0m_n122), .B(
        c0nm_b0m_v0m_n123), .S0(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n218) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u90 ( .A0(c0nm_b0m_v0m_buffers0_0_), .A1(
        c0nm_b0m_v0m_n120), .B0(c0nm_b0m_v0m_buffers2_0_), .B1(
        c0nm_b0m_v0m_n121), .Y(c0nm_b0m_v0m_n117) );
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u89 ( .A0(c0nm_b0m_v0m_n119), .A1(
        c0nm_b0m_v0m_n114), .B0(flitin_0[0]), .B1(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n118) );
  OAI211_X0P5M_A12TR c0nm_b0m_v0m_u88 ( .A0(c0nm_b0m_v0m_n116), .A1(
        c0nm_b0m_v0m_n23), .B0(c0nm_b0m_v0m_n117), .C0(c0nm_b0m_v0m_n118), .Y(
        c0nm_b0m_v0m_n25) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u87 ( .A0(c0nm_b0m_v0m_n113), .A1(
        c0nm_b0m_v0m_n114), .B0(c0nm_b0m_v0m_buffers0_0_), .B1(
        c0nm_b0m_v0m_n115), .C0(debitout_0), .Y(c0nm_b0m_v0m_n112) );
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u86 ( .A0(c0nm_b0m_v0m_n110), .A1(
        c0nm_b0m_v0m_n105), .B0(c0nm_b0m_v0m_n111), .B1(c0nm_b0m_v0m_n23), 
        .C0(c0nm_b0m_v0m_n112), .Y(c0nm_b0m_v0m_n27) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u85 ( .A0(c0nm_b0m_v0m_n108), .A1(
        c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n109), .B1(c0nm_b0m_v0m_n27), .C0(
        reset), .Y(c0nm_b0m_v0m_n106) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u84 ( .A(c0nm_b0m_v0m_n105), .B(
        c0nm_b0m_v0m_n106), .S0(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n219) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u83 ( .A(c0nm_b0m_v0m_n93), .Y(c0nm_b0m_v0m_n99) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u82 ( .A(c0nm_b0m_v0m_n99), .B(
        c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n102) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u81 ( .A(c0nm_b0m_v0m_n93), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n104), .Y(c0nm_b0m_v0m_n98) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u80 ( .A(c0nm_b0m_v0m_n95), .B(
        c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n100) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u79 ( .A(c0nm_b0m_v0m_n98), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n100), .Y(c0nm_b0m_v0m_n103) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u78 ( .A0(c0nm_b0m_v0m_n19), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n50), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n220) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u77 ( .A0(c0nm_b0m_v0m_n70), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n51), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n221) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u76 ( .A0(c0nm_b0m_v0m_n67), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n52), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n222) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u75 ( .A0(c0nm_b0m_v0m_n64), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n53), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n223) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u74 ( .A0(c0nm_b0m_v0m_n49), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n54), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n224) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u73 ( .A0(c0nm_b0m_v0m_n46), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n55), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n225) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u72 ( .A0(c0nm_b0m_v0m_n43), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n56), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n226) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u71 ( .A0(c0nm_b0m_v0m_n40), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n57), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n227) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u70 ( .A0(c0nm_b0m_v0m_n37), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n58), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n228) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u69 ( .A0(c0nm_b0m_v0m_n34), .A1(
        c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n103), 
        .C0(c0nm_b0m_v0m_n59), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n229) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u68 ( .A0(c0nm_b0m_v0m_n99), .A1(
        c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n100), .B1(c0nm_b0m_v0m_n32), .C0(
        reset), .Y(c0nm_b0m_v0m_n101) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u67 ( .A(c0nm_b0m_v0m_n60), .B(
        c0nm_b0m_v0m_n101), .S0(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n230) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u66 ( .A0(c0nm_b0m_v0m_n99), .A1(
        c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n100), .B1(c0nm_b0m_v0m_n27), .C0(
        reset), .Y(c0nm_b0m_v0m_n97) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u65 ( .A(c0nm_b0m_v0m_n61), .B(
        c0nm_b0m_v0m_n97), .S0(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n231) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u64 ( .A(c0nm_b0m_v0m_n95), .Y(c0nm_b0m_v0m_n77) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u63 ( .A(c0nm_b0m_v0m_n77), .B(
        c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n81) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u62 ( .A(c0nm_b0m_v0m_n95), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n96), .Y(c0nm_b0m_v0m_n76) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u61 ( .A(c0nm_b0m_v0m_n93), .B(
        c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n78) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u60 ( .A(c0nm_b0m_v0m_n76), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n78), .Y(c0nm_b0m_v0m_n82) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u59 ( .A(c0nm_b0m_v0m_buffers0_11_), .Y(
        c0nm_b0m_v0m_n92) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u58 ( .A0(c0nm_b0m_v0m_n19), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n92), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n232) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u57 ( .A(c0nm_b0m_v0m_buffers0_10_), .Y(
        c0nm_b0m_v0m_n91) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u56 ( .A0(c0nm_b0m_v0m_n70), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n91), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n233) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u55 ( .A(c0nm_b0m_v0m_buffers0_9_), .Y(
        c0nm_b0m_v0m_n90) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u54 ( .A0(c0nm_b0m_v0m_n67), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n90), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n234) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u53 ( .A(c0nm_b0m_v0m_buffers0_8_), .Y(
        c0nm_b0m_v0m_n89) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u52 ( .A0(c0nm_b0m_v0m_n64), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n89), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n235) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u51 ( .A(c0nm_b0m_v0m_buffers0_7_), .Y(
        c0nm_b0m_v0m_n88) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u50 ( .A0(c0nm_b0m_v0m_n49), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n88), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n236) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u49 ( .A(c0nm_b0m_v0m_buffers0_6_), .Y(
        c0nm_b0m_v0m_n87) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u48 ( .A0(c0nm_b0m_v0m_n46), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n87), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n237) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u47 ( .A(c0nm_b0m_v0m_buffers0_5_), .Y(
        c0nm_b0m_v0m_n86) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u46 ( .A0(c0nm_b0m_v0m_n43), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n86), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n238) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u45 ( .A(c0nm_b0m_v0m_buffers0_4_), .Y(
        c0nm_b0m_v0m_n85) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u44 ( .A0(c0nm_b0m_v0m_n40), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n85), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n239) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u43 ( .A(c0nm_b0m_v0m_buffers0_3_), .Y(
        c0nm_b0m_v0m_n84) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u42 ( .A0(c0nm_b0m_v0m_n37), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n84), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n240) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u41 ( .A(c0nm_b0m_v0m_buffers0_2_), .Y(
        c0nm_b0m_v0m_n83) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u40 ( .A0(c0nm_b0m_v0m_n34), .A1(
        c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n82), .C0(
        c0nm_b0m_v0m_n83), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n241) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u39 ( .A(c0nm_b0m_v0m_buffers0_1_), .Y(
        c0nm_b0m_v0m_n79) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u38 ( .A0(c0nm_b0m_v0m_n77), .A1(
        c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n78), .B1(c0nm_b0m_v0m_n32), .C0(
        reset), .Y(c0nm_b0m_v0m_n80) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u37 ( .A(c0nm_b0m_v0m_n79), .B(
        c0nm_b0m_v0m_n80), .S0(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n242) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u36 ( .A(c0nm_b0m_v0m_buffers0_0_), .Y(
        c0nm_b0m_v0m_n74) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u35 ( .A0(c0nm_b0m_v0m_n77), .A1(
        c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n78), .B1(c0nm_b0m_v0m_n27), .C0(
        reset), .Y(c0nm_b0m_v0m_n75) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u34 ( .A(c0nm_b0m_v0m_n74), .B(
        c0nm_b0m_v0m_n75), .S0(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n243) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u33 ( .A(c0nm_b0m_v0m_n72), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n73), .Y(c0nm_b0m_v0m_n22) );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u32 ( .A(c0nm_b0m_v0m_n22), .B(
        c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n28), .Y(c0nm_b0m_v0m_n18) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u31 ( .A(c0nm_b0m_v0m_n26), .B(
        c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n20) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u30 ( .A0(c0nm_b0m_v0m_n69), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n70), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n71), .Y(c0nm_b0m_v0m_n244) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u29 ( .A0(c0nm_b0m_v0m_n66), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n67), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n68), .Y(c0nm_b0m_v0m_n245) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u28 ( .A0(c0nm_b0m_v0m_n63), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n64), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n65), .Y(c0nm_b0m_v0m_n246) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u27 ( .A0(c0nm_b0m_v0m_n48), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n49), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n62), .Y(c0nm_b0m_v0m_n247) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u26 ( .A0(c0nm_b0m_v0m_n45), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n46), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n47), .Y(c0nm_b0m_v0m_n248) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u25 ( .A0(c0nm_b0m_v0m_n42), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n43), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n44), .Y(c0nm_b0m_v0m_n249) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u24 ( .A0(c0nm_b0m_v0m_n39), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n40), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n41), .Y(c0nm_b0m_v0m_n250) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u23 ( .A0(c0nm_b0m_v0m_n36), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n37), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n38), .Y(c0nm_b0m_v0m_n251) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u22 ( .A0(c0nm_b0m_v0m_n33), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n34), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n35), .Y(c0nm_b0m_v0m_n252) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u21 ( .A0(c0nm_b0m_v0m_n31), .A1(
        c0nm_b0m_v0m_n26), .B0(c0nm_b0m_v0m_n32), .B1(c0nm_b0m_v0m_n28), .C0(
        reset), .Y(c0nm_b0m_v0m_n30) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u20 ( .A(c0nm_b0m_v0m_n29), .B(
        c0nm_b0m_v0m_n30), .S0(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n253) );
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u19 ( .A0(c0nm_b0m_v0m_n25), .A1(
        c0nm_b0m_v0m_n26), .B0(c0nm_b0m_v0m_n27), .B1(c0nm_b0m_v0m_n28), .C0(
        reset), .Y(c0nm_b0m_v0m_n24) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u18 ( .A(c0nm_b0m_v0m_n23), .B(
        c0nm_b0m_v0m_n24), .S0(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n254) );
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u17 ( .A0(c0nm_b0m_v0m_n17), .A1(
        c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n19), .B1(c0nm_b0m_v0m_n20), .C0(
        c0nm_b0m_v0m_n21), .C1(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n255) );
  AOI21_X0P5M_A12TR c0nm_b0m_v0m_u16 ( .A0(c0nm_b0m_v0m_n4), .A1(
        c0nm_b0m_v0m_n16), .B0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n12) );
  OA21A1OI2_X0P5M_A12TR c0nm_b0m_v0m_u15 ( .A0(reset), .A1(
        c0nm_b0m_v0m_head_1_), .B0(c0nm_b0m_v0m_n12), .C0(c0nm_b0m_v0m_n15), 
        .Y(c0nm_b0m_v0m_n256) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u14 ( .A(c0nm_b0m_v0m_n10), .B(
        c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n13) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u13 ( .A(c0nm_b0m_v0m_head_1_), .Y(
        c0nm_b0m_v0m_n14) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u12 ( .A(c0nm_b0m_v0m_n12), .B(
        c0nm_b0m_v0m_n13), .S0(c0nm_b0m_v0m_n14), .Y(c0nm_b0m_v0m_n257) );
  MXT2_X0P5M_A12TR c0nm_b0m_v0m_u11 ( .A(c0nm_b0m_v0m_n10), .B(
        c0nm_b0m_v0m_n11), .S0(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n258) );
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u10 ( .A(reset), .B(c0nm_b0m_n1), .Y(
        c0nm_b0m_v0m_n8) );
  AOI21_X0P5M_A12TR c0nm_b0m_v0m_u9 ( .A0(c0nm_b0m_v0m_n3), .A1(
        c0nm_b0m_v0m_n4), .B0(c0nm_b0m_v0m_n8), .Y(c0nm_b0m_v0m_n5) );
  OA21A1OI2_X0P5M_A12TR c0nm_b0m_v0m_u8 ( .A0(c0nm_b0m_v0m_tail_1_), .A1(reset), .B0(c0nm_b0m_v0m_n5), .C0(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n259) );
  INV_X0P5B_A12TR c0nm_b0m_v0m_u7 ( .A(c0nm_b0m_v0m_n8), .Y(c0nm_b0m_v0m_n1)
         );
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u6 ( .A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), 
        .C(c0nm_b0m_v0m_tail_0_), .Y(c0nm_b0m_v0m_n6) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u5 ( .A(c0nm_b0m_v0m_n5), .B(c0nm_b0m_v0m_n6), 
        .S0(c0nm_b0m_v0m_n7), .Y(c0nm_b0m_v0m_n260) );
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u4 ( .A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), 
        .Y(c0nm_b0m_v0m_n2) );
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u3 ( .A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n2), 
        .S0(c0nm_b0m_v0m_n3), .Y(c0nm_b0m_v0m_n261) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_tail_reg_2_ ( .D(c0nm_b0m_v0m_n259), .CK(clk), 
        .QN(c0nm_b0m_v0m_n9) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_2_ ( .D(c0nm_b0m_v0m_n229), .CK(
        clk), .QN(c0nm_b0m_v0m_n59) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_3_ ( .D(c0nm_b0m_v0m_n228), .CK(
        clk), .QN(c0nm_b0m_v0m_n58) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_4_ ( .D(c0nm_b0m_v0m_n227), .CK(
        clk), .QN(c0nm_b0m_v0m_n57) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_5_ ( .D(c0nm_b0m_v0m_n226), .CK(
        clk), .QN(c0nm_b0m_v0m_n56) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_6_ ( .D(c0nm_b0m_v0m_n225), .CK(
        clk), .QN(c0nm_b0m_v0m_n55) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_7_ ( .D(c0nm_b0m_v0m_n224), .CK(
        clk), .QN(c0nm_b0m_v0m_n54) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_8_ ( .D(c0nm_b0m_v0m_n223), .CK(
        clk), .QN(c0nm_b0m_v0m_n53) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_9_ ( .D(c0nm_b0m_v0m_n222), .CK(
        clk), .QN(c0nm_b0m_v0m_n52) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_10_ ( .D(c0nm_b0m_v0m_n221), .CK(
        clk), .QN(c0nm_b0m_v0m_n51) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_11_ ( .D(c0nm_b0m_v0m_n220), .CK(
        clk), .QN(c0nm_b0m_v0m_n50) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_0_ ( .D(c0nm_b0m_v0m_n231), .CK(
        clk), .QN(c0nm_b0m_v0m_n61) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_1_ ( .D(c0nm_b0m_v0m_n230), .CK(
        clk), .QN(c0nm_b0m_v0m_n60) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_1_ ( .D(c0nm_b0m_v0m_n257), .CK(clk), 
        .Q(c0nm_b0m_v0m_head_1_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_0_ ( .D(c0nm_b0m_v0m_n258), .CK(clk), 
        .Q(c0nm_b0m_v0m_head_0_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_tailout_reg ( .D(c0nm_b0m_v0m_n1710), .CK(clk), 
        .Q(tailout_0) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_11_ ( .D(c0nm_b0m_v0m_n232), .CK(
        clk), .Q(c0nm_b0m_v0m_buffers0_11_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_0_ ( .D(c0nm_b0m_v0m_n243), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_0_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_1_ ( .D(c0nm_b0m_v0m_n242), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_1_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_2_ ( .D(c0nm_b0m_v0m_n241), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_2_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_3_ ( .D(c0nm_b0m_v0m_n240), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_3_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_4_ ( .D(c0nm_b0m_v0m_n239), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_4_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_5_ ( .D(c0nm_b0m_v0m_n238), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_5_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_6_ ( .D(c0nm_b0m_v0m_n237), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_6_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_7_ ( .D(c0nm_b0m_v0m_n236), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_7_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_8_ ( .D(c0nm_b0m_v0m_n235), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_8_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_9_ ( .D(c0nm_b0m_v0m_n234), .CK(clk), .Q(c0nm_b0m_v0m_buffers0_9_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_10_ ( .D(c0nm_b0m_v0m_n233), .CK(
        clk), .Q(c0nm_b0m_v0m_buffers0_10_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_2_ ( .D(c0nm_b0m_v0m_n256), .CK(clk), 
        .Q(c0nm_b0m_v0m_head_2_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_tail_reg_0_ ( .D(c0nm_b0m_v0m_n261), .CK(clk), 
        .Q(c0nm_b0m_v0m_tail_0_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_tail_reg_1_ ( .D(c0nm_b0m_v0m_n260), .CK(clk), 
        .Q(c0nm_b0m_v0m_tail_1_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_2_ ( .D(c0nm_b0m_v0m_n217), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_2_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_2_ ( .D(c0nm_b0m_v0m_n252), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_2_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_3_ ( .D(c0nm_b0m_v0m_n216), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_3_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_3_ ( .D(c0nm_b0m_v0m_n251), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_3_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_4_ ( .D(c0nm_b0m_v0m_n215), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_4_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_4_ ( .D(c0nm_b0m_v0m_n250), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_4_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_5_ ( .D(c0nm_b0m_v0m_n214), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_5_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_5_ ( .D(c0nm_b0m_v0m_n249), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_5_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_6_ ( .D(c0nm_b0m_v0m_n213), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_6_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_6_ ( .D(c0nm_b0m_v0m_n248), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_6_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_7_ ( .D(c0nm_b0m_v0m_n212), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_7_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_7_ ( .D(c0nm_b0m_v0m_n247), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_7_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_8_ ( .D(c0nm_b0m_v0m_n211), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_8_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_8_ ( .D(c0nm_b0m_v0m_n246), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_8_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_9_ ( .D(c0nm_b0m_v0m_n210), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_9_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_9_ ( .D(c0nm_b0m_v0m_n245), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_9_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_10_ ( .D(c0nm_b0m_v0m_n209), .CK(
        clk), .Q(c0nm_b0m_v0m_buffers2_10_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_10_ ( .D(c0nm_b0m_v0m_n244), .CK(
        clk), .Q(c0nm_b0m_v0m_buffers3_10_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_11_ ( .D(c0nm_b0m_v0m_n208), .CK(
        clk), .Q(c0nm_b0m_v0m_buffers2_11_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_11_ ( .D(c0nm_b0m_v0m_n255), .CK(
        clk), .Q(c0nm_b0m_v0m_buffers3_11_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_0_ ( .D(c0nm_b0m_v0m_n219), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_0_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_1_ ( .D(c0nm_b0m_v0m_n218), .CK(clk), .Q(c0nm_b0m_v0m_buffers2_1_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_0_ ( .D(c0nm_b0m_v0m_n207), .CK(clk), 
        .Q(c0nm_b0m_rdata[0]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_1_ ( .D(c0nm_b0m_v0m_n206), .CK(clk), 
        .Q(c0nm_b0m_rdata[1]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_10_ ( .D(c0nm_b0m_v0m_n197), .CK(clk), 
        .Q(c0nm_b0m_rdata[10]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_11_ ( .D(c0nm_b0m_v0m_n196), .CK(clk), 
        .Q(c0nm_b0m_rdata[11]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_2_ ( .D(c0nm_b0m_v0m_n205), .CK(clk), 
        .Q(c0nm_b0m_rdata[2]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_3_ ( .D(c0nm_b0m_v0m_n204), .CK(clk), 
        .Q(c0nm_b0m_rdata[3]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_4_ ( .D(c0nm_b0m_v0m_n203), .CK(clk), 
        .Q(c0nm_b0m_rdata[4]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_5_ ( .D(c0nm_b0m_v0m_n202), .CK(clk), 
        .Q(c0nm_b0m_rdata[5]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_6_ ( .D(c0nm_b0m_v0m_n201), .CK(clk), 
        .Q(c0nm_b0m_rdata[6]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_7_ ( .D(c0nm_b0m_v0m_n200), .CK(clk), 
        .Q(c0nm_b0m_rdata[7]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_8_ ( .D(c0nm_b0m_v0m_n199), .CK(clk), 
        .Q(c0nm_b0m_rdata[8]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_9_ ( .D(c0nm_b0m_v0m_n198), .CK(clk), 
        .Q(c0nm_b0m_rdata[9]) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_0_ ( .D(c0nm_b0m_v0m_n254), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_0_) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_1_ ( .D(c0nm_b0m_v0m_n253), .CK(clk), .Q(c0nm_b0m_v0m_buffers3_1_) );
  INV_X0P5B_A12TR c0nm_r0m_u20 ( .A(currx[2]), .Y(c0nm_r0m_n4) );
  INV_X0P5B_A12TR c0nm_r0m_u19 ( .A(c0nm_headflit[5]), .Y(c0nm_r0m_n9) );
  OR2_X0P5M_A12TR c0nm_r0m_u18 ( .A(currx[0]), .B(c0nm_r0m_n9), .Y(
        c0nm_r0m_n15) );
  INV_X0P5B_A12TR c0nm_r0m_u17 ( .A(c0nm_headflit[6]), .Y(c0nm_r0m_n8) );
  AND2_X0P5M_A12TR c0nm_r0m_u16 ( .A(c0nm_r0m_n15), .B(currx[1]), .Y(
        c0nm_r0m_n16) );
  OA21A1OI2_X0P5M_A12TR c0nm_r0m_u15 ( .A0(currx[1]), .A1(c0nm_r0m_n15), .B0(
        c0nm_r0m_n8), .C0(c0nm_r0m_n16), .Y(c0nm_r0m_n6) );
  AOI2XB1_X0P5M_A12TR c0nm_r0m_u14 ( .A1N(curry[1]), .A0(c0nm_headflit[3]), 
        .B0(c0nm_headflit[2]), .Y(c0nm_r0m_n13) );
  INV_X0P5B_A12TR c0nm_r0m_u13 ( .A(c0nm_headflit[3]), .Y(c0nm_r0m_n14) );
  AOI22_X0P5M_A12TR c0nm_r0m_u12 ( .A0(c0nm_r0m_n13), .A1(curry[0]), .B0(
        curry[1]), .B1(c0nm_r0m_n14), .Y(c0nm_r0m_n12) );
  AOI2XB1_X0P5M_A12TR c0nm_r0m_u11 ( .A1N(curry[2]), .A0(c0nm_headflit[4]), 
        .B0(c0nm_r0m_n12), .Y(c0nm_r0m_n11) );
  AOI2XB1_X0P5M_A12TR c0nm_r0m_u10 ( .A1N(c0nm_headflit[4]), .A0(curry[2]), 
        .B0(c0nm_r0m_n11), .Y(c0nm_r0m_n10) );
  AOI221_X0P5M_A12TR c0nm_r0m_u9 ( .A0(currx[1]), .A1(c0nm_r0m_n8), .B0(
        currx[0]), .B1(c0nm_r0m_n9), .C0(c0nm_r0m_n10), .Y(c0nm_r0m_n7) );
  OAI22_X0P5M_A12TR c0nm_r0m_u8 ( .A0(c0nm_r0m_n6), .A1(c0nm_r0m_n7), .B0(
        c0nm_headflit[7]), .B1(c0nm_r0m_n4), .Y(c0nm_r0m_n5) );
  AO1B2_X0P5M_A12TR c0nm_r0m_u7 ( .B0(c0nm_r0m_n4), .B1(c0nm_headflit[7]), 
        .A0N(c0nm_r0m_n5), .Y(c0nm_r0m_n3) );
  INV_X0P5B_A12TR c0nm_r0m_u6 ( .A(c0nm_n1), .Y(c0nm_r0m_n1) );
  NOR3_X0P5A_A12TR c0nm_r0m_u5 ( .A(c0nm_r0m_n3), .B(reset), .C(c0nm_r0m_n1), 
        .Y(c0nm_r0m_n100) );
  INV_X0P5B_A12TR c0nm_r0m_u4 ( .A(c0nm_r0m_n3), .Y(c0nm_r0m_n2) );
  NOR3_X0P5A_A12TR c0nm_r0m_u3 ( .A(c0nm_r0m_n1), .B(reset), .C(c0nm_r0m_n2), 
        .Y(c0nm_r0m_n110) );
  DFFQ_X1M_A12TR c0nm_r0m_vc_req_reg_0_ ( .D(c0nm_r0m_n100), .CK(clk), .Q(
        c0nm_routewire[0]) );
  DFFQ_X1M_A12TR c0nm_r0m_vc_req_reg_1_ ( .D(c0nm_r0m_n110), .CK(clk), .Q(
        c0nm_routewire[1]) );
  INV_X0P5B_A12TR c0nm_v0m_u40 ( .A(c0nm_v0m_state_status_1_), .Y(c0nm_v0m_n29) );
  OAI211_X0P5M_A12TR c0nm_v0m_u39 ( .A0(swalloc_resp_0[1]), .A1(
        swalloc_resp_0[0]), .B0(c0nm_v0m_n29), .C0(c0nm_v0m_state_status_0_), 
        .Y(c0nm_v0m_n5) );
  NOR2_X0P5A_A12TR c0nm_v0m_u38 ( .A(reset), .B(tailout_0), .Y(c0nm_v0m_n8) );
  AO1B2_X0P5M_A12TR c0nm_v0m_u37 ( .B0(c0nm_v0m_n5), .B1(
        c0nm_v0m_state_status_0_), .A0N(c0nm_v0m_n8), .Y(c0nm_v0m_n57) );
  OA211_X0P5M_A12TR c0nm_v0m_u36 ( .A0(c0nm_routewire[1]), .A1(
        c0nm_routewire[0]), .B0(c0nm_v0m_state_status_0_), .C0(
        c0nm_v0m_state_status_1_), .Y(c0nm_v0m_n4) );
  AO21A1AI2_X0P5M_A12TR c0nm_v0m_u35 ( .A0(c0nm_v0m_n29), .A1(c0nm_v0m_n5), 
        .B0(c0nm_v0m_n4), .C0(c0nm_v0m_n8), .Y(c0nm_v0m_n58) );
  INV_X0P5B_A12TR c0nm_v0m_u34 ( .A(c0nm_v0m_state_queuelen_0_), .Y(
        c0nm_v0m_n23) );
  INV_X0P5B_A12TR c0nm_v0m_u33 ( .A(c0nm_v0m_full), .Y(c0nm_v0m_n26) );
  OAI31_X0P5M_A12TR c0nm_v0m_u32 ( .A0(c0nm_v0m_n29), .A1(tailout_0), .A2(
        c0nm_v0m_state_status_0_), .B0(c0nm_v0m_n5), .Y(c0nm_v0m_n28) );
  OAI31_X0P5M_A12TR c0nm_v0m_u31 ( .A0(c0nm_v0m_state_queuelen_0_), .A1(
        c0nm_v0m_state_queuelen_2_), .A2(c0nm_v0m_state_queuelen_1_), .B0(
        c0nm_v0m_n28), .Y(c0nm_v0m_n9) );
  NOR2_X0P5A_A12TR c0nm_v0m_u30 ( .A(c0nm_v0m_n9), .B(c0nm_n2), .Y(
        c0nm_v0m_n13) );
  INV_X0P5B_A12TR c0nm_v0m_u29 ( .A(c0nm_v0m_state_queuelen_2_), .Y(
        c0nm_v0m_n17) );
  NAND3_X0P5A_A12TR c0nm_v0m_u28 ( .A(c0nm_v0m_state_queuelen_0_), .B(
        c0nm_v0m_n17), .C(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n14) );
  NAND3_X0P5A_A12TR c0nm_v0m_u27 ( .A(c0nm_v0m_n14), .B(c0nm_v0m_n9), .C(
        c0nm_n2), .Y(c0nm_v0m_n18) );
  INV_X0P5B_A12TR c0nm_v0m_u26 ( .A(c0nm_v0m_n18), .Y(c0nm_v0m_n22) );
  AOI21_X0P5M_A12TR c0nm_v0m_u25 ( .A0(c0nm_v0m_n26), .A1(c0nm_v0m_n13), .B0(
        c0nm_v0m_n22), .Y(c0nm_v0m_n24) );
  XNOR2_X0P5M_A12TR c0nm_v0m_u24 ( .A(c0nm_v0m_n23), .B(c0nm_v0m_n24), .Y(
        c0nm_v0m_n27) );
  NOR2_X0P5A_A12TR c0nm_v0m_u23 ( .A(reset), .B(c0nm_v0m_n27), .Y(c0nm_v0m_n61) );
  NAND2_X0P5A_A12TR c0nm_v0m_u22 ( .A(c0nm_v0m_n13), .B(c0nm_v0m_n26), .Y(
        c0nm_v0m_n25) );
  MXIT2_X0P5M_A12TR c0nm_v0m_u21 ( .A(c0nm_v0m_n18), .B(c0nm_v0m_n25), .S0(
        c0nm_v0m_n23), .Y(c0nm_v0m_n20) );
  AOI21_X0P5M_A12TR c0nm_v0m_u20 ( .A0(c0nm_v0m_n23), .A1(c0nm_v0m_n22), .B0(
        c0nm_v0m_n24), .Y(c0nm_v0m_n16) );
  OAI21_X0P5M_A12TR c0nm_v0m_u19 ( .A0(c0nm_v0m_n22), .A1(c0nm_v0m_n23), .B0(
        c0nm_v0m_n16), .Y(c0nm_v0m_n21) );
  MXIT2_X0P5M_A12TR c0nm_v0m_u18 ( .A(c0nm_v0m_n20), .B(c0nm_v0m_n21), .S0(
        c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n19) );
  NOR2_X0P5A_A12TR c0nm_v0m_u17 ( .A(reset), .B(c0nm_v0m_n19), .Y(c0nm_v0m_n62) );
  MXIT2_X0P5M_A12TR c0nm_v0m_u16 ( .A(c0nm_v0m_state_queuelen_0_), .B(
        c0nm_v0m_n18), .S0(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n15) );
  AOI211_X0P5M_A12TR c0nm_v0m_u15 ( .A0(c0nm_v0m_n15), .A1(c0nm_v0m_n16), .B0(
        c0nm_v0m_n17), .C0(reset), .Y(c0nm_v0m_n63) );
  INV_X0P5B_A12TR c0nm_v0m_u14 ( .A(c0nm_v0m_n14), .Y(c0nm_v0m_n11) );
  INV_X0P5B_A12TR c0nm_v0m_u13 ( .A(c0nm_v0m_n13), .Y(c0nm_v0m_n12) );
  AOI32_X0P5M_A12TR c0nm_v0m_u12 ( .A0(c0nm_v0m_n11), .A1(c0nm_v0m_n9), .A2(
        c0nm_n2), .B0(c0nm_v0m_full), .B1(c0nm_v0m_n12), .Y(c0nm_v0m_n10) );
  NOR2_X0P5A_A12TR c0nm_v0m_u11 ( .A(reset), .B(c0nm_v0m_n10), .Y(c0nm_v0m_n64) );
  INV_X0P5B_A12TR c0nm_v0m_u10 ( .A(c0nm_v0m_n9), .Y(debitout_0) );
  INV_X0P5B_A12TR c0nm_v0m_u9 ( .A(c0nm_v0m_n8), .Y(c0nm_v0m_n1) );
  AND2_X0P5M_A12TR c0nm_v0m_u8 ( .A(swalloc_req_0[0]), .B(c0nm_v0m_n5), .Y(
        c0nm_v0m_n7) );
  MXIT2_X0P5M_A12TR c0nm_v0m_u7 ( .A(c0nm_v0m_n7), .B(c0nm_routewire[0]), .S0(
        c0nm_v0m_n4), .Y(c0nm_v0m_n6) );
  NOR2_X0P5A_A12TR c0nm_v0m_u6 ( .A(c0nm_v0m_n1), .B(c0nm_v0m_n6), .Y(
        c0nm_v0m_n30) );
  AND2_X0P5M_A12TR c0nm_v0m_u5 ( .A(swalloc_req_0[1]), .B(c0nm_v0m_n5), .Y(
        c0nm_v0m_n3) );
  MXIT2_X0P5M_A12TR c0nm_v0m_u4 ( .A(c0nm_v0m_n3), .B(c0nm_routewire[1]), .S0(
        c0nm_v0m_n4), .Y(c0nm_v0m_n2) );
  NOR2_X0P5A_A12TR c0nm_v0m_u3 ( .A(c0nm_v0m_n1), .B(c0nm_v0m_n2), .Y(
        c0nm_v0m_n31) );
  DFFQ_X1M_A12TR c0nm_v0m_state_queuelen_reg_1_ ( .D(c0nm_v0m_n62), .CK(clk), 
        .Q(c0nm_v0m_state_queuelen_1_) );
  DFFQ_X1M_A12TR c0nm_v0m_state_queuelen_reg_0_ ( .D(c0nm_v0m_n61), .CK(clk), 
        .Q(c0nm_v0m_state_queuelen_0_) );
  DFFQ_X1M_A12TR c0nm_v0m_state_status_reg_0_ ( .D(c0nm_v0m_n57), .CK(clk), 
        .Q(c0nm_v0m_state_status_0_) );
  DFFQ_X1M_A12TR c0nm_v0m_state_swreq_reg_1_ ( .D(c0nm_v0m_n31), .CK(clk), .Q(
        swalloc_req_0[1]) );
  DFFQ_X1M_A12TR c0nm_v0m_state_swreq_reg_0_ ( .D(c0nm_v0m_n30), .CK(clk), .Q(
        swalloc_req_0[0]) );
  DFFQ_X1M_A12TR c0nm_v0m_state_queuelen_reg_2_ ( .D(c0nm_v0m_n63), .CK(clk), 
        .Q(c0nm_v0m_state_queuelen_2_) );
  DFFQ_X1M_A12TR c0nm_v0m_full_reg ( .D(c0nm_v0m_n64), .CK(clk), .Q(
        c0nm_v0m_full) );
  DFFQ_X1M_A12TR c0nm_v0m_state_status_reg_1_ ( .D(c0nm_v0m_n58), .CK(clk), 
        .Q(c0nm_v0m_state_status_1_) );
  NOR2B_X0P5M_A12TR c0sm_u5 ( .AN(debitout_1), .B(reset), .Y(creditout_1) );
  NOR2B_X0P5M_A12TR c0sm_u4 ( .AN(c0sm_headflit[1]), .B(c0sm_headflit[0]), .Y(
        c0sm_n4) );
  NAND2_X0P5A_A12TR c0sm_u3 ( .A(flitin_1[1]), .B(flitin_1[0]), .Y(c0sm_n3) );
  TIELO_X1M_A12TR c0sm_u2 ( .Y(c0sm__logic0_) );
  NOR2B_X0P5M_A12TR c0sm_b0m_u27 ( .AN(debitout_1), .B(reset), .Y(c0sm_b0m_n9)
         );
  NAND2B_X0P5M_A12TR c0sm_b0m_u26 ( .AN(c0sm_b0m_rdata[0]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[0]) );
  AND2_X0P5M_A12TR c0sm_b0m_u25 ( .A(c0sm_b0m_rdata[10]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[10]) );
  AND2_X0P5M_A12TR c0sm_b0m_u24 ( .A(c0sm_b0m_rdata[11]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[11]) );
  NAND2B_X0P5M_A12TR c0sm_b0m_u23 ( .AN(c0sm_b0m_rdata[1]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[1]) );
  AND2_X0P5M_A12TR c0sm_b0m_u22 ( .A(c0sm_b0m_rdata[2]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[2]) );
  AND2_X0P5M_A12TR c0sm_b0m_u21 ( .A(c0sm_b0m_rdata[3]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[3]) );
  AND2_X0P5M_A12TR c0sm_b0m_u20 ( .A(c0sm_b0m_rdata[4]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[4]) );
  AND2_X0P5M_A12TR c0sm_b0m_u19 ( .A(c0sm_b0m_rdata[5]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[5]) );
  AND2_X0P5M_A12TR c0sm_b0m_u18 ( .A(c0sm_b0m_rdata[6]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[6]) );
  AND2_X0P5M_A12TR c0sm_b0m_u17 ( .A(c0sm_b0m_rdata[7]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[7]) );
  AND2_X0P5M_A12TR c0sm_b0m_u16 ( .A(c0sm_b0m_rdata[8]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[8]) );
  AND2_X0P5M_A12TR c0sm_b0m_u15 ( .A(c0sm_b0m_rdata[9]), .B(
        c0sm_b0m_dqenablereg), .Y(flitout_switch_1[9]) );
  NAND2_X0P5A_A12TR c0sm_b0m_u14 ( .A(flitin_1[1]), .B(flitin_1[0]), .Y(
        c0sm_b0m_n2) );
  AND2_X0P5M_A12TR c0sm_b0m_u13 ( .A(flitin_1[10]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_10_) );
  AND2_X0P5M_A12TR c0sm_b0m_u12 ( .A(flitin_1[11]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_11_) );
  AND2_X0P5M_A12TR c0sm_b0m_u11 ( .A(flitin_1[2]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_2_) );
  AND2_X0P5M_A12TR c0sm_b0m_u10 ( .A(flitin_1[3]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_3_) );
  AND2_X0P5M_A12TR c0sm_b0m_u9 ( .A(flitin_1[4]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_4_) );
  AND2_X0P5M_A12TR c0sm_b0m_u8 ( .A(flitin_1[5]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_5_) );
  AND2_X0P5M_A12TR c0sm_b0m_u7 ( .A(flitin_1[6]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_6_) );
  AND2_X0P5M_A12TR c0sm_b0m_u6 ( .A(flitin_1[7]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_7_) );
  AND2_X0P5M_A12TR c0sm_b0m_u5 ( .A(flitin_1[8]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_8_) );
  AND2_X0P5M_A12TR c0sm_b0m_u4 ( .A(flitin_1[9]), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_wdata_9_) );
  TIELO_X1M_A12TR c0sm_b0m_u3 ( .Y(c0sm_b0m__logic0_) );
  DFFQ_X1M_A12TR c0sm_b0m_dqenablereg_reg ( .D(c0sm_b0m_n9), .CK(clk), .Q(
        c0sm_b0m_dqenablereg) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u278 ( .A(c0sm_b0m_v0m_head_0_), .Y(
        c0sm_b0m_v0m_n16) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u277 ( .A(c0sm_b0m_v0m_head_2_), .Y(
        c0sm_b0m_v0m_n15) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u276 ( .A(c0sm_b0m_v0m_n16), .B(
        c0sm_b0m_v0m_n15), .C(c0sm_b0m_v0m_head_1_), .Y(c0sm_b0m_v0m_n187) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u275 ( .A(c0sm_b0m_v0m_buffers2_0_), .Y(
        c0sm_b0m_v0m_n105) );
  AOI21_X0P5M_A12TR c0sm_b0m_v0m_u274 ( .A0(c0sm_b0m_v0m_head_0_), .A1(
        c0sm_b0m_v0m_head_1_), .B0(c0sm_b0m_v0m_head_2_), .Y(c0sm_b0m_v0m_n73)
         );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u273 ( .A(c0sm_b0m_v0m_buffers3_0_), .Y(
        c0sm_b0m_v0m_n23) );
  NOR3_X0P5A_A12TR c0sm_b0m_v0m_u272 ( .A(c0sm_b0m_v0m_head_1_), .B(
        c0sm_b0m_v0m_head_2_), .C(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n193)
         );
  NOR3_X0P5A_A12TR c0sm_b0m_v0m_u271 ( .A(c0sm_b0m_v0m_head_1_), .B(
        c0sm_b0m_v0m_head_2_), .C(c0sm_b0m_v0m_n16), .Y(c0sm_b0m_v0m_n192) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u270 ( .A(c0sm_b0m_v0m_n343), .Y(
        c0sm_b0m_v0m_n114) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u269 ( .A0(c0sm_b0m_v0m_buffers0_0_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n114), 
        .Y(c0sm_b0m_v0m_n276) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u268 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n105), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n23), .C0(
        c0sm_b0m_v0m_n276), .Y(c0sm_headflit[0]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u267 ( .A(c0sm_b0m_v0m_buffers2_1_), .Y(
        c0sm_b0m_v0m_n122) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u266 ( .A(c0sm_b0m_v0m_buffers3_1_), .Y(
        c0sm_b0m_v0m_n29) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u265 ( .A(c0sm_b0m_v0m_n344), .Y(
        c0sm_b0m_v0m_n125) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u264 ( .A0(c0sm_b0m_v0m_buffers0_1_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n125), 
        .Y(c0sm_b0m_v0m_n275) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u263 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n122), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n29), .C0(
        c0sm_b0m_v0m_n275), .Y(c0sm_headflit[1]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u262 ( .A(c0sm_headflit[1]), .Y(
        c0sm_b0m_v0m_n264) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u261 ( .A(reset), .Y(c0sm_b0m_v0m_n4) );
  AND4_X0P5M_A12TR c0sm_b0m_v0m_u260 ( .A(debitout_1), .B(c0sm_headflit[0]), 
        .C(c0sm_b0m_v0m_n264), .D(c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n1710) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u259 ( .A(c0sm_b0m_v0m_buffers2_10_), .Y(
        c0sm_b0m_v0m_n180) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u258 ( .A(c0sm_b0m_v0m_buffers3_10_), .Y(
        c0sm_b0m_v0m_n71) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u257 ( .A(c0sm_b0m_v0m_n353), .Y(
        c0sm_b0m_v0m_n183) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u256 ( .A0(c0sm_b0m_v0m_buffers0_10_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n183), 
        .Y(c0sm_b0m_v0m_n274) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u255 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n180), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n71), .C0(
        c0sm_b0m_v0m_n274), .Y(c0sm_b0m_headflit_10_) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u254 ( .A(c0sm_b0m_v0m_buffers2_11_), .Y(
        c0sm_b0m_v0m_n186) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u253 ( .A(c0sm_b0m_v0m_buffers3_11_), .Y(
        c0sm_b0m_v0m_n21) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u252 ( .A(c0sm_b0m_v0m_n354), .Y(
        c0sm_b0m_v0m_n190) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u251 ( .A0(c0sm_b0m_v0m_n193), .A1(
        c0sm_b0m_v0m_buffers0_11_), .B0(c0sm_b0m_v0m_n192), .B1(
        c0sm_b0m_v0m_n190), .Y(c0sm_b0m_v0m_n273) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u250 ( .A0(c0sm_b0m_v0m_n186), .A1(
        c0sm_b0m_v0m_n187), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n21), .C0(
        c0sm_b0m_v0m_n273), .Y(c0sm_b0m_headflit_11_) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u249 ( .A(c0sm_b0m_v0m_buffers2_2_), .Y(
        c0sm_b0m_v0m_n131) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u248 ( .A(c0sm_b0m_v0m_buffers3_2_), .Y(
        c0sm_b0m_v0m_n35) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u247 ( .A(c0sm_b0m_v0m_n345), .Y(
        c0sm_b0m_v0m_n134) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u246 ( .A0(c0sm_b0m_v0m_buffers0_2_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n134), 
        .Y(c0sm_b0m_v0m_n272) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u245 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n131), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n35), .C0(
        c0sm_b0m_v0m_n272), .Y(c0sm_headflit[2]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u244 ( .A(c0sm_b0m_v0m_buffers2_3_), .Y(
        c0sm_b0m_v0m_n138) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u243 ( .A(c0sm_b0m_v0m_buffers3_3_), .Y(
        c0sm_b0m_v0m_n38) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u242 ( .A(c0sm_b0m_v0m_n346), .Y(
        c0sm_b0m_v0m_n141) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u241 ( .A0(c0sm_b0m_v0m_buffers0_3_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n141), 
        .Y(c0sm_b0m_v0m_n271) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u240 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n138), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n38), .C0(
        c0sm_b0m_v0m_n271), .Y(c0sm_headflit[3]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u239 ( .A(c0sm_b0m_v0m_buffers2_4_), .Y(
        c0sm_b0m_v0m_n144) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u238 ( .A(c0sm_b0m_v0m_buffers3_4_), .Y(
        c0sm_b0m_v0m_n41) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u237 ( .A(c0sm_b0m_v0m_n347), .Y(
        c0sm_b0m_v0m_n147) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u236 ( .A0(c0sm_b0m_v0m_buffers0_4_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n147), 
        .Y(c0sm_b0m_v0m_n270) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u235 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n144), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n41), .C0(
        c0sm_b0m_v0m_n270), .Y(c0sm_headflit[4]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u234 ( .A(c0sm_b0m_v0m_buffers2_5_), .Y(
        c0sm_b0m_v0m_n150) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u233 ( .A(c0sm_b0m_v0m_buffers3_5_), .Y(
        c0sm_b0m_v0m_n44) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u232 ( .A(c0sm_b0m_v0m_n348), .Y(
        c0sm_b0m_v0m_n153) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u231 ( .A0(c0sm_b0m_v0m_buffers0_5_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n153), 
        .Y(c0sm_b0m_v0m_n269) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u230 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n150), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n44), .C0(
        c0sm_b0m_v0m_n269), .Y(c0sm_headflit[5]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u229 ( .A(c0sm_b0m_v0m_buffers2_6_), .Y(
        c0sm_b0m_v0m_n156) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u228 ( .A(c0sm_b0m_v0m_buffers3_6_), .Y(
        c0sm_b0m_v0m_n47) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u227 ( .A(c0sm_b0m_v0m_n349), .Y(
        c0sm_b0m_v0m_n159) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u226 ( .A0(c0sm_b0m_v0m_buffers0_6_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n159), 
        .Y(c0sm_b0m_v0m_n268) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u225 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n156), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n47), .C0(
        c0sm_b0m_v0m_n268), .Y(c0sm_headflit[6]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u224 ( .A(c0sm_b0m_v0m_buffers2_7_), .Y(
        c0sm_b0m_v0m_n162) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u223 ( .A(c0sm_b0m_v0m_buffers3_7_), .Y(
        c0sm_b0m_v0m_n62) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u222 ( .A(c0sm_b0m_v0m_n350), .Y(
        c0sm_b0m_v0m_n165) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u221 ( .A0(c0sm_b0m_v0m_buffers0_7_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n165), 
        .Y(c0sm_b0m_v0m_n267) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u220 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n162), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n62), .C0(
        c0sm_b0m_v0m_n267), .Y(c0sm_headflit[7]) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u219 ( .A(c0sm_b0m_v0m_buffers2_8_), .Y(
        c0sm_b0m_v0m_n168) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u218 ( .A(c0sm_b0m_v0m_buffers3_8_), .Y(
        c0sm_b0m_v0m_n65) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u217 ( .A(c0sm_b0m_v0m_n351), .Y(
        c0sm_b0m_v0m_n171) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u216 ( .A0(c0sm_b0m_v0m_buffers0_8_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n171), 
        .Y(c0sm_b0m_v0m_n266) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u215 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n168), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n65), .C0(
        c0sm_b0m_v0m_n266), .Y(c0sm_b0m_headflit_8_) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u214 ( .A(c0sm_b0m_v0m_buffers2_9_), .Y(
        c0sm_b0m_v0m_n174) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u213 ( .A(c0sm_b0m_v0m_buffers3_9_), .Y(
        c0sm_b0m_v0m_n68) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u212 ( .A(c0sm_b0m_v0m_n352), .Y(
        c0sm_b0m_v0m_n177) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u211 ( .A0(c0sm_b0m_v0m_buffers0_9_), .A1(
        c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n177), 
        .Y(c0sm_b0m_v0m_n265) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u210 ( .A0(c0sm_b0m_v0m_n187), .A1(
        c0sm_b0m_v0m_n174), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n68), .C0(
        c0sm_b0m_v0m_n265), .Y(c0sm_b0m_headflit_9_) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u209 ( .A(debitout_1), .B(reset), .Y(
        c0sm_b0m_v0m_n11) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u208 ( .A(c0sm_b0m_v0m_n11), .B(reset), .Y(
        c0sm_b0m_v0m_n10) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u207 ( .A0(c0sm_b0m_rdata[11]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_11_), 
        .Y(c0sm_b0m_v0m_n342) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u206 ( .A0(c0sm_b0m_rdata[10]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_10_), 
        .Y(c0sm_b0m_v0m_n341) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u205 ( .A0(c0sm_b0m_rdata[9]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_9_), 
        .Y(c0sm_b0m_v0m_n340) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u204 ( .A0(c0sm_b0m_rdata[8]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_8_), 
        .Y(c0sm_b0m_v0m_n339) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u203 ( .A0(c0sm_b0m_rdata[7]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[7]), .Y(
        c0sm_b0m_v0m_n338) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u202 ( .A0(c0sm_b0m_rdata[6]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[6]), .Y(
        c0sm_b0m_v0m_n337) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u201 ( .A0(c0sm_b0m_rdata[5]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[5]), .Y(
        c0sm_b0m_v0m_n336) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u200 ( .A0(c0sm_b0m_rdata[4]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[4]), .Y(
        c0sm_b0m_v0m_n335) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u199 ( .A0(c0sm_b0m_rdata[3]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[3]), .Y(
        c0sm_b0m_v0m_n334) );
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u198 ( .A0(c0sm_b0m_rdata[2]), .A1(
        c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[2]), .Y(
        c0sm_b0m_v0m_n333) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u197 ( .A(c0sm_b0m_v0m_n264), .B(
        c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n263) );
  MXT2_X0P5M_A12TR c0sm_b0m_v0m_u196 ( .A(c0sm_b0m_v0m_n263), .B(
        c0sm_b0m_rdata[1]), .S0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n332) );
  NAND2B_X0P5M_A12TR c0sm_b0m_v0m_u195 ( .AN(c0sm_headflit[0]), .B(
        c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n262) );
  MXT2_X0P5M_A12TR c0sm_b0m_v0m_u194 ( .A(c0sm_b0m_v0m_n262), .B(
        c0sm_b0m_rdata[0]), .S0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n331) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u193 ( .A(c0sm_b0m_v0m_tail_1_), .Y(
        c0sm_b0m_v0m_n7) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u192 ( .A(c0sm_b0m_v0m_tail_0_), .B(
        c0sm_b0m_v0m_n7), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n93) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u191 ( .A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_n2), 
        .Y(c0sm_b0m_v0m_n119) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u190 ( .A(c0sm_b0m_v0m_n119), .Y(
        c0sm_b0m_v0m_n135) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u189 ( .A(c0sm_b0m_v0m_tail_0_), .Y(
        c0sm_b0m_v0m_n3) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u188 ( .A(c0sm_b0m_v0m_tail_1_), .B(
        c0sm_b0m_v0m_n3), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n94) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u187 ( .A(c0sm_b0m_v0m_n94), .B(c0sm_b0m_n2), 
        .Y(c0sm_b0m_v0m_n121) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u186 ( .A(c0sm_b0m_v0m_n3), .B(
        c0sm_b0m_v0m_n7), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n95) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u185 ( .A(c0sm_b0m_v0m_n95), .B(c0sm_b0m_n2), 
        .Y(c0sm_b0m_v0m_n120) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u184 ( .A0(c0sm_b0m_v0m_buffers2_11_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_11_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n194) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u183 ( .A(c0sm_b0m_v0m_n95), .B(
        c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n93), .Y(c0sm_b0m_v0m_n28) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u182 ( .A(c0sm_b0m_v0m_n28), .B(c0sm_b0m_n2), 
        .Y(c0sm_b0m_v0m_n128) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u181 ( .A0(c0sm_b0m_v0m_buffers3_11_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_n2), .B1(c0sm_b0m_wdata_11_), .Y(
        c0sm_b0m_v0m_n195) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u180 ( .A0(c0sm_b0m_v0m_n354), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n194), .C0(c0sm_b0m_v0m_n195), 
        .Y(c0sm_b0m_v0m_n19) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u179 ( .A(c0sm_b0m_v0m_n94), .Y(
        c0sm_b0m_v0m_n108) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u178 ( .A(c0sm_b0m_v0m_n108), .B(
        c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n129) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u177 ( .A(c0sm_b0m_v0m_n193), .Y(
        c0sm_b0m_v0m_n96) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u176 ( .A(c0sm_b0m_v0m_n192), .Y(
        c0sm_b0m_v0m_n104) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u175 ( .A(debitout_1), .Y(c0sm_b0m_v0m_n191) );
  NAND4_X0P5A_A12TR c0sm_b0m_v0m_u174 ( .A(c0sm_b0m_v0m_n96), .B(
        c0sm_b0m_v0m_n104), .C(c0sm_b0m_v0m_n187), .D(c0sm_b0m_v0m_n191), .Y(
        c0sm_b0m_v0m_n111) );
  OR2_X0P5M_A12TR c0sm_b0m_v0m_u173 ( .A(c0sm_b0m_v0m_n187), .B(debitout_1), 
        .Y(c0sm_b0m_v0m_n110) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u172 ( .A(c0sm_b0m_v0m_n96), .B(debitout_1), 
        .Y(c0sm_b0m_v0m_n115) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u171 ( .A(c0sm_b0m_v0m_n104), .B(debitout_1), 
        .Y(c0sm_b0m_v0m_n113) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u170 ( .A0(c0sm_b0m_v0m_n115), .A1(
        c0sm_b0m_v0m_buffers0_11_), .B0(c0sm_b0m_v0m_n113), .B1(
        c0sm_b0m_v0m_n190), .Y(c0sm_b0m_v0m_n189) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u169 ( .A0(c0sm_b0m_v0m_n21), .A1(
        c0sm_b0m_v0m_n111), .B0(c0sm_b0m_v0m_n186), .B1(c0sm_b0m_v0m_n110), 
        .C0(c0sm_b0m_v0m_n189), .Y(c0sm_b0m_v0m_n188) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u168 ( .A(c0sm_b0m_v0m_n188), .Y(
        c0sm_b0m_v0m_n17) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u167 ( .A(c0sm_b0m_v0m_n187), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n94), .Y(c0sm_b0m_v0m_n107) );
  OAI21_X0P5M_A12TR c0sm_b0m_v0m_u166 ( .A0(c0sm_b0m_v0m_n3), .A1(
        c0sm_b0m_v0m_n7), .B0(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n26) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u165 ( .A(c0sm_b0m_v0m_n26), .Y(
        c0sm_b0m_v0m_n72) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u164 ( .A(c0sm_b0m_v0m_n93), .B(
        c0sm_b0m_v0m_n95), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n109) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u163 ( .A(c0sm_b0m_v0m_n107), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n109), .Y(c0sm_b0m_v0m_n130) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u162 ( .A0(c0sm_b0m_v0m_n19), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n186), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n330)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u161 ( .A0(c0sm_b0m_v0m_buffers2_10_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_10_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n184) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u160 ( .A0(c0sm_b0m_v0m_buffers3_10_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_10_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n185) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u159 ( .A0(c0sm_b0m_v0m_n353), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n184), .C0(c0sm_b0m_v0m_n185), 
        .Y(c0sm_b0m_v0m_n70) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u158 ( .A0(c0sm_b0m_v0m_buffers0_10_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n183), 
        .Y(c0sm_b0m_v0m_n182) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u157 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n71), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n180), 
        .C0(c0sm_b0m_v0m_n182), .Y(c0sm_b0m_v0m_n181) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u156 ( .A(c0sm_b0m_v0m_n181), .Y(
        c0sm_b0m_v0m_n69) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u155 ( .A0(c0sm_b0m_v0m_n70), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n180), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n329)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u154 ( .A0(c0sm_b0m_v0m_buffers2_9_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_9_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n178) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u153 ( .A0(c0sm_b0m_v0m_buffers3_9_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_9_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n179) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u152 ( .A0(c0sm_b0m_v0m_n352), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n178), .C0(c0sm_b0m_v0m_n179), 
        .Y(c0sm_b0m_v0m_n67) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u151 ( .A0(c0sm_b0m_v0m_buffers0_9_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n177), 
        .Y(c0sm_b0m_v0m_n176) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u150 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n68), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n174), 
        .C0(c0sm_b0m_v0m_n176), .Y(c0sm_b0m_v0m_n175) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u149 ( .A(c0sm_b0m_v0m_n175), .Y(
        c0sm_b0m_v0m_n66) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u148 ( .A0(c0sm_b0m_v0m_n67), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n174), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n328)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u147 ( .A0(c0sm_b0m_v0m_buffers2_8_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_8_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n172) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u146 ( .A0(c0sm_b0m_v0m_buffers3_8_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_8_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n173) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u145 ( .A0(c0sm_b0m_v0m_n351), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n172), .C0(c0sm_b0m_v0m_n173), 
        .Y(c0sm_b0m_v0m_n64) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u144 ( .A0(c0sm_b0m_v0m_buffers0_8_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n171), 
        .Y(c0sm_b0m_v0m_n170) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u143 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n65), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n168), 
        .C0(c0sm_b0m_v0m_n170), .Y(c0sm_b0m_v0m_n169) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u142 ( .A(c0sm_b0m_v0m_n169), .Y(
        c0sm_b0m_v0m_n63) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u141 ( .A0(c0sm_b0m_v0m_n64), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n168), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n327)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u140 ( .A0(c0sm_b0m_v0m_buffers2_7_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_7_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n166) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u139 ( .A0(c0sm_b0m_v0m_buffers3_7_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_7_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n167) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u138 ( .A0(c0sm_b0m_v0m_n350), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n166), .C0(c0sm_b0m_v0m_n167), 
        .Y(c0sm_b0m_v0m_n49) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u137 ( .A0(c0sm_b0m_v0m_buffers0_7_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n165), 
        .Y(c0sm_b0m_v0m_n164) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u136 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n62), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n162), 
        .C0(c0sm_b0m_v0m_n164), .Y(c0sm_b0m_v0m_n163) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u135 ( .A(c0sm_b0m_v0m_n163), .Y(
        c0sm_b0m_v0m_n48) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u134 ( .A0(c0sm_b0m_v0m_n49), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n162), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n326)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u133 ( .A0(c0sm_b0m_v0m_buffers2_6_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_6_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n160) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u132 ( .A0(c0sm_b0m_v0m_buffers3_6_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_6_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n161) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u131 ( .A0(c0sm_b0m_v0m_n349), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n160), .C0(c0sm_b0m_v0m_n161), 
        .Y(c0sm_b0m_v0m_n46) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u130 ( .A0(c0sm_b0m_v0m_buffers0_6_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n159), 
        .Y(c0sm_b0m_v0m_n158) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u129 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n47), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n156), 
        .C0(c0sm_b0m_v0m_n158), .Y(c0sm_b0m_v0m_n157) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u128 ( .A(c0sm_b0m_v0m_n157), .Y(
        c0sm_b0m_v0m_n45) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u127 ( .A0(c0sm_b0m_v0m_n46), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n156), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n325)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u126 ( .A0(c0sm_b0m_v0m_buffers2_5_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_5_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n154) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u125 ( .A0(c0sm_b0m_v0m_buffers3_5_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_5_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n155) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u124 ( .A0(c0sm_b0m_v0m_n348), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n154), .C0(c0sm_b0m_v0m_n155), 
        .Y(c0sm_b0m_v0m_n43) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u123 ( .A0(c0sm_b0m_v0m_buffers0_5_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n153), 
        .Y(c0sm_b0m_v0m_n152) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u122 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n44), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n150), 
        .C0(c0sm_b0m_v0m_n152), .Y(c0sm_b0m_v0m_n151) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u121 ( .A(c0sm_b0m_v0m_n151), .Y(
        c0sm_b0m_v0m_n42) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u120 ( .A0(c0sm_b0m_v0m_n43), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n150), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n324)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u119 ( .A0(c0sm_b0m_v0m_buffers2_4_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_4_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n148) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u118 ( .A0(c0sm_b0m_v0m_buffers3_4_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_4_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n149) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u117 ( .A0(c0sm_b0m_v0m_n347), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n148), .C0(c0sm_b0m_v0m_n149), 
        .Y(c0sm_b0m_v0m_n40) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u116 ( .A0(c0sm_b0m_v0m_buffers0_4_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n147), 
        .Y(c0sm_b0m_v0m_n146) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u115 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n41), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n144), 
        .C0(c0sm_b0m_v0m_n146), .Y(c0sm_b0m_v0m_n145) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u114 ( .A(c0sm_b0m_v0m_n145), .Y(
        c0sm_b0m_v0m_n39) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u113 ( .A0(c0sm_b0m_v0m_n40), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n144), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n323)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u112 ( .A0(c0sm_b0m_v0m_buffers2_3_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_3_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n142) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u111 ( .A0(c0sm_b0m_v0m_buffers3_3_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_3_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n143) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u110 ( .A0(c0sm_b0m_v0m_n346), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n142), .C0(c0sm_b0m_v0m_n143), 
        .Y(c0sm_b0m_v0m_n37) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u109 ( .A0(c0sm_b0m_v0m_buffers0_3_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n141), 
        .Y(c0sm_b0m_v0m_n140) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u108 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n38), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n138), 
        .C0(c0sm_b0m_v0m_n140), .Y(c0sm_b0m_v0m_n139) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u107 ( .A(c0sm_b0m_v0m_n139), .Y(
        c0sm_b0m_v0m_n36) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u106 ( .A0(c0sm_b0m_v0m_n37), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n138), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n322)
         );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u105 ( .A0(c0sm_b0m_v0m_buffers2_2_), .A1(
        c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_2_), .B1(
        c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n136) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u104 ( .A0(c0sm_b0m_v0m_buffers3_2_), .A1(
        c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_2_), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n137) );
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u103 ( .A0(c0sm_b0m_v0m_n345), .A1(
        c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n136), .C0(c0sm_b0m_v0m_n137), 
        .Y(c0sm_b0m_v0m_n34) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u102 ( .A0(c0sm_b0m_v0m_buffers0_2_), .A1(
        c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n134), 
        .Y(c0sm_b0m_v0m_n133) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u101 ( .A0(c0sm_b0m_v0m_n111), .A1(
        c0sm_b0m_v0m_n35), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n131), 
        .C0(c0sm_b0m_v0m_n133), .Y(c0sm_b0m_v0m_n132) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u100 ( .A(c0sm_b0m_v0m_n132), .Y(
        c0sm_b0m_v0m_n33) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u99 ( .A0(c0sm_b0m_v0m_n34), .A1(
        c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n130), 
        .C0(c0sm_b0m_v0m_n131), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n321)
         );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u98 ( .A(c0sm_b0m_v0m_n128), .Y(
        c0sm_b0m_v0m_n116) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u97 ( .A0(c0sm_b0m_v0m_buffers0_1_), .A1(
        c0sm_b0m_v0m_n120), .B0(c0sm_b0m_v0m_buffers2_1_), .B1(
        c0sm_b0m_v0m_n121), .Y(c0sm_b0m_v0m_n126) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u96 ( .A0(c0sm_b0m_v0m_n119), .A1(
        c0sm_b0m_v0m_n125), .B0(flitin_1[1]), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n127) );
  OAI211_X0P5M_A12TR c0sm_b0m_v0m_u95 ( .A0(c0sm_b0m_v0m_n116), .A1(
        c0sm_b0m_v0m_n29), .B0(c0sm_b0m_v0m_n126), .C0(c0sm_b0m_v0m_n127), .Y(
        c0sm_b0m_v0m_n31) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u94 ( .A0(c0sm_b0m_v0m_n113), .A1(
        c0sm_b0m_v0m_n125), .B0(c0sm_b0m_v0m_buffers0_1_), .B1(
        c0sm_b0m_v0m_n115), .C0(debitout_1), .Y(c0sm_b0m_v0m_n124) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u93 ( .A0(c0sm_b0m_v0m_n110), .A1(
        c0sm_b0m_v0m_n122), .B0(c0sm_b0m_v0m_n111), .B1(c0sm_b0m_v0m_n29), 
        .C0(c0sm_b0m_v0m_n124), .Y(c0sm_b0m_v0m_n32) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u92 ( .A0(c0sm_b0m_v0m_n108), .A1(
        c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n109), .B1(c0sm_b0m_v0m_n32), .C0(
        reset), .Y(c0sm_b0m_v0m_n123) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u91 ( .A(c0sm_b0m_v0m_n122), .B(
        c0sm_b0m_v0m_n123), .S0(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n320) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u90 ( .A0(c0sm_b0m_v0m_buffers0_0_), .A1(
        c0sm_b0m_v0m_n120), .B0(c0sm_b0m_v0m_buffers2_0_), .B1(
        c0sm_b0m_v0m_n121), .Y(c0sm_b0m_v0m_n117) );
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u89 ( .A0(c0sm_b0m_v0m_n119), .A1(
        c0sm_b0m_v0m_n114), .B0(flitin_1[0]), .B1(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n118) );
  OAI211_X0P5M_A12TR c0sm_b0m_v0m_u88 ( .A0(c0sm_b0m_v0m_n116), .A1(
        c0sm_b0m_v0m_n23), .B0(c0sm_b0m_v0m_n117), .C0(c0sm_b0m_v0m_n118), .Y(
        c0sm_b0m_v0m_n25) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u87 ( .A0(c0sm_b0m_v0m_n113), .A1(
        c0sm_b0m_v0m_n114), .B0(c0sm_b0m_v0m_buffers0_0_), .B1(
        c0sm_b0m_v0m_n115), .C0(debitout_1), .Y(c0sm_b0m_v0m_n112) );
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u86 ( .A0(c0sm_b0m_v0m_n110), .A1(
        c0sm_b0m_v0m_n105), .B0(c0sm_b0m_v0m_n111), .B1(c0sm_b0m_v0m_n23), 
        .C0(c0sm_b0m_v0m_n112), .Y(c0sm_b0m_v0m_n27) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u85 ( .A0(c0sm_b0m_v0m_n108), .A1(
        c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n109), .B1(c0sm_b0m_v0m_n27), .C0(
        reset), .Y(c0sm_b0m_v0m_n106) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u84 ( .A(c0sm_b0m_v0m_n105), .B(
        c0sm_b0m_v0m_n106), .S0(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n319) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u83 ( .A(c0sm_b0m_v0m_n93), .Y(c0sm_b0m_v0m_n99) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u82 ( .A(c0sm_b0m_v0m_n99), .B(
        c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n102) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u81 ( .A(c0sm_b0m_v0m_n93), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n104), .Y(c0sm_b0m_v0m_n98) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u80 ( .A(c0sm_b0m_v0m_n95), .B(
        c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n100) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u79 ( .A(c0sm_b0m_v0m_n98), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n100), .Y(c0sm_b0m_v0m_n103) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u78 ( .A0(c0sm_b0m_v0m_n19), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n354), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n318)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u77 ( .A0(c0sm_b0m_v0m_n70), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n353), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n317)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u76 ( .A0(c0sm_b0m_v0m_n67), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n352), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n316)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u75 ( .A0(c0sm_b0m_v0m_n64), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n351), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n315)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u74 ( .A0(c0sm_b0m_v0m_n49), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n350), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n314)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u73 ( .A0(c0sm_b0m_v0m_n46), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n349), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n313)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u72 ( .A0(c0sm_b0m_v0m_n43), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n348), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n312)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u71 ( .A0(c0sm_b0m_v0m_n40), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n347), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n311)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u70 ( .A0(c0sm_b0m_v0m_n37), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n346), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n310)
         );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u69 ( .A0(c0sm_b0m_v0m_n34), .A1(
        c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n103), 
        .C0(c0sm_b0m_v0m_n345), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n309)
         );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u68 ( .A0(c0sm_b0m_v0m_n99), .A1(
        c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n100), .B1(c0sm_b0m_v0m_n32), .C0(
        reset), .Y(c0sm_b0m_v0m_n101) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u67 ( .A(c0sm_b0m_v0m_n344), .B(
        c0sm_b0m_v0m_n101), .S0(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n308) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u66 ( .A0(c0sm_b0m_v0m_n99), .A1(
        c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n100), .B1(c0sm_b0m_v0m_n27), .C0(
        reset), .Y(c0sm_b0m_v0m_n97) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u65 ( .A(c0sm_b0m_v0m_n343), .B(
        c0sm_b0m_v0m_n97), .S0(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n307) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u64 ( .A(c0sm_b0m_v0m_n95), .Y(c0sm_b0m_v0m_n77) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u63 ( .A(c0sm_b0m_v0m_n77), .B(
        c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n81) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u62 ( .A(c0sm_b0m_v0m_n95), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n96), .Y(c0sm_b0m_v0m_n76) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u61 ( .A(c0sm_b0m_v0m_n93), .B(
        c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n78) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u60 ( .A(c0sm_b0m_v0m_n76), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n78), .Y(c0sm_b0m_v0m_n82) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u59 ( .A(c0sm_b0m_v0m_buffers0_11_), .Y(
        c0sm_b0m_v0m_n92) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u58 ( .A0(c0sm_b0m_v0m_n19), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n92), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n306) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u57 ( .A(c0sm_b0m_v0m_buffers0_10_), .Y(
        c0sm_b0m_v0m_n91) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u56 ( .A0(c0sm_b0m_v0m_n70), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n91), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n305) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u55 ( .A(c0sm_b0m_v0m_buffers0_9_), .Y(
        c0sm_b0m_v0m_n90) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u54 ( .A0(c0sm_b0m_v0m_n67), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n90), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n304) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u53 ( .A(c0sm_b0m_v0m_buffers0_8_), .Y(
        c0sm_b0m_v0m_n89) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u52 ( .A0(c0sm_b0m_v0m_n64), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n89), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n303) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u51 ( .A(c0sm_b0m_v0m_buffers0_7_), .Y(
        c0sm_b0m_v0m_n88) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u50 ( .A0(c0sm_b0m_v0m_n49), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n88), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n302) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u49 ( .A(c0sm_b0m_v0m_buffers0_6_), .Y(
        c0sm_b0m_v0m_n87) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u48 ( .A0(c0sm_b0m_v0m_n46), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n87), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n301) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u47 ( .A(c0sm_b0m_v0m_buffers0_5_), .Y(
        c0sm_b0m_v0m_n86) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u46 ( .A0(c0sm_b0m_v0m_n43), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n86), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n300) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u45 ( .A(c0sm_b0m_v0m_buffers0_4_), .Y(
        c0sm_b0m_v0m_n85) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u44 ( .A0(c0sm_b0m_v0m_n40), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n85), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n299) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u43 ( .A(c0sm_b0m_v0m_buffers0_3_), .Y(
        c0sm_b0m_v0m_n84) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u42 ( .A0(c0sm_b0m_v0m_n37), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n84), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n298) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u41 ( .A(c0sm_b0m_v0m_buffers0_2_), .Y(
        c0sm_b0m_v0m_n83) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u40 ( .A0(c0sm_b0m_v0m_n34), .A1(
        c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n82), .C0(
        c0sm_b0m_v0m_n83), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n297) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u39 ( .A(c0sm_b0m_v0m_buffers0_1_), .Y(
        c0sm_b0m_v0m_n79) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u38 ( .A0(c0sm_b0m_v0m_n77), .A1(
        c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n78), .B1(c0sm_b0m_v0m_n32), .C0(
        reset), .Y(c0sm_b0m_v0m_n80) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u37 ( .A(c0sm_b0m_v0m_n79), .B(
        c0sm_b0m_v0m_n80), .S0(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n296) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u36 ( .A(c0sm_b0m_v0m_buffers0_0_), .Y(
        c0sm_b0m_v0m_n74) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u35 ( .A0(c0sm_b0m_v0m_n77), .A1(
        c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n78), .B1(c0sm_b0m_v0m_n27), .C0(
        reset), .Y(c0sm_b0m_v0m_n75) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u34 ( .A(c0sm_b0m_v0m_n74), .B(
        c0sm_b0m_v0m_n75), .S0(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n295) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u33 ( .A(c0sm_b0m_v0m_n72), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n73), .Y(c0sm_b0m_v0m_n22) );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u32 ( .A(c0sm_b0m_v0m_n22), .B(
        c0sm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n28), .Y(c0sm_b0m_v0m_n18) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u31 ( .A(c0sm_b0m_v0m_n26), .B(
        c0sm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n20) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u30 ( .A0(c0sm_b0m_v0m_n69), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n70), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n71), .Y(c0sm_b0m_v0m_n294) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u29 ( .A0(c0sm_b0m_v0m_n66), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n67), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n68), .Y(c0sm_b0m_v0m_n293) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u28 ( .A0(c0sm_b0m_v0m_n63), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n64), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n65), .Y(c0sm_b0m_v0m_n292) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u27 ( .A0(c0sm_b0m_v0m_n48), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n49), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n62), .Y(c0sm_b0m_v0m_n291) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u26 ( .A0(c0sm_b0m_v0m_n45), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n46), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n47), .Y(c0sm_b0m_v0m_n290) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u25 ( .A0(c0sm_b0m_v0m_n42), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n43), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n44), .Y(c0sm_b0m_v0m_n289) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u24 ( .A0(c0sm_b0m_v0m_n39), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n40), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n41), .Y(c0sm_b0m_v0m_n288) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u23 ( .A0(c0sm_b0m_v0m_n36), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n37), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n38), .Y(c0sm_b0m_v0m_n287) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u22 ( .A0(c0sm_b0m_v0m_n33), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n34), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n35), .Y(c0sm_b0m_v0m_n286) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u21 ( .A0(c0sm_b0m_v0m_n31), .A1(
        c0sm_b0m_v0m_n26), .B0(c0sm_b0m_v0m_n32), .B1(c0sm_b0m_v0m_n28), .C0(
        reset), .Y(c0sm_b0m_v0m_n30) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u20 ( .A(c0sm_b0m_v0m_n29), .B(
        c0sm_b0m_v0m_n30), .S0(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n285) );
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u19 ( .A0(c0sm_b0m_v0m_n25), .A1(
        c0sm_b0m_v0m_n26), .B0(c0sm_b0m_v0m_n27), .B1(c0sm_b0m_v0m_n28), .C0(
        reset), .Y(c0sm_b0m_v0m_n24) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u18 ( .A(c0sm_b0m_v0m_n23), .B(
        c0sm_b0m_v0m_n24), .S0(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n284) );
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u17 ( .A0(c0sm_b0m_v0m_n17), .A1(
        c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n19), .B1(c0sm_b0m_v0m_n20), .C0(
        c0sm_b0m_v0m_n21), .C1(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n283) );
  AOI21_X0P5M_A12TR c0sm_b0m_v0m_u16 ( .A0(c0sm_b0m_v0m_n4), .A1(
        c0sm_b0m_v0m_n16), .B0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n12) );
  OA21A1OI2_X0P5M_A12TR c0sm_b0m_v0m_u15 ( .A0(reset), .A1(
        c0sm_b0m_v0m_head_1_), .B0(c0sm_b0m_v0m_n12), .C0(c0sm_b0m_v0m_n15), 
        .Y(c0sm_b0m_v0m_n282) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u14 ( .A(c0sm_b0m_v0m_n10), .B(
        c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n13) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u13 ( .A(c0sm_b0m_v0m_head_1_), .Y(
        c0sm_b0m_v0m_n14) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u12 ( .A(c0sm_b0m_v0m_n12), .B(
        c0sm_b0m_v0m_n13), .S0(c0sm_b0m_v0m_n14), .Y(c0sm_b0m_v0m_n281) );
  MXT2_X0P5M_A12TR c0sm_b0m_v0m_u11 ( .A(c0sm_b0m_v0m_n10), .B(
        c0sm_b0m_v0m_n11), .S0(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n280) );
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u10 ( .A(reset), .B(c0sm_b0m_n2), .Y(
        c0sm_b0m_v0m_n8) );
  AOI21_X0P5M_A12TR c0sm_b0m_v0m_u9 ( .A0(c0sm_b0m_v0m_n3), .A1(
        c0sm_b0m_v0m_n4), .B0(c0sm_b0m_v0m_n8), .Y(c0sm_b0m_v0m_n5) );
  OA21A1OI2_X0P5M_A12TR c0sm_b0m_v0m_u8 ( .A0(c0sm_b0m_v0m_tail_1_), .A1(reset), .B0(c0sm_b0m_v0m_n5), .C0(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n279) );
  INV_X0P5B_A12TR c0sm_b0m_v0m_u7 ( .A(c0sm_b0m_v0m_n8), .Y(c0sm_b0m_v0m_n1)
         );
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u6 ( .A(c0sm_b0m_v0m_n1), .B(c0sm_b0m_v0m_n4), 
        .C(c0sm_b0m_v0m_tail_0_), .Y(c0sm_b0m_v0m_n6) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u5 ( .A(c0sm_b0m_v0m_n5), .B(c0sm_b0m_v0m_n6), 
        .S0(c0sm_b0m_v0m_n7), .Y(c0sm_b0m_v0m_n278) );
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u4 ( .A(c0sm_b0m_v0m_n1), .B(c0sm_b0m_v0m_n4), 
        .Y(c0sm_b0m_v0m_n2) );
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u3 ( .A(c0sm_b0m_v0m_n1), .B(c0sm_b0m_v0m_n2), 
        .S0(c0sm_b0m_v0m_n3), .Y(c0sm_b0m_v0m_n277) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_tail_reg_2_ ( .D(c0sm_b0m_v0m_n279), .CK(clk), 
        .QN(c0sm_b0m_v0m_n355) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_2_ ( .D(c0sm_b0m_v0m_n309), .CK(
        clk), .QN(c0sm_b0m_v0m_n345) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_3_ ( .D(c0sm_b0m_v0m_n310), .CK(
        clk), .QN(c0sm_b0m_v0m_n346) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_4_ ( .D(c0sm_b0m_v0m_n311), .CK(
        clk), .QN(c0sm_b0m_v0m_n347) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_5_ ( .D(c0sm_b0m_v0m_n312), .CK(
        clk), .QN(c0sm_b0m_v0m_n348) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_6_ ( .D(c0sm_b0m_v0m_n313), .CK(
        clk), .QN(c0sm_b0m_v0m_n349) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_7_ ( .D(c0sm_b0m_v0m_n314), .CK(
        clk), .QN(c0sm_b0m_v0m_n350) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_8_ ( .D(c0sm_b0m_v0m_n315), .CK(
        clk), .QN(c0sm_b0m_v0m_n351) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_9_ ( .D(c0sm_b0m_v0m_n316), .CK(
        clk), .QN(c0sm_b0m_v0m_n352) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_10_ ( .D(c0sm_b0m_v0m_n317), .CK(
        clk), .QN(c0sm_b0m_v0m_n353) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_11_ ( .D(c0sm_b0m_v0m_n318), .CK(
        clk), .QN(c0sm_b0m_v0m_n354) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_0_ ( .D(c0sm_b0m_v0m_n307), .CK(
        clk), .QN(c0sm_b0m_v0m_n343) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_1_ ( .D(c0sm_b0m_v0m_n308), .CK(
        clk), .QN(c0sm_b0m_v0m_n344) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_1_ ( .D(c0sm_b0m_v0m_n281), .CK(clk), 
        .Q(c0sm_b0m_v0m_head_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_0_ ( .D(c0sm_b0m_v0m_n280), .CK(clk), 
        .Q(c0sm_b0m_v0m_head_0_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_tailout_reg ( .D(c0sm_b0m_v0m_n1710), .CK(clk), 
        .Q(tailout_1) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_11_ ( .D(c0sm_b0m_v0m_n306), .CK(
        clk), .Q(c0sm_b0m_v0m_buffers0_11_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_0_ ( .D(c0sm_b0m_v0m_n295), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_0_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_1_ ( .D(c0sm_b0m_v0m_n296), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_2_ ( .D(c0sm_b0m_v0m_n297), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_2_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_3_ ( .D(c0sm_b0m_v0m_n298), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_3_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_4_ ( .D(c0sm_b0m_v0m_n299), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_4_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_5_ ( .D(c0sm_b0m_v0m_n300), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_5_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_6_ ( .D(c0sm_b0m_v0m_n301), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_6_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_7_ ( .D(c0sm_b0m_v0m_n302), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_7_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_8_ ( .D(c0sm_b0m_v0m_n303), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_8_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_9_ ( .D(c0sm_b0m_v0m_n304), .CK(clk), .Q(c0sm_b0m_v0m_buffers0_9_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_10_ ( .D(c0sm_b0m_v0m_n305), .CK(
        clk), .Q(c0sm_b0m_v0m_buffers0_10_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_2_ ( .D(c0sm_b0m_v0m_n282), .CK(clk), 
        .Q(c0sm_b0m_v0m_head_2_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_tail_reg_0_ ( .D(c0sm_b0m_v0m_n277), .CK(clk), 
        .Q(c0sm_b0m_v0m_tail_0_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_tail_reg_1_ ( .D(c0sm_b0m_v0m_n278), .CK(clk), 
        .Q(c0sm_b0m_v0m_tail_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_2_ ( .D(c0sm_b0m_v0m_n321), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_2_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_2_ ( .D(c0sm_b0m_v0m_n286), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_2_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_3_ ( .D(c0sm_b0m_v0m_n322), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_3_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_3_ ( .D(c0sm_b0m_v0m_n287), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_3_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_4_ ( .D(c0sm_b0m_v0m_n323), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_4_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_4_ ( .D(c0sm_b0m_v0m_n288), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_4_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_5_ ( .D(c0sm_b0m_v0m_n324), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_5_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_5_ ( .D(c0sm_b0m_v0m_n289), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_5_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_6_ ( .D(c0sm_b0m_v0m_n325), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_6_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_6_ ( .D(c0sm_b0m_v0m_n290), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_6_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_7_ ( .D(c0sm_b0m_v0m_n326), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_7_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_7_ ( .D(c0sm_b0m_v0m_n291), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_7_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_8_ ( .D(c0sm_b0m_v0m_n327), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_8_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_8_ ( .D(c0sm_b0m_v0m_n292), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_8_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_9_ ( .D(c0sm_b0m_v0m_n328), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_9_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_9_ ( .D(c0sm_b0m_v0m_n293), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_9_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_10_ ( .D(c0sm_b0m_v0m_n329), .CK(
        clk), .Q(c0sm_b0m_v0m_buffers2_10_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_10_ ( .D(c0sm_b0m_v0m_n294), .CK(
        clk), .Q(c0sm_b0m_v0m_buffers3_10_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_11_ ( .D(c0sm_b0m_v0m_n330), .CK(
        clk), .Q(c0sm_b0m_v0m_buffers2_11_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_11_ ( .D(c0sm_b0m_v0m_n283), .CK(
        clk), .Q(c0sm_b0m_v0m_buffers3_11_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_0_ ( .D(c0sm_b0m_v0m_n319), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_0_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_1_ ( .D(c0sm_b0m_v0m_n320), .CK(clk), .Q(c0sm_b0m_v0m_buffers2_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_0_ ( .D(c0sm_b0m_v0m_n331), .CK(clk), 
        .Q(c0sm_b0m_rdata[0]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_1_ ( .D(c0sm_b0m_v0m_n332), .CK(clk), 
        .Q(c0sm_b0m_rdata[1]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_10_ ( .D(c0sm_b0m_v0m_n341), .CK(clk), 
        .Q(c0sm_b0m_rdata[10]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_11_ ( .D(c0sm_b0m_v0m_n342), .CK(clk), 
        .Q(c0sm_b0m_rdata[11]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_2_ ( .D(c0sm_b0m_v0m_n333), .CK(clk), 
        .Q(c0sm_b0m_rdata[2]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_3_ ( .D(c0sm_b0m_v0m_n334), .CK(clk), 
        .Q(c0sm_b0m_rdata[3]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_4_ ( .D(c0sm_b0m_v0m_n335), .CK(clk), 
        .Q(c0sm_b0m_rdata[4]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_5_ ( .D(c0sm_b0m_v0m_n336), .CK(clk), 
        .Q(c0sm_b0m_rdata[5]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_6_ ( .D(c0sm_b0m_v0m_n337), .CK(clk), 
        .Q(c0sm_b0m_rdata[6]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_7_ ( .D(c0sm_b0m_v0m_n338), .CK(clk), 
        .Q(c0sm_b0m_rdata[7]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_8_ ( .D(c0sm_b0m_v0m_n339), .CK(clk), 
        .Q(c0sm_b0m_rdata[8]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_9_ ( .D(c0sm_b0m_v0m_n340), .CK(clk), 
        .Q(c0sm_b0m_rdata[9]) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_0_ ( .D(c0sm_b0m_v0m_n284), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_0_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_1_ ( .D(c0sm_b0m_v0m_n285), .CK(clk), .Q(c0sm_b0m_v0m_buffers3_1_) );
  INV_X0P5B_A12TR c0sm_r0m_u20 ( .A(currx[2]), .Y(c0sm_r0m_n4) );
  INV_X0P5B_A12TR c0sm_r0m_u19 ( .A(c0sm_headflit[5]), .Y(c0sm_r0m_n9) );
  OR2_X0P5M_A12TR c0sm_r0m_u18 ( .A(currx[0]), .B(c0sm_r0m_n9), .Y(
        c0sm_r0m_n15) );
  INV_X0P5B_A12TR c0sm_r0m_u17 ( .A(c0sm_headflit[6]), .Y(c0sm_r0m_n8) );
  AND2_X0P5M_A12TR c0sm_r0m_u16 ( .A(c0sm_r0m_n15), .B(currx[1]), .Y(
        c0sm_r0m_n16) );
  OA21A1OI2_X0P5M_A12TR c0sm_r0m_u15 ( .A0(currx[1]), .A1(c0sm_r0m_n15), .B0(
        c0sm_r0m_n8), .C0(c0sm_r0m_n16), .Y(c0sm_r0m_n6) );
  AOI2XB1_X0P5M_A12TR c0sm_r0m_u14 ( .A1N(curry[1]), .A0(c0sm_headflit[3]), 
        .B0(c0sm_headflit[2]), .Y(c0sm_r0m_n13) );
  INV_X0P5B_A12TR c0sm_r0m_u13 ( .A(c0sm_headflit[3]), .Y(c0sm_r0m_n14) );
  AOI22_X0P5M_A12TR c0sm_r0m_u12 ( .A0(c0sm_r0m_n13), .A1(curry[0]), .B0(
        curry[1]), .B1(c0sm_r0m_n14), .Y(c0sm_r0m_n12) );
  AOI2XB1_X0P5M_A12TR c0sm_r0m_u11 ( .A1N(curry[2]), .A0(c0sm_headflit[4]), 
        .B0(c0sm_r0m_n12), .Y(c0sm_r0m_n11) );
  AOI2XB1_X0P5M_A12TR c0sm_r0m_u10 ( .A1N(c0sm_headflit[4]), .A0(curry[2]), 
        .B0(c0sm_r0m_n11), .Y(c0sm_r0m_n10) );
  AOI221_X0P5M_A12TR c0sm_r0m_u9 ( .A0(currx[1]), .A1(c0sm_r0m_n8), .B0(
        currx[0]), .B1(c0sm_r0m_n9), .C0(c0sm_r0m_n10), .Y(c0sm_r0m_n7) );
  OAI22_X0P5M_A12TR c0sm_r0m_u8 ( .A0(c0sm_r0m_n6), .A1(c0sm_r0m_n7), .B0(
        c0sm_headflit[7]), .B1(c0sm_r0m_n4), .Y(c0sm_r0m_n5) );
  AO1B2_X0P5M_A12TR c0sm_r0m_u7 ( .B0(c0sm_r0m_n4), .B1(c0sm_headflit[7]), 
        .A0N(c0sm_r0m_n5), .Y(c0sm_r0m_n3) );
  INV_X0P5B_A12TR c0sm_r0m_u6 ( .A(c0sm_n4), .Y(c0sm_r0m_n1) );
  NOR3_X0P5A_A12TR c0sm_r0m_u5 ( .A(c0sm_r0m_n3), .B(reset), .C(c0sm_r0m_n1), 
        .Y(c0sm_r0m_n100) );
  INV_X0P5B_A12TR c0sm_r0m_u4 ( .A(c0sm_r0m_n3), .Y(c0sm_r0m_n2) );
  NOR3_X0P5A_A12TR c0sm_r0m_u3 ( .A(c0sm_r0m_n1), .B(reset), .C(c0sm_r0m_n2), 
        .Y(c0sm_r0m_n110) );
  DFFQ_X1M_A12TR c0sm_r0m_vc_req_reg_0_ ( .D(c0sm_r0m_n100), .CK(clk), .Q(
        c0sm_routewire[0]) );
  DFFQ_X1M_A12TR c0sm_r0m_vc_req_reg_1_ ( .D(c0sm_r0m_n110), .CK(clk), .Q(
        c0sm_routewire[1]) );
  INV_X0P5B_A12TR c0sm_v0m_u40 ( .A(c0sm_v0m_state_status_1_), .Y(c0sm_v0m_n29) );
  OAI211_X0P5M_A12TR c0sm_v0m_u39 ( .A0(swalloc_resp_1[1]), .A1(
        swalloc_resp_1[0]), .B0(c0sm_v0m_n29), .C0(c0sm_v0m_state_status_0_), 
        .Y(c0sm_v0m_n5) );
  NOR2_X0P5A_A12TR c0sm_v0m_u38 ( .A(reset), .B(tailout_1), .Y(c0sm_v0m_n8) );
  AO1B2_X0P5M_A12TR c0sm_v0m_u37 ( .B0(c0sm_v0m_n5), .B1(
        c0sm_v0m_state_status_0_), .A0N(c0sm_v0m_n8), .Y(c0sm_v0m_n57) );
  OA211_X0P5M_A12TR c0sm_v0m_u36 ( .A0(c0sm_routewire[1]), .A1(
        c0sm_routewire[0]), .B0(c0sm_v0m_state_status_0_), .C0(
        c0sm_v0m_state_status_1_), .Y(c0sm_v0m_n4) );
  AO21A1AI2_X0P5M_A12TR c0sm_v0m_u35 ( .A0(c0sm_v0m_n29), .A1(c0sm_v0m_n5), 
        .B0(c0sm_v0m_n4), .C0(c0sm_v0m_n8), .Y(c0sm_v0m_n58) );
  INV_X0P5B_A12TR c0sm_v0m_u34 ( .A(c0sm_v0m_state_queuelen_0_), .Y(
        c0sm_v0m_n23) );
  INV_X0P5B_A12TR c0sm_v0m_u33 ( .A(c0sm_v0m_full), .Y(c0sm_v0m_n26) );
  OAI31_X0P5M_A12TR c0sm_v0m_u32 ( .A0(c0sm_v0m_n29), .A1(tailout_1), .A2(
        c0sm_v0m_state_status_0_), .B0(c0sm_v0m_n5), .Y(c0sm_v0m_n28) );
  OAI31_X0P5M_A12TR c0sm_v0m_u31 ( .A0(c0sm_v0m_state_queuelen_0_), .A1(
        c0sm_v0m_state_queuelen_2_), .A2(c0sm_v0m_state_queuelen_1_), .B0(
        c0sm_v0m_n28), .Y(c0sm_v0m_n9) );
  NOR2_X0P5A_A12TR c0sm_v0m_u30 ( .A(c0sm_v0m_n9), .B(c0sm_n3), .Y(
        c0sm_v0m_n13) );
  INV_X0P5B_A12TR c0sm_v0m_u29 ( .A(c0sm_v0m_state_queuelen_2_), .Y(
        c0sm_v0m_n17) );
  NAND3_X0P5A_A12TR c0sm_v0m_u28 ( .A(c0sm_v0m_state_queuelen_0_), .B(
        c0sm_v0m_n17), .C(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n14) );
  NAND3_X0P5A_A12TR c0sm_v0m_u27 ( .A(c0sm_v0m_n14), .B(c0sm_v0m_n9), .C(
        c0sm_n3), .Y(c0sm_v0m_n18) );
  INV_X0P5B_A12TR c0sm_v0m_u26 ( .A(c0sm_v0m_n18), .Y(c0sm_v0m_n22) );
  AOI21_X0P5M_A12TR c0sm_v0m_u25 ( .A0(c0sm_v0m_n26), .A1(c0sm_v0m_n13), .B0(
        c0sm_v0m_n22), .Y(c0sm_v0m_n24) );
  XNOR2_X0P5M_A12TR c0sm_v0m_u24 ( .A(c0sm_v0m_n23), .B(c0sm_v0m_n24), .Y(
        c0sm_v0m_n27) );
  NOR2_X0P5A_A12TR c0sm_v0m_u23 ( .A(reset), .B(c0sm_v0m_n27), .Y(c0sm_v0m_n61) );
  NAND2_X0P5A_A12TR c0sm_v0m_u22 ( .A(c0sm_v0m_n13), .B(c0sm_v0m_n26), .Y(
        c0sm_v0m_n25) );
  MXIT2_X0P5M_A12TR c0sm_v0m_u21 ( .A(c0sm_v0m_n18), .B(c0sm_v0m_n25), .S0(
        c0sm_v0m_n23), .Y(c0sm_v0m_n20) );
  AOI21_X0P5M_A12TR c0sm_v0m_u20 ( .A0(c0sm_v0m_n23), .A1(c0sm_v0m_n22), .B0(
        c0sm_v0m_n24), .Y(c0sm_v0m_n16) );
  OAI21_X0P5M_A12TR c0sm_v0m_u19 ( .A0(c0sm_v0m_n22), .A1(c0sm_v0m_n23), .B0(
        c0sm_v0m_n16), .Y(c0sm_v0m_n21) );
  MXIT2_X0P5M_A12TR c0sm_v0m_u18 ( .A(c0sm_v0m_n20), .B(c0sm_v0m_n21), .S0(
        c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n19) );
  NOR2_X0P5A_A12TR c0sm_v0m_u17 ( .A(reset), .B(c0sm_v0m_n19), .Y(c0sm_v0m_n62) );
  MXIT2_X0P5M_A12TR c0sm_v0m_u16 ( .A(c0sm_v0m_state_queuelen_0_), .B(
        c0sm_v0m_n18), .S0(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n15) );
  AOI211_X0P5M_A12TR c0sm_v0m_u15 ( .A0(c0sm_v0m_n15), .A1(c0sm_v0m_n16), .B0(
        c0sm_v0m_n17), .C0(reset), .Y(c0sm_v0m_n63) );
  INV_X0P5B_A12TR c0sm_v0m_u14 ( .A(c0sm_v0m_n14), .Y(c0sm_v0m_n11) );
  INV_X0P5B_A12TR c0sm_v0m_u13 ( .A(c0sm_v0m_n13), .Y(c0sm_v0m_n12) );
  AOI32_X0P5M_A12TR c0sm_v0m_u12 ( .A0(c0sm_v0m_n11), .A1(c0sm_v0m_n9), .A2(
        c0sm_n3), .B0(c0sm_v0m_full), .B1(c0sm_v0m_n12), .Y(c0sm_v0m_n10) );
  NOR2_X0P5A_A12TR c0sm_v0m_u11 ( .A(reset), .B(c0sm_v0m_n10), .Y(c0sm_v0m_n64) );
  INV_X0P5B_A12TR c0sm_v0m_u10 ( .A(c0sm_v0m_n9), .Y(debitout_1) );
  INV_X0P5B_A12TR c0sm_v0m_u9 ( .A(c0sm_v0m_n8), .Y(c0sm_v0m_n1) );
  AND2_X0P5M_A12TR c0sm_v0m_u8 ( .A(swalloc_req_1[0]), .B(c0sm_v0m_n5), .Y(
        c0sm_v0m_n7) );
  MXIT2_X0P5M_A12TR c0sm_v0m_u7 ( .A(c0sm_v0m_n7), .B(c0sm_routewire[0]), .S0(
        c0sm_v0m_n4), .Y(c0sm_v0m_n6) );
  NOR2_X0P5A_A12TR c0sm_v0m_u6 ( .A(c0sm_v0m_n1), .B(c0sm_v0m_n6), .Y(
        c0sm_v0m_n33) );
  AND2_X0P5M_A12TR c0sm_v0m_u5 ( .A(swalloc_req_1[1]), .B(c0sm_v0m_n5), .Y(
        c0sm_v0m_n3) );
  MXIT2_X0P5M_A12TR c0sm_v0m_u4 ( .A(c0sm_v0m_n3), .B(c0sm_routewire[1]), .S0(
        c0sm_v0m_n4), .Y(c0sm_v0m_n2) );
  NOR2_X0P5A_A12TR c0sm_v0m_u3 ( .A(c0sm_v0m_n1), .B(c0sm_v0m_n2), .Y(
        c0sm_v0m_n32) );
  DFFQ_X1M_A12TR c0sm_v0m_state_queuelen_reg_1_ ( .D(c0sm_v0m_n62), .CK(clk), 
        .Q(c0sm_v0m_state_queuelen_1_) );
  DFFQ_X1M_A12TR c0sm_v0m_state_queuelen_reg_0_ ( .D(c0sm_v0m_n61), .CK(clk), 
        .Q(c0sm_v0m_state_queuelen_0_) );
  DFFQ_X1M_A12TR c0sm_v0m_state_status_reg_0_ ( .D(c0sm_v0m_n57), .CK(clk), 
        .Q(c0sm_v0m_state_status_0_) );
  DFFQ_X1M_A12TR c0sm_v0m_state_swreq_reg_1_ ( .D(c0sm_v0m_n32), .CK(clk), .Q(
        swalloc_req_1[1]) );
  DFFQ_X1M_A12TR c0sm_v0m_state_swreq_reg_0_ ( .D(c0sm_v0m_n33), .CK(clk), .Q(
        swalloc_req_1[0]) );
  DFFQ_X1M_A12TR c0sm_v0m_state_queuelen_reg_2_ ( .D(c0sm_v0m_n63), .CK(clk), 
        .Q(c0sm_v0m_state_queuelen_2_) );
  DFFQ_X1M_A12TR c0sm_v0m_full_reg ( .D(c0sm_v0m_n64), .CK(clk), .Q(
        c0sm_v0m_full) );
  DFFQ_X1M_A12TR c0sm_v0m_state_status_reg_1_ ( .D(c0sm_v0m_n58), .CK(clk), 
        .Q(c0sm_v0m_state_status_1_) );
  NAND2_X0P5A_A12TR s0m_u38 ( .A(debitout_1), .B(s0m_state_invc0_1_), .Y(
        s0m_n26) );
  INV_X0P5B_A12TR s0m_u37 ( .A(debitout_0), .Y(s0m_n21) );
  MXIT2_X0P5M_A12TR s0m_u36 ( .A(s0m_n26), .B(s0m_n21), .S0(s0m_state_invc0_0_), .Y(s0m_debit_outvc0) );
  NAND2_X0P5A_A12TR s0m_u35 ( .A(debitout_1), .B(s0m_state_invc1_1_), .Y(
        s0m_n20) );
  MXIT2_X0P5M_A12TR s0m_u34 ( .A(s0m_n20), .B(s0m_n21), .S0(s0m_state_invc1_0_), .Y(s0m_debit_outvc1) );
  INV_X0P5B_A12TR s0m_u33 ( .A(swalloc_resp_1[1]), .Y(s0m_n17) );
  NOR2_X0P5A_A12TR s0m_u32 ( .A(reset), .B(tailout_1), .Y(s0m_n16) );
  NAND2_X0P5A_A12TR s0m_u31 ( .A(s0m_outb1_1_), .B(s0m_n16), .Y(s0m_n18) );
  NOR2_X0P5A_A12TR s0m_u30 ( .A(swalloc_req_1[1]), .B(swalloc_req_1[0]), .Y(
        s0m_n19) );
  OAI31_X0P5M_A12TR s0m_u29 ( .A0(s0m_n19), .A1(swalloc_resp_1[1]), .A2(
        swalloc_resp_1[0]), .B0(s0m_n16), .Y(s0m_n15) );
  MXIT2_X0P5M_A12TR s0m_u28 ( .A(s0m_n17), .B(s0m_n18), .S0(s0m_n15), .Y(
        s0m_n22) );
  INV_X0P5B_A12TR s0m_u27 ( .A(swalloc_resp_1[0]), .Y(s0m_n13) );
  NAND2_X0P5A_A12TR s0m_u26 ( .A(s0m_outb0_1_), .B(s0m_n16), .Y(s0m_n14) );
  MXIT2_X0P5M_A12TR s0m_u25 ( .A(s0m_n13), .B(s0m_n14), .S0(s0m_n15), .Y(
        s0m_n23) );
  INV_X0P5B_A12TR s0m_u24 ( .A(swalloc_resp_0[1]), .Y(s0m_n10) );
  NOR2_X0P5A_A12TR s0m_u23 ( .A(reset), .B(tailout_0), .Y(s0m_n9) );
  NAND2_X0P5A_A12TR s0m_u22 ( .A(s0m_outb1_0_), .B(s0m_n9), .Y(s0m_n11) );
  NOR2_X0P5A_A12TR s0m_u21 ( .A(swalloc_req_0[1]), .B(swalloc_req_0[0]), .Y(
        s0m_n12) );
  OAI31_X0P5M_A12TR s0m_u20 ( .A0(s0m_n12), .A1(swalloc_resp_0[1]), .A2(
        swalloc_resp_0[0]), .B0(s0m_n9), .Y(s0m_n8) );
  MXIT2_X0P5M_A12TR s0m_u19 ( .A(s0m_n10), .B(s0m_n11), .S0(s0m_n8), .Y(
        s0m_n24) );
  INV_X0P5B_A12TR s0m_u18 ( .A(swalloc_resp_0[0]), .Y(s0m_n6) );
  NAND2_X0P5A_A12TR s0m_u17 ( .A(s0m_outb0_0_), .B(s0m_n9), .Y(s0m_n7) );
  MXIT2_X0P5M_A12TR s0m_u16 ( .A(s0m_n6), .B(s0m_n7), .S0(s0m_n8), .Y(s0m_n25)
         );
  INV_X0P5B_A12TR s0m_u15 ( .A(s0m_no_bufs1), .Y(s0m_n4) );
  INV_X0P5B_A12TR s0m_u14 ( .A(s0m_no_bufs0), .Y(s0m_n5) );
  MXIT2_X0P5M_A12TR s0m_u13 ( .A(s0m_n4), .B(s0m_n5), .S0(s0m_state_invc0_0_), 
        .Y(nomorebufs_0) );
  MXIT2_X0P5M_A12TR s0m_u12 ( .A(s0m_n4), .B(s0m_n5), .S0(s0m_state_invc0_1_), 
        .Y(nomorebufs_1) );
  AND2_X0P5M_A12TR s0m_u11 ( .A(s0m_elig_0_), .B(swalloc_req_0[0]), .Y(
        s0m_request0[0]) );
  AND2_X0P5M_A12TR s0m_u10 ( .A(s0m_elig_1_), .B(swalloc_req_0[1]), .Y(
        s0m_request0[1]) );
  AND2_X0P5M_A12TR s0m_u9 ( .A(s0m_elig_0_), .B(swalloc_req_1[0]), .Y(
        s0m_request1[0]) );
  AND2_X0P5M_A12TR s0m_u8 ( .A(s0m_elig_1_), .B(swalloc_req_1[1]), .Y(
        s0m_request1[1]) );
  NAND2_X0P5A_A12TR s0m_u7 ( .A(s0m_state_invc0_1_), .B(tailout_1), .Y(s0m_n3)
         );
  INV_X0P5B_A12TR s0m_u6 ( .A(tailout_0), .Y(s0m_n2) );
  MXIT2_X0P5M_A12TR s0m_u5 ( .A(s0m_n3), .B(s0m_n2), .S0(s0m_state_invc0_0_), 
        .Y(s0m_tail_outvc0) );
  NAND2_X0P5A_A12TR s0m_u4 ( .A(tailout_1), .B(s0m_state_invc1_1_), .Y(s0m_n1)
         );
  MXIT2_X0P5M_A12TR s0m_u3 ( .A(s0m_n1), .B(s0m_n2), .S0(s0m_state_invc1_0_), 
        .Y(s0m_tail_outvc1) );
  TIELO_X1M_A12TR s0m_u2 ( .Y(s0m__logic0_) );
  DFFQ_X1M_A12TR s0m_resp0_reg_0_ ( .D(s0m_n25), .CK(clk), .Q(
        swalloc_resp_0[0]) );
  DFFQ_X1M_A12TR s0m_resp0_reg_1_ ( .D(s0m_n24), .CK(clk), .Q(
        swalloc_resp_0[1]) );
  DFFQ_X1M_A12TR s0m_resp1_reg_0_ ( .D(s0m_n23), .CK(clk), .Q(
        swalloc_resp_1[0]) );
  DFFQ_X1M_A12TR s0m_resp1_reg_1_ ( .D(s0m_n22), .CK(clk), .Q(
        swalloc_resp_1[1]) );
  INV_X0P5B_A12TR s0m_m0m_u8 ( .A(s0m_request0[0]), .Y(s0m_m0m_n1) );
  AOI21_X0P5M_A12TR s0m_m0m_u7 ( .A0(s0m_request1[0]), .A1(s0m_m0m_row1_0_), 
        .B0(s0m_m0m_n1), .Y(s0m_outb0_0_) );
  AOI2XB1_X0P5M_A12TR s0m_m0m_u6 ( .A1N(s0m_request1[0]), .A0(s0m_m0m_row1_0_), 
        .B0(s0m_outb0_0_), .Y(s0m_m0m_n3) );
  XOR2_X0P5M_A12TR s0m_m0m_u5 ( .A(s0m__logic0_), .B(s0m_m0m_n3), .Y(
        s0m_m0m_n2) );
  NOR2_X0P5A_A12TR s0m_m0m_u4 ( .A(reset), .B(s0m_m0m_n2), .Y(s0m_m0m_n10) );
  OA21_X0P5M_A12TR s0m_m0m_u3 ( .A0(s0m_m0m_n1), .A1(s0m_m0m_row1_0_), .B0(
        s0m_request1[0]), .Y(s0m_outb0_1_) );
  DFFQ_X1M_A12TR s0m_m0m_state1_reg ( .D(s0m_m0m_n10), .CK(clk), .Q(
        s0m_m0m_row1_0_) );
  INV_X0P5B_A12TR s0m_m1m_u8 ( .A(s0m_request0[1]), .Y(s0m_m1m_n1) );
  AOI21_X0P5M_A12TR s0m_m1m_u7 ( .A0(s0m_request1[1]), .A1(s0m_m1m_row1_0_), 
        .B0(s0m_m1m_n1), .Y(s0m_outb1_0_) );
  AOI2XB1_X0P5M_A12TR s0m_m1m_u6 ( .A1N(s0m_request1[1]), .A0(s0m_m1m_row1_0_), 
        .B0(s0m_outb1_0_), .Y(s0m_m1m_n3) );
  XOR2_X0P5M_A12TR s0m_m1m_u5 ( .A(s0m__logic0_), .B(s0m_m1m_n3), .Y(
        s0m_m1m_n2) );
  NOR2_X0P5A_A12TR s0m_m1m_u4 ( .A(reset), .B(s0m_m1m_n2), .Y(s0m_m1m_n10) );
  OA21_X0P5M_A12TR s0m_m1m_u3 ( .A0(s0m_m1m_n1), .A1(s0m_m1m_row1_0_), .B0(
        s0m_request1[1]), .Y(s0m_outb1_1_) );
  DFFQ_X1M_A12TR s0m_m1m_state1_reg ( .D(s0m_m1m_n10), .CK(clk), .Q(
        s0m_m1m_row1_0_) );
  NOR2_X0P5A_A12TR s0m_o0nm_u35 ( .A(s0m_tail_outvc0), .B(reset), .Y(
        s0m_o0nm_n3) );
  OAI31_X0P5M_A12TR s0m_o0nm_u34 ( .A0(s0m_outb0_0_), .A1(
        s0m_o0nm_state_assigned), .A2(s0m_outb0_1_), .B0(s0m_o0nm_n3), .Y(
        s0m_o0nm_n25) );
  INV_X0P5B_A12TR s0m_o0nm_u33 ( .A(s0m_o0nm_n25), .Y(s0m_o0nm_n35) );
  NOR3_X0P5A_A12TR s0m_o0nm_u32 ( .A(s0m_outb0_1_), .B(s0m_outb0_0_), .C(
        s0m_debit_outvc0), .Y(s0m_o0nm_n9) );
  INV_X0P5B_A12TR s0m_o0nm_u31 ( .A(s0m_no_bufs0), .Y(s0m_o0nm_n10) );
  AND3_X0P5M_A12TR s0m_o0nm_u30 ( .A(s0m_o0nm_n9), .B(s0m_o0nm_n10), .C(
        creditin_0), .Y(s0m_o0nm_n23) );
  OR2_X0P5M_A12TR s0m_o0nm_u29 ( .A(s0m_o0nm_state_credits_1_), .B(
        s0m_o0nm_state_credits_0_), .Y(s0m_o0nm_n22) );
  NOR2_X0P5A_A12TR s0m_o0nm_u28 ( .A(s0m_o0nm_state_credits_2_), .B(
        s0m_o0nm_n22), .Y(s0m_o0nm_n12) );
  NOR3_X0P5A_A12TR s0m_o0nm_u27 ( .A(s0m_o0nm_n9), .B(creditin_0), .C(
        s0m_o0nm_n12), .Y(s0m_o0nm_n20) );
  NOR2_X0P5A_A12TR s0m_o0nm_u26 ( .A(s0m_o0nm_n23), .B(s0m_o0nm_n20), .Y(
        s0m_o0nm_n16) );
  XOR2_X0P5M_A12TR s0m_o0nm_u25 ( .A(s0m_o0nm_state_credits_0_), .B(
        s0m_o0nm_n16), .Y(s0m_o0nm_n24) );
  INV_X0P5B_A12TR s0m_o0nm_u24 ( .A(reset), .Y(s0m_o0nm_n8) );
  NAND2_X0P5A_A12TR s0m_o0nm_u23 ( .A(s0m_o0nm_n24), .B(s0m_o0nm_n8), .Y(
        s0m_o0nm_n36) );
  NAND2_X0P5A_A12TR s0m_o0nm_u22 ( .A(s0m_o0nm_state_credits_1_), .B(
        s0m_o0nm_state_credits_0_), .Y(s0m_o0nm_n18) );
  AO1B2_X0P5M_A12TR s0m_o0nm_u21 ( .B0(s0m_o0nm_n18), .B1(s0m_o0nm_n22), .A0N(
        s0m_o0nm_n20), .Y(s0m_o0nm_n19) );
  AOI32_X0P5M_A12TR s0m_o0nm_u20 ( .A0(s0m_o0nm_n22), .A1(s0m_o0nm_n18), .A2(
        s0m_o0nm_n23), .B0(s0m_o0nm_n16), .B1(s0m_o0nm_state_credits_1_), .Y(
        s0m_o0nm_n21) );
  NAND3_X0P5A_A12TR s0m_o0nm_u19 ( .A(s0m_o0nm_n19), .B(s0m_o0nm_n8), .C(
        s0m_o0nm_n21), .Y(s0m_o0nm_n37) );
  NOR3_X0P5A_A12TR s0m_o0nm_u18 ( .A(s0m_o0nm_n18), .B(s0m_o0nm_n20), .C(
        s0m_o0nm_n16), .Y(s0m_o0nm_n14) );
  XOR2_X0P5M_A12TR s0m_o0nm_u17 ( .A(s0m_o0nm_n18), .B(s0m_o0nm_n19), .Y(
        s0m_o0nm_n17) );
  NAND2B_X0P5M_A12TR s0m_o0nm_u16 ( .AN(s0m_o0nm_n16), .B(s0m_o0nm_n17), .Y(
        s0m_o0nm_n15) );
  MXIT2_X0P5M_A12TR s0m_o0nm_u15 ( .A(s0m_o0nm_n14), .B(s0m_o0nm_n15), .S0(
        s0m_o0nm_state_credits_2_), .Y(s0m_o0nm_n13) );
  NOR2_X0P5A_A12TR s0m_o0nm_u14 ( .A(reset), .B(s0m_o0nm_n13), .Y(s0m_o0nm_n38) );
  INV_X0P5B_A12TR s0m_o0nm_u13 ( .A(s0m_o0nm_n12), .Y(s0m_o0nm_n11) );
  NOR3_X0P5A_A12TR s0m_o0nm_u12 ( .A(s0m_o0nm_n11), .B(creditin_0), .C(
        s0m_o0nm_n9), .Y(s0m_o0nm_n6) );
  AOI21_X0P5M_A12TR s0m_o0nm_u11 ( .A0(creditin_0), .A1(s0m_o0nm_n9), .B0(
        s0m_o0nm_n10), .Y(s0m_o0nm_n7) );
  OA21_X0P5M_A12TR s0m_o0nm_u10 ( .A0(s0m_o0nm_n6), .A1(s0m_o0nm_n7), .B0(
        s0m_o0nm_n8), .Y(s0m_o0nm_n42) );
  NOR2_X0P5A_A12TR s0m_o0nm_u9 ( .A(s0m_o0nm_n42), .B(s0m_o0nm_n35), .Y(
        s0m_o0nm_n41) );
  INV_X0P5B_A12TR s0m_o0nm_u8 ( .A(s0m_outb0_1_), .Y(s0m_o0nm_n5) );
  AO21A1AI2_X0P5M_A12TR s0m_o0nm_u7 ( .A0(s0m_o0nm_n5), .A1(s0m_state_invc0_0_), .B0(s0m_outb0_0_), .C0(s0m_o0nm_n3), .Y(s0m_o0nm_n4) );
  INV_X0P5B_A12TR s0m_o0nm_u6 ( .A(s0m_o0nm_n4), .Y(s0m_o0nm_n30) );
  INV_X0P5B_A12TR s0m_o0nm_u5 ( .A(s0m_outb0_0_), .Y(s0m_o0nm_n2) );
  AO21A1AI2_X0P5M_A12TR s0m_o0nm_u4 ( .A0(s0m_o0nm_n2), .A1(s0m_state_invc0_1_), .B0(s0m_outb0_1_), .C0(s0m_o0nm_n3), .Y(s0m_o0nm_n1) );
  INV_X0P5B_A12TR s0m_o0nm_u3 ( .A(s0m_o0nm_n1), .Y(s0m_o0nm_n31) );
  DFFQ_X1M_A12TR s0m_o0nm_state_invc_reg_0_ ( .D(s0m_o0nm_n30), .CK(clk), .Q(
        s0m_state_invc0_0_) );
  DFFQ_X1M_A12TR s0m_o0nm_state_invc_reg_1_ ( .D(s0m_o0nm_n31), .CK(clk), .Q(
        s0m_state_invc0_1_) );
  DFFQ_X1M_A12TR s0m_o0nm_state_credits_reg_0_ ( .D(s0m_o0nm_n36), .CK(clk), 
        .Q(s0m_o0nm_state_credits_0_) );
  DFFQ_X1M_A12TR s0m_o0nm_state_credits_reg_1_ ( .D(s0m_o0nm_n37), .CK(clk), 
        .Q(s0m_o0nm_state_credits_1_) );
  DFFQ_X1M_A12TR s0m_o0nm_state_credits_reg_2_ ( .D(s0m_o0nm_n38), .CK(clk), 
        .Q(s0m_o0nm_state_credits_2_) );
  DFFQ_X1M_A12TR s0m_o0nm_no_bufs_reg ( .D(s0m_o0nm_n42), .CK(clk), .Q(
        s0m_no_bufs0) );
  DFFQ_X1M_A12TR s0m_o0nm_eligible_reg ( .D(s0m_o0nm_n41), .CK(clk), .Q(
        s0m_elig_0_) );
  DFFQ_X1M_A12TR s0m_o0nm_state_assigned_reg ( .D(s0m_o0nm_n35), .CK(clk), .Q(
        s0m_o0nm_state_assigned) );
  NOR2_X0P5A_A12TR s0m_o0sm_u35 ( .A(s0m_tail_outvc1), .B(reset), .Y(
        s0m_o0sm_n3) );
  OAI31_X0P5M_A12TR s0m_o0sm_u34 ( .A0(s0m_outb1_0_), .A1(
        s0m_o0sm_state_assigned), .A2(s0m_outb1_1_), .B0(s0m_o0sm_n3), .Y(
        s0m_o0sm_n25) );
  INV_X0P5B_A12TR s0m_o0sm_u33 ( .A(s0m_o0sm_n25), .Y(s0m_o0sm_n35) );
  NOR3_X0P5A_A12TR s0m_o0sm_u32 ( .A(s0m_outb1_1_), .B(s0m_outb1_0_), .C(
        s0m_debit_outvc1), .Y(s0m_o0sm_n9) );
  INV_X0P5B_A12TR s0m_o0sm_u31 ( .A(s0m_no_bufs1), .Y(s0m_o0sm_n10) );
  AND3_X0P5M_A12TR s0m_o0sm_u30 ( .A(s0m_o0sm_n9), .B(s0m_o0sm_n10), .C(
        creditin_1), .Y(s0m_o0sm_n23) );
  OR2_X0P5M_A12TR s0m_o0sm_u29 ( .A(s0m_o0sm_state_credits_1_), .B(
        s0m_o0sm_state_credits_0_), .Y(s0m_o0sm_n22) );
  NOR2_X0P5A_A12TR s0m_o0sm_u28 ( .A(s0m_o0sm_state_credits_2_), .B(
        s0m_o0sm_n22), .Y(s0m_o0sm_n12) );
  NOR3_X0P5A_A12TR s0m_o0sm_u27 ( .A(s0m_o0sm_n9), .B(creditin_1), .C(
        s0m_o0sm_n12), .Y(s0m_o0sm_n20) );
  NOR2_X0P5A_A12TR s0m_o0sm_u26 ( .A(s0m_o0sm_n23), .B(s0m_o0sm_n20), .Y(
        s0m_o0sm_n16) );
  XOR2_X0P5M_A12TR s0m_o0sm_u25 ( .A(s0m_o0sm_state_credits_0_), .B(
        s0m_o0sm_n16), .Y(s0m_o0sm_n24) );
  INV_X0P5B_A12TR s0m_o0sm_u24 ( .A(reset), .Y(s0m_o0sm_n8) );
  NAND2_X0P5A_A12TR s0m_o0sm_u23 ( .A(s0m_o0sm_n24), .B(s0m_o0sm_n8), .Y(
        s0m_o0sm_n36) );
  NAND2_X0P5A_A12TR s0m_o0sm_u22 ( .A(s0m_o0sm_state_credits_1_), .B(
        s0m_o0sm_state_credits_0_), .Y(s0m_o0sm_n18) );
  AO1B2_X0P5M_A12TR s0m_o0sm_u21 ( .B0(s0m_o0sm_n18), .B1(s0m_o0sm_n22), .A0N(
        s0m_o0sm_n20), .Y(s0m_o0sm_n19) );
  AOI32_X0P5M_A12TR s0m_o0sm_u20 ( .A0(s0m_o0sm_n22), .A1(s0m_o0sm_n18), .A2(
        s0m_o0sm_n23), .B0(s0m_o0sm_n16), .B1(s0m_o0sm_state_credits_1_), .Y(
        s0m_o0sm_n21) );
  NAND3_X0P5A_A12TR s0m_o0sm_u19 ( .A(s0m_o0sm_n19), .B(s0m_o0sm_n8), .C(
        s0m_o0sm_n21), .Y(s0m_o0sm_n37) );
  NOR3_X0P5A_A12TR s0m_o0sm_u18 ( .A(s0m_o0sm_n18), .B(s0m_o0sm_n20), .C(
        s0m_o0sm_n16), .Y(s0m_o0sm_n14) );
  XOR2_X0P5M_A12TR s0m_o0sm_u17 ( .A(s0m_o0sm_n18), .B(s0m_o0sm_n19), .Y(
        s0m_o0sm_n17) );
  NAND2B_X0P5M_A12TR s0m_o0sm_u16 ( .AN(s0m_o0sm_n16), .B(s0m_o0sm_n17), .Y(
        s0m_o0sm_n15) );
  MXIT2_X0P5M_A12TR s0m_o0sm_u15 ( .A(s0m_o0sm_n14), .B(s0m_o0sm_n15), .S0(
        s0m_o0sm_state_credits_2_), .Y(s0m_o0sm_n13) );
  NOR2_X0P5A_A12TR s0m_o0sm_u14 ( .A(reset), .B(s0m_o0sm_n13), .Y(s0m_o0sm_n38) );
  INV_X0P5B_A12TR s0m_o0sm_u13 ( .A(s0m_o0sm_n12), .Y(s0m_o0sm_n11) );
  NOR3_X0P5A_A12TR s0m_o0sm_u12 ( .A(s0m_o0sm_n11), .B(creditin_1), .C(
        s0m_o0sm_n9), .Y(s0m_o0sm_n6) );
  AOI21_X0P5M_A12TR s0m_o0sm_u11 ( .A0(creditin_1), .A1(s0m_o0sm_n9), .B0(
        s0m_o0sm_n10), .Y(s0m_o0sm_n7) );
  OA21_X0P5M_A12TR s0m_o0sm_u10 ( .A0(s0m_o0sm_n6), .A1(s0m_o0sm_n7), .B0(
        s0m_o0sm_n8), .Y(s0m_o0sm_n42) );
  NOR2_X0P5A_A12TR s0m_o0sm_u9 ( .A(s0m_o0sm_n42), .B(s0m_o0sm_n35), .Y(
        s0m_o0sm_n41) );
  INV_X0P5B_A12TR s0m_o0sm_u8 ( .A(s0m_outb1_1_), .Y(s0m_o0sm_n5) );
  AO21A1AI2_X0P5M_A12TR s0m_o0sm_u7 ( .A0(s0m_o0sm_n5), .A1(s0m_state_invc1_0_), .B0(s0m_outb1_0_), .C0(s0m_o0sm_n3), .Y(s0m_o0sm_n4) );
  INV_X0P5B_A12TR s0m_o0sm_u6 ( .A(s0m_o0sm_n4), .Y(s0m_o0sm_n27) );
  INV_X0P5B_A12TR s0m_o0sm_u5 ( .A(s0m_outb1_0_), .Y(s0m_o0sm_n2) );
  AO21A1AI2_X0P5M_A12TR s0m_o0sm_u4 ( .A0(s0m_o0sm_n2), .A1(s0m_state_invc1_1_), .B0(s0m_outb1_1_), .C0(s0m_o0sm_n3), .Y(s0m_o0sm_n1) );
  INV_X0P5B_A12TR s0m_o0sm_u3 ( .A(s0m_o0sm_n1), .Y(s0m_o0sm_n26) );
  DFFQ_X1M_A12TR s0m_o0sm_state_invc_reg_0_ ( .D(s0m_o0sm_n27), .CK(clk), .Q(
        s0m_state_invc1_0_) );
  DFFQ_X1M_A12TR s0m_o0sm_state_credits_reg_0_ ( .D(s0m_o0sm_n36), .CK(clk), 
        .Q(s0m_o0sm_state_credits_0_) );
  DFFQ_X1M_A12TR s0m_o0sm_state_invc_reg_1_ ( .D(s0m_o0sm_n26), .CK(clk), .Q(
        s0m_state_invc1_1_) );
  DFFQ_X1M_A12TR s0m_o0sm_state_credits_reg_1_ ( .D(s0m_o0sm_n37), .CK(clk), 
        .Q(s0m_o0sm_state_credits_1_) );
  DFFQ_X1M_A12TR s0m_o0sm_state_credits_reg_2_ ( .D(s0m_o0sm_n38), .CK(clk), 
        .Q(s0m_o0sm_state_credits_2_) );
  DFFQ_X1M_A12TR s0m_o0sm_no_bufs_reg ( .D(s0m_o0sm_n42), .CK(clk), .Q(
        s0m_no_bufs1) );
  DFFQ_X1M_A12TR s0m_o0sm_eligible_reg ( .D(s0m_o0sm_n41), .CK(clk), .Q(
        s0m_elig_1_) );
  DFFQ_X1M_A12TR s0m_o0sm_state_assigned_reg ( .D(s0m_o0sm_n35), .CK(clk), .Q(
        s0m_o0sm_state_assigned) );
  NAND2B_X0P5M_A12TR d0m_u2 ( .AN(swalloc_resp_1[0]), .B(swalloc_resp_0[0]), 
        .Y(colsel0[0]) );
  NOR2_X0P5A_A12TR d0m_u1 ( .A(swalloc_resp_1[0]), .B(swalloc_resp_0[0]), .Y(
        colsel0[1]) );
  NAND2B_X0P5M_A12TR d1m_u2 ( .AN(swalloc_resp_1[1]), .B(swalloc_resp_0[1]), 
        .Y(colsel1[0]) );
  NOR2_X0P5A_A12TR d1m_u1 ( .A(swalloc_resp_1[1]), .B(swalloc_resp_0[1]), .Y(
        colsel1[1]) );
  OR2_X0P5M_A12TR x0m_u8 ( .A(colsel0[0]), .B(reset), .Y(x0m_n3) );
  OR2_X0P5M_A12TR x0m_u7 ( .A(colsel0[1]), .B(reset), .Y(x0m_n4) );
  OR2_X0P5M_A12TR x0m_u6 ( .A(colsel1[0]), .B(reset), .Y(x0m_n5) );
  OR2_X0P5M_A12TR x0m_u5 ( .A(colsel1[1]), .B(reset), .Y(x0m_n6) );
  TIEHI_X1M_A12TR x0m_u4 ( .Y(x0m__logic1_) );
  TIELO_X1M_A12TR x0m_u3 ( .Y(x0m__logic0_) );
  DFFQ_X1M_A12TR x0m_colsel0reg_reg_0_ ( .D(x0m_n3), .CK(clk), .Q(
        x0m_colsel0reg_0_) );
  DFFQ_X1M_A12TR x0m_colsel0reg_reg_1_ ( .D(x0m_n4), .CK(clk), .Q(
        x0m_colsel0reg_1_) );
  DFFQ_X1M_A12TR x0m_colsel1reg_reg_0_ ( .D(x0m_n5), .CK(clk), .Q(
        x0m_colsel1reg_0_) );
  DFFQ_X1M_A12TR x0m_colsel1reg_reg_1_ ( .D(x0m_n6), .CK(clk), .Q(
        x0m_colsel1reg_1_) );
  MXT2_X0P5M_A12TR x0m_bx0m_m0m_m0m_u1 ( .A(flitout_switch_0[0]), .B(
        flitout_switch_1[0]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx0m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx0m_m0m_m4m_u1 ( .A(x0m_bx0m_m0m_int01), .B(
        x0m__logic1_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[0]) );
  MXT2_X0P5M_A12TR x0m_bx0m_m1m_m0m_u1 ( .A(flitout_switch_0[0]), .B(
        flitout_switch_1[0]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx0m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx0m_m1m_m4m_u1 ( .A(x0m_bx0m_m1m_int01), .B(
        x0m__logic1_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[0]) );
  MXT2_X0P5M_A12TR x0m_bx1m_m0m_m0m_u1 ( .A(flitout_switch_0[1]), .B(
        flitout_switch_1[1]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx1m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx1m_m0m_m4m_u1 ( .A(x0m_bx1m_m0m_int01), .B(
        x0m__logic1_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[1]) );
  MXT2_X0P5M_A12TR x0m_bx1m_m1m_m0m_u1 ( .A(flitout_switch_0[1]), .B(
        flitout_switch_1[1]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx1m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx1m_m1m_m4m_u1 ( .A(x0m_bx1m_m1m_int01), .B(
        x0m__logic1_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[1]) );
  MXT2_X0P5M_A12TR x0m_bx2m_m0m_m0m_u1 ( .A(flitout_switch_0[2]), .B(
        flitout_switch_1[2]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx2m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx2m_m0m_m4m_u1 ( .A(x0m_bx2m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[2]) );
  MXT2_X0P5M_A12TR x0m_bx2m_m1m_m0m_u1 ( .A(flitout_switch_0[2]), .B(
        flitout_switch_1[2]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx2m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx2m_m1m_m4m_u1 ( .A(x0m_bx2m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[2]) );
  MXT2_X0P5M_A12TR x0m_bx3m_m0m_m0m_u1 ( .A(flitout_switch_0[3]), .B(
        flitout_switch_1[3]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx3m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx3m_m0m_m4m_u1 ( .A(x0m_bx3m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[3]) );
  MXT2_X0P5M_A12TR x0m_bx3m_m1m_m0m_u1 ( .A(flitout_switch_0[3]), .B(
        flitout_switch_1[3]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx3m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx3m_m1m_m4m_u1 ( .A(x0m_bx3m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[3]) );
  MXT2_X0P5M_A12TR x0m_bx4m_m0m_m0m_u1 ( .A(flitout_switch_0[4]), .B(
        flitout_switch_1[4]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx4m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx4m_m0m_m4m_u1 ( .A(x0m_bx4m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[4]) );
  MXT2_X0P5M_A12TR x0m_bx4m_m1m_m0m_u1 ( .A(flitout_switch_0[4]), .B(
        flitout_switch_1[4]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx4m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx4m_m1m_m4m_u1 ( .A(x0m_bx4m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[4]) );
  MXT2_X0P5M_A12TR x0m_bx5m_m0m_m0m_u1 ( .A(flitout_switch_0[5]), .B(
        flitout_switch_1[5]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx5m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx5m_m0m_m4m_u1 ( .A(x0m_bx5m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[5]) );
  MXT2_X0P5M_A12TR x0m_bx5m_m1m_m0m_u1 ( .A(flitout_switch_0[5]), .B(
        flitout_switch_1[5]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx5m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx5m_m1m_m4m_u1 ( .A(x0m_bx5m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[5]) );
  MXT2_X0P5M_A12TR x0m_bx6m_m0m_m0m_u1 ( .A(flitout_switch_0[6]), .B(
        flitout_switch_1[6]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx6m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx6m_m0m_m4m_u1 ( .A(x0m_bx6m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[6]) );
  MXT2_X0P5M_A12TR x0m_bx6m_m1m_m0m_u1 ( .A(flitout_switch_0[6]), .B(
        flitout_switch_1[6]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx6m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx6m_m1m_m4m_u1 ( .A(x0m_bx6m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[6]) );
  MXT2_X0P5M_A12TR x0m_bx7m_m0m_m0m_u1 ( .A(flitout_switch_0[7]), .B(
        flitout_switch_1[7]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx7m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx7m_m0m_m4m_u1 ( .A(x0m_bx7m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[7]) );
  MXT2_X0P5M_A12TR x0m_bx7m_m1m_m0m_u1 ( .A(flitout_switch_0[7]), .B(
        flitout_switch_1[7]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx7m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx7m_m1m_m4m_u1 ( .A(x0m_bx7m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[7]) );
  MXT2_X0P5M_A12TR x0m_bx8m_m0m_m0m_u1 ( .A(flitout_switch_0[8]), .B(
        flitout_switch_1[8]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx8m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx8m_m0m_m4m_u1 ( .A(x0m_bx8m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[8]) );
  MXT2_X0P5M_A12TR x0m_bx8m_m1m_m0m_u1 ( .A(flitout_switch_0[8]), .B(
        flitout_switch_1[8]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx8m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx8m_m1m_m4m_u1 ( .A(x0m_bx8m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[8]) );
  MXT2_X0P5M_A12TR x0m_bx9m_m0m_m0m_u1 ( .A(flitout_switch_0[9]), .B(
        flitout_switch_1[9]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx9m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx9m_m0m_m4m_u1 ( .A(x0m_bx9m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[9]) );
  MXT2_X0P5M_A12TR x0m_bx9m_m1m_m0m_u1 ( .A(flitout_switch_0[9]), .B(
        flitout_switch_1[9]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx9m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx9m_m1m_m4m_u1 ( .A(x0m_bx9m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[9]) );
  MXT2_X0P5M_A12TR x0m_bx10m_m0m_m0m_u1 ( .A(flitout_switch_0[10]), .B(
        flitout_switch_1[10]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx10m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx10m_m0m_m4m_u1 ( .A(x0m_bx10m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[10]) );
  MXT2_X0P5M_A12TR x0m_bx10m_m1m_m0m_u1 ( .A(flitout_switch_0[10]), .B(
        flitout_switch_1[10]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx10m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx10m_m1m_m4m_u1 ( .A(x0m_bx10m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[10]) );
  MXT2_X0P5M_A12TR x0m_bx11m_m0m_m0m_u1 ( .A(flitout_switch_0[11]), .B(
        flitout_switch_1[11]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx11m_m0m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx11m_m0m_m4m_u1 ( .A(x0m_bx11m_m0m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[11]) );
  MXT2_X0P5M_A12TR x0m_bx11m_m1m_m0m_u1 ( .A(flitout_switch_0[11]), .B(
        flitout_switch_1[11]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx11m_m1m_int01)
         );
  MXT2_X0P5M_A12TR x0m_bx11m_m1m_m4m_u1 ( .A(x0m_bx11m_m1m_int01), .B(
        x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[11]) );
endmodule

