
module ae18_core ( wb_clk_o, wb_rst_o, iwb_adr_o, iwb_dat_o, iwb_stb_o, 
        iwb_we_o, iwb_sel_o, dwb_adr_o, dwb_dat_o, dwb_stb_o, dwb_we_o, 
        iwb_dat_i, iwb_ack_i, dwb_dat_i, dwb_ack_i, int_i, inte_i, clk_i, 
        rst_i );
  output [19:0] iwb_adr_o;
  output [15:0] iwb_dat_o;
  output [1:0] iwb_sel_o;
  output [11:0] dwb_adr_o;
  output [7:0] dwb_dat_o;
  input [15:0] iwb_dat_i;
  input [7:0] dwb_dat_i;
  input [1:0] int_i;
  input [7:6] inte_i;
  input iwb_ack_i, dwb_ack_i, clk_i, rst_i;
  output wb_clk_o, wb_rst_o, iwb_stb_o, iwb_we_o, dwb_stb_o, dwb_we_o;
  wire   n214, n215, n216, n217, n218, wb_clk_o, qrst, rclrwdt, rsleep,
         rswdten, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n262, rpcu_4_, rpcl_0_,
         rnskp, rbcc, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, rsfrstb, wrrc_7_, rc_,
         rclrwdt_, rsleep_, n845, n846, rreset_, rz, rov, rn, rstkptr_5_, rdc,
         rstkful, rstkunf, n17820, n1783, n17840, n1785, n1786, n17870, n1788,
         n1789, n17900, n1791, n1792, n1793, n1794, n1795, n1796, n17970,
         n1413, n1414, n1415, n1416, n1417, n1419, n1420, n1421, n1423, n1426,
         n1427, n1428, n1430, n1433, n1434, n1435, n1437, n1440, n1443, n1444,
         n1446, n1448, n1450, n1452, n1454, n1456, n1458, n1459, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1471, n1481, n1495,
         n1497, n1499, n1501, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1513, n1514, n1516, n1517, n1519, n1520, n1522, n1523,
         n1525, n1526, n1528, n1529, n1531, n1532, n1534, n1535, n1537, n1538,
         n1540, n1541, n1543, n1544, n1546, n1547, n1548, n1550, n1552, n1553,
         n1555, n1556, n1558, n1559, n1560, n1562, n1563, n1564, n1566, n1567,
         n1568, n1570, n1571, n1572, n1574, n1575, n1576, n1578, n1579, n1580,
         n1582, n1583, n1584, n1586, n1587, n1588, n1589, n1591, n1592, n1594,
         n1595, n1597, n1599, n1601, n1603, n1605, n1607, n1608, n1610, n1611,
         n1613, n1614, n1616, n1617, n1619, n1620, n1622, n1623, n1625, n1626,
         n1628, n1629, n1631, n1632, n1634, n1636, n1638, n1640, n1642, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1658, n1660, n1662, n1676, n1678, n1680, n1682, n1684,
         n1691, n1693, n1695, n1697, n1699, n1701, n1703, n1705, n1708, n1710,
         n1713, n1715, n1717, n1719, n1722, n1724, n1727, n1730, n1733, n1736,
         n1739, n1741, n1743, n1747, n1749, n1751, n1753, n1755, n1757, n1759,
         n1762, n1764, n1766, n1768, n1770, n1772, n1774, n1776, n1778, n1780,
         n17821, n17841, n17871, n17901, n17971, n1799, n1801, n1803, n1805,
         n1807, n1809, n1829, n1831, n1833, n1835, n1836, n1838, n1840, n1843,
         n1846, n1847, n1849, n1851, n1853, n1854, n1856, n1858, n1861, n1862,
         n1864, n1866, n1868, n1869, n1870, n1871, n1872, n1873, n1875, n1877,
         n1879, n1881, n1883, n1885, n1887, n1889, n1891, n1893, n1895, n1897,
         n1899, n1901, n1902, n1904, n1906, n3, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1940, n1941, n1942, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, sub_1479_n10, sub_1479_n9,
         sub_1479_n8, sub_1479_n7, sub_1479_n6, sub_1479_n5, sub_1479_n4,
         sub_1479_n3, sub_1479_n2, sub_1479_n1, sub_1552_n18, sub_1552_n17,
         sub_1552_n16, sub_1552_n15, sub_1552_n14, sub_1552_n13, sub_1552_n12,
         sub_1552_n11, sub_1552_n10, sub_1552_n9, sub_1552_n8, sub_1552_n7,
         sub_1552_n6, sub_1552_n5, sub_1552_n4, sub_1552_n3, sub_1552_n2,
         sub_1552_n1, sub_1478_n10, sub_1478_n9, sub_1478_n8, sub_1478_n7,
         sub_1478_n6, sub_1478_n5, sub_1478_n4, sub_1478_n3, sub_1478_n2,
         sub_1478_n1, add_1151_n4, add_1151_n3, add_1151_n2, add_1151_n1,
         add_1151_carry_2_, add_1151_carry_3_, add_1151_carry_4_,
         add_1151_carry_5_, add_1151_carry_6_, add_1151_carry_7_,
         add_1151_carry_8_, add_1150_n4, add_1150_n3, add_1150_n2, add_1150_n1,
         add_1150_carry_2_, add_1150_carry_3_, add_1150_carry_4_,
         add_1150_carry_5_, add_1150_carry_6_, add_1150_carry_7_,
         add_1150_carry_8_, sub_1006_n10, sub_1006_n9, sub_1006_n8,
         sub_1006_n7, sub_1006_n6, sub_1006_n5, sub_1006_n4, sub_1006_n3,
         sub_1006_n1, add_1004_n1, add_436_n1, sub_1477_n10, sub_1477_n9,
         sub_1477_n8, sub_1477_n7, sub_1477_n6, sub_1477_n5, sub_1477_n4,
         sub_1477_n3, sub_1477_n2, sub_1477_n1, add_1152_n4, add_1152_n3,
         add_1152_n2, add_1152_n1, add_1152_carry_2_, add_1152_carry_3_,
         add_1152_carry_4_, add_1152_carry_5_, add_1152_carry_6_,
         add_1152_carry_7_, add_1152_carry_8_, mult_1536_n177, mult_1536_n176,
         mult_1536_n175, mult_1536_n174, mult_1536_n173, mult_1536_n172,
         mult_1536_n171, mult_1536_n170, mult_1536_n169, mult_1536_n168,
         mult_1536_n167, mult_1536_n166, mult_1536_n165, mult_1536_n164,
         mult_1536_n163, mult_1536_n162, mult_1536_n161, mult_1536_n160,
         mult_1536_n159, mult_1536_n158, mult_1536_n157, mult_1536_n156,
         mult_1536_n155, mult_1536_n154, mult_1536_n153, mult_1536_n152,
         mult_1536_n151, mult_1536_n150, mult_1536_n149, mult_1536_n148,
         mult_1536_n147, mult_1536_n146, mult_1536_n145, mult_1536_n144,
         mult_1536_n143, mult_1536_n142, mult_1536_n141, mult_1536_n140,
         mult_1536_n139, mult_1536_n138, mult_1536_n137, mult_1536_n136,
         mult_1536_n135, mult_1536_n134, mult_1536_n133, mult_1536_n132,
         mult_1536_n131, mult_1536_n130, mult_1536_n129, mult_1536_n128,
         mult_1536_n127, mult_1536_n126, mult_1536_n125, mult_1536_n124,
         mult_1536_n123, mult_1536_n122, mult_1536_n121, mult_1536_n120,
         mult_1536_n119, mult_1536_n118, mult_1536_n117, mult_1536_n116,
         mult_1536_n115, mult_1536_n114, mult_1536_n113, mult_1536_n112,
         mult_1536_n111, mult_1536_n110, mult_1536_n109, mult_1536_n108,
         mult_1536_n107, mult_1536_n106, mult_1536_n105, mult_1536_n104,
         mult_1536_n103, mult_1536_n102, mult_1536_n101, mult_1536_n100,
         mult_1536_n99, mult_1536_n98, mult_1536_n97, mult_1536_n96,
         mult_1536_n95, mult_1536_n94, mult_1536_n93, mult_1536_n92,
         mult_1536_n91, mult_1536_n90, mult_1536_n89, mult_1536_n88,
         mult_1536_n87, mult_1536_n86, mult_1536_n85, mult_1536_n84,
         mult_1536_n83, mult_1536_n82, mult_1536_n81, mult_1536_n80,
         mult_1536_n79, mult_1536_n78, mult_1536_n77, mult_1536_n76,
         mult_1536_n75, mult_1536_n74, mult_1536_n73, mult_1536_n72,
         mult_1536_n71, mult_1536_n70, mult_1536_n69, mult_1536_n68,
         mult_1536_n67, mult_1536_n66, mult_1536_n65, mult_1536_n64,
         mult_1536_n63, mult_1536_n62, mult_1536_n61, mult_1536_n60,
         mult_1536_n59, mult_1536_n58, mult_1536_n57, mult_1536_n56,
         mult_1536_n55, mult_1536_n54, mult_1536_n53, mult_1536_n52,
         mult_1536_n51, mult_1536_n50, mult_1536_n49, mult_1536_n48,
         mult_1536_n47, mult_1536_n46, mult_1536_n45, mult_1536_n44,
         mult_1536_n43, mult_1536_n42, mult_1536_n41, mult_1536_n40,
         mult_1536_n39, mult_1536_n38, mult_1536_n37, mult_1536_n36,
         mult_1536_n35, mult_1536_n34, mult_1536_n33, mult_1536_n32,
         mult_1536_n31, mult_1536_n30, mult_1536_n29, mult_1536_n28,
         mult_1536_n27, mult_1536_n26, mult_1536_n25, mult_1536_n24,
         mult_1536_n23, mult_1536_n22, mult_1536_n21, mult_1536_n20,
         mult_1536_n19, mult_1536_n18, mult_1536_n17, mult_1536_n16,
         mult_1536_n15, mult_1536_n14, mult_1536_n13, mult_1536_n12,
         mult_1536_n11, mult_1536_n10, mult_1536_n9, mult_1536_n8,
         mult_1536_n7, mult_1536_n6, mult_1536_n5, mult_1536_n4, mult_1536_n3,
         mult_1536_n2;
  wire   [16:0] rwdt;
  wire   [7:0] rprng;
  wire   [1:0] rfsm;
  wire   [3:0] qena;
  wire   [1:0] qfsm;
  wire   [2:0] rinth;
  wire   [2:0] rintl;
  wire   [1:0] rintf;
  wire   [1:0] rnxt;
  wire   [18:0] wpclat;
  wire   [18:0] rpcnxt;
  wire   [3:0] rmxtbl;
  wire   [7:4] rtblptru;
  wire   [18:0] wpcinc;
  wire   [10:0] rireg;
  wire   [15:0] rromlat;
  wire   [7:4] rtosu;
  wire   [2:0] rmxnpc;
  wire   [7:0] rilat;
  wire   [15:0] reaptr;
  wire   [1:0] rmxbsr;
  wire   [3:0] rmxalu;
  wire   [2:0] rmxbcc;
  wire   [1:0] rmxdst;
  wire   [3:0] rmxfsr;
  wire   [1:0] rmxsha;
  wire   [2:0] rmxskp;
  wire   [1:0] rmxsrc;
  wire   [2:0] rmxsta;
  wire   [1:0] rmxstk;
  wire   [1:0] rmxtgt;
  wire   [15:8] wfilebsr;
  wire   [7:0] rmask;
  wire   [7:0] rsfrdat;
  wire   [7:0] rwreg;
  wire   [7:0] rsrc;
  wire   [7:1] rtgt;
  wire   [8:0] wadd;
  wire   [8:0] waddc;
  wire   [8:0] wsub;
  wire   [8:0] wsubc;
  wire   [7:0] wneg;
  wire   [15:12] rdwbadr;
  wire   [7:0] rfsr0h;
  wire   [7:0] rfsr0l;
  wire   [11:0] wfsrinc0;
  wire   [7:0] rfsr1h;
  wire   [7:0] rfsr1l;
  wire   [11:0] wfsrinc1;
  wire   [4:0] rfsr2h;
  wire   [7:0] rfsr2l;
  wire   [11:0] wfsrinc2;
  wire   [11:0] wfsrplusw0;
  wire   [11:0] wfsrplusw1;
  wire   [11:0] wfsrplusw2;
  wire   [19:0] wstkw;
  wire   [639:0] rstkram;
  wire   [4:0] rstkptr_;
  wire   [7:0] rprodl;
  wire   [7:0] rprodh;
  wire   [7:0] rpclath;
  wire   [7:0] rpclatu;
  wire   [4:1] wstkinc;
  wire   [4:1] wstkdec;
  wire   [7:0] rbsr_;
  wire   [4:0] rstatus_;
  wire   [7:0] rwreg_;
  wire   [2:0] rmxstal;
  wire   [11:0] wfsrdec0;
  wire   [11:0] wfsrdec1;
  wire   [11:0] wfsrdec2;
  wire   [19:0] wtblinc;
  wire   [19:0] wtblat;
  wire   [19:0] wtbldec;
  wire   [18:2] add_434_carry;
  wire   [5:2] add_1310_carry;
  wire   [19:2] add_1550_carry;
  wire   [11:2] add_1149_carry;
  wire   [11:2] add_1148_carry;
  wire   [11:2] add_1147_carry;
  wire   [8:2] sub_1006_carry;
  wire   [7:2] add_1004_carry;
  wire   [18:2] add_436_carry;
  wire   [18:2] add_433_carry;
  wire   [16:2] add_276_carry;
  assign wb_clk_o = clk_i;
  assign iwb_dat_o[6] = iwb_dat_o[14];
  assign iwb_dat_o[5] = iwb_dat_o[13];
  assign iwb_dat_o[4] = iwb_dat_o[12];
  assign iwb_dat_o[3] = iwb_dat_o[11];
  assign iwb_dat_o[2] = iwb_dat_o[10];
  assign iwb_dat_o[1] = iwb_dat_o[9];
  assign iwb_dat_o[0] = iwb_dat_o[8];
  assign iwb_dat_o[7] = iwb_dat_o[15];

  DFFRPQ_X4M_A12TR rstkptr_reg_1_ ( .D(n1415), .CK(wb_clk_o), .R(n2803), .Q(
        n215) );
  ADDF_X1M_A12TR add_434_u1_1 ( .A(iwb_adr_o[2]), .B(rireg[1]), .CI(n2786), 
        .CO(add_434_carry[2]), .S(n367) );
  ADDF_X1M_A12TR add_434_u1_2 ( .A(iwb_adr_o[3]), .B(rireg[2]), .CI(
        add_434_carry[2]), .CO(add_434_carry[3]), .S(n368) );
  ADDF_X1M_A12TR add_434_u1_3 ( .A(iwb_adr_o[4]), .B(rireg[3]), .CI(
        add_434_carry[3]), .CO(add_434_carry[4]), .S(n369) );
  ADDF_X1M_A12TR add_434_u1_4 ( .A(iwb_adr_o[5]), .B(rireg[4]), .CI(
        add_434_carry[4]), .CO(add_434_carry[5]), .S(n370) );
  ADDF_X1M_A12TR add_434_u1_5 ( .A(iwb_adr_o[6]), .B(rireg[5]), .CI(
        add_434_carry[5]), .CO(add_434_carry[6]), .S(n371) );
  ADDF_X1M_A12TR add_434_u1_6 ( .A(iwb_adr_o[7]), .B(rireg[6]), .CI(
        add_434_carry[6]), .CO(add_434_carry[7]), .S(n372) );
  ADDF_X1M_A12TR add_434_u1_7 ( .A(iwb_adr_o[8]), .B(rireg[7]), .CI(
        add_434_carry[7]), .CO(add_434_carry[8]), .S(n373) );
  ADDF_X1M_A12TR add_434_u1_8 ( .A(iwb_adr_o[9]), .B(rireg[7]), .CI(
        add_434_carry[8]), .CO(add_434_carry[9]), .S(n374) );
  ADDF_X1M_A12TR add_434_u1_9 ( .A(iwb_adr_o[10]), .B(rireg[7]), .CI(
        add_434_carry[9]), .CO(add_434_carry[10]), .S(n375) );
  ADDF_X1M_A12TR add_434_u1_10 ( .A(iwb_adr_o[11]), .B(rireg[7]), .CI(
        add_434_carry[10]), .CO(add_434_carry[11]), .S(n376) );
  ADDF_X1M_A12TR add_434_u1_11 ( .A(iwb_adr_o[12]), .B(rireg[7]), .CI(
        add_434_carry[11]), .CO(add_434_carry[12]), .S(n377) );
  ADDF_X1M_A12TR add_434_u1_12 ( .A(iwb_adr_o[13]), .B(rireg[7]), .CI(
        add_434_carry[12]), .CO(add_434_carry[13]), .S(n378) );
  ADDF_X1M_A12TR add_434_u1_13 ( .A(iwb_adr_o[14]), .B(rireg[7]), .CI(
        add_434_carry[13]), .CO(add_434_carry[14]), .S(n379) );
  ADDF_X1M_A12TR add_434_u1_14 ( .A(iwb_adr_o[15]), .B(rireg[7]), .CI(
        add_434_carry[14]), .CO(add_434_carry[15]), .S(n380) );
  ADDF_X1M_A12TR add_434_u1_15 ( .A(iwb_adr_o[16]), .B(rireg[7]), .CI(
        add_434_carry[15]), .CO(add_434_carry[16]), .S(n381) );
  ADDF_X1M_A12TR add_434_u1_16 ( .A(iwb_adr_o[17]), .B(rireg[7]), .CI(
        add_434_carry[16]), .CO(add_434_carry[17]), .S(n382) );
  ADDF_X1M_A12TR add_434_u1_17 ( .A(iwb_adr_o[18]), .B(rireg[7]), .CI(
        add_434_carry[17]), .CO(add_434_carry[18]), .S(n383) );
  ADDF_X1M_A12TR add_434_u1_18 ( .A(iwb_adr_o[19]), .B(rireg[7]), .CI(
        add_434_carry[18]), .CO(), .S(n384) );
  DFFQ_X1M_A12TR rstkram_reg_31__3_ ( .D(n2190), .CK(wb_clk_o), .Q(rstkram[3])
         );
  DFFQ_X1M_A12TR rstkram_reg_31__2_ ( .D(n2222), .CK(wb_clk_o), .Q(rstkram[2])
         );
  DFFQ_X1M_A12TR rstkram_reg_31__14_ ( .D(n2350), .CK(wb_clk_o), .Q(
        rstkram[14]) );
  DFFQ_X1M_A12TR rstkram_reg_31__19_ ( .D(n2574), .CK(wb_clk_o), .Q(
        rstkram[19]) );
  DFFQ_X1M_A12TR rstkram_reg_27__3_ ( .D(n2194), .CK(wb_clk_o), .Q(rstkram[83]) );
  DFFQ_X1M_A12TR rstkram_reg_27__2_ ( .D(n2226), .CK(wb_clk_o), .Q(rstkram[82]) );
  DFFQ_X1M_A12TR rstkram_reg_27__14_ ( .D(n2354), .CK(wb_clk_o), .Q(
        rstkram[94]) );
  DFFQ_X1M_A12TR rstkram_reg_27__19_ ( .D(n2578), .CK(wb_clk_o), .Q(
        rstkram[99]) );
  DFFQ_X1M_A12TR rstkram_reg_23__3_ ( .D(n2198), .CK(wb_clk_o), .Q(
        rstkram[163]) );
  DFFQ_X1M_A12TR rstkram_reg_23__2_ ( .D(n2230), .CK(wb_clk_o), .Q(
        rstkram[162]) );
  DFFQ_X1M_A12TR rstkram_reg_23__14_ ( .D(n2358), .CK(wb_clk_o), .Q(
        rstkram[174]) );
  DFFQ_X1M_A12TR rstkram_reg_23__19_ ( .D(n2582), .CK(wb_clk_o), .Q(
        rstkram[179]) );
  DFFQ_X1M_A12TR rstkram_reg_19__3_ ( .D(n2202), .CK(wb_clk_o), .Q(
        rstkram[243]) );
  DFFQ_X1M_A12TR rstkram_reg_19__2_ ( .D(n2234), .CK(wb_clk_o), .Q(
        rstkram[242]) );
  DFFQ_X1M_A12TR rstkram_reg_19__14_ ( .D(n2362), .CK(wb_clk_o), .Q(
        rstkram[254]) );
  DFFQ_X1M_A12TR rstkram_reg_19__19_ ( .D(n2586), .CK(wb_clk_o), .Q(
        rstkram[259]) );
  DFFQ_X1M_A12TR rstkram_reg_15__3_ ( .D(n2206), .CK(wb_clk_o), .Q(
        rstkram[323]) );
  DFFQ_X1M_A12TR rstkram_reg_15__2_ ( .D(n2238), .CK(wb_clk_o), .Q(
        rstkram[322]) );
  DFFQ_X1M_A12TR rstkram_reg_15__14_ ( .D(n2366), .CK(wb_clk_o), .Q(
        rstkram[334]) );
  DFFQ_X1M_A12TR rstkram_reg_15__19_ ( .D(n2590), .CK(wb_clk_o), .Q(
        rstkram[339]) );
  DFFQ_X1M_A12TR rstkram_reg_11__3_ ( .D(n2210), .CK(wb_clk_o), .Q(
        rstkram[403]) );
  DFFQ_X1M_A12TR rstkram_reg_11__2_ ( .D(n2242), .CK(wb_clk_o), .Q(
        rstkram[402]) );
  DFFQ_X1M_A12TR rstkram_reg_11__14_ ( .D(n2370), .CK(wb_clk_o), .Q(
        rstkram[414]) );
  DFFQ_X1M_A12TR rstkram_reg_11__19_ ( .D(n2594), .CK(wb_clk_o), .Q(
        rstkram[419]) );
  DFFQ_X1M_A12TR rstkram_reg_7__3_ ( .D(n2214), .CK(wb_clk_o), .Q(rstkram[483]) );
  DFFQ_X1M_A12TR rstkram_reg_7__2_ ( .D(n2246), .CK(wb_clk_o), .Q(rstkram[482]) );
  DFFQ_X1M_A12TR rstkram_reg_7__14_ ( .D(n2374), .CK(wb_clk_o), .Q(
        rstkram[494]) );
  DFFQ_X1M_A12TR rstkram_reg_7__19_ ( .D(n2598), .CK(wb_clk_o), .Q(
        rstkram[499]) );
  DFFQ_X1M_A12TR rstkram_reg_3__3_ ( .D(n2218), .CK(wb_clk_o), .Q(rstkram[563]) );
  DFFQ_X1M_A12TR rstkram_reg_3__2_ ( .D(n2250), .CK(wb_clk_o), .Q(rstkram[562]) );
  DFFQ_X1M_A12TR rstkram_reg_3__14_ ( .D(n2378), .CK(wb_clk_o), .Q(
        rstkram[574]) );
  DFFQ_X1M_A12TR rstkram_reg_3__19_ ( .D(n2602), .CK(wb_clk_o), .Q(
        rstkram[579]) );
  DFFQ_X1M_A12TR rstkram_reg_31__7_ ( .D(n2062), .CK(wb_clk_o), .Q(rstkram[7])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__7_ ( .D(n2066), .CK(wb_clk_o), .Q(rstkram[87]) );
  DFFQ_X1M_A12TR rstkram_reg_23__7_ ( .D(n2070), .CK(wb_clk_o), .Q(
        rstkram[167]) );
  DFFQ_X1M_A12TR rstkram_reg_19__7_ ( .D(n2074), .CK(wb_clk_o), .Q(
        rstkram[247]) );
  DFFQ_X1M_A12TR rstkram_reg_15__7_ ( .D(n2078), .CK(wb_clk_o), .Q(
        rstkram[327]) );
  DFFQ_X1M_A12TR rstkram_reg_11__7_ ( .D(n2082), .CK(wb_clk_o), .Q(
        rstkram[407]) );
  DFFQ_X1M_A12TR rstkram_reg_7__7_ ( .D(n2086), .CK(wb_clk_o), .Q(rstkram[487]) );
  DFFQ_X1M_A12TR rstkram_reg_3__7_ ( .D(n2090), .CK(wb_clk_o), .Q(rstkram[567]) );
  DFFQ_X1M_A12TR rstkram_reg_31__5_ ( .D(n2126), .CK(wb_clk_o), .Q(rstkram[5])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__5_ ( .D(n2130), .CK(wb_clk_o), .Q(rstkram[85]) );
  DFFQ_X1M_A12TR rstkram_reg_23__5_ ( .D(n2134), .CK(wb_clk_o), .Q(
        rstkram[165]) );
  DFFQ_X1M_A12TR rstkram_reg_19__5_ ( .D(n2138), .CK(wb_clk_o), .Q(
        rstkram[245]) );
  DFFQ_X1M_A12TR rstkram_reg_15__5_ ( .D(n2142), .CK(wb_clk_o), .Q(
        rstkram[325]) );
  DFFQ_X1M_A12TR rstkram_reg_11__5_ ( .D(n2146), .CK(wb_clk_o), .Q(
        rstkram[405]) );
  DFFQ_X1M_A12TR rstkram_reg_7__5_ ( .D(n2150), .CK(wb_clk_o), .Q(rstkram[485]) );
  DFFQ_X1M_A12TR rstkram_reg_3__5_ ( .D(n2154), .CK(wb_clk_o), .Q(rstkram[565]) );
  DFFQ_X1M_A12TR rstkram_reg_31__1_ ( .D(n2254), .CK(wb_clk_o), .Q(rstkram[1])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__1_ ( .D(n2258), .CK(wb_clk_o), .Q(rstkram[81]) );
  DFFQ_X1M_A12TR rstkram_reg_23__1_ ( .D(n2262), .CK(wb_clk_o), .Q(
        rstkram[161]) );
  DFFQ_X1M_A12TR rstkram_reg_19__1_ ( .D(n2266), .CK(wb_clk_o), .Q(
        rstkram[241]) );
  DFFQ_X1M_A12TR rstkram_reg_15__1_ ( .D(n2270), .CK(wb_clk_o), .Q(
        rstkram[321]) );
  DFFQ_X1M_A12TR rstkram_reg_11__1_ ( .D(n2274), .CK(wb_clk_o), .Q(
        rstkram[401]) );
  DFFQ_X1M_A12TR rstkram_reg_7__1_ ( .D(n2278), .CK(wb_clk_o), .Q(rstkram[481]) );
  DFFQ_X1M_A12TR rstkram_reg_3__1_ ( .D(n2282), .CK(wb_clk_o), .Q(rstkram[561]) );
  DFFQ_X1M_A12TR rstkram_reg_31__4_ ( .D(n2158), .CK(wb_clk_o), .Q(rstkram[4])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__4_ ( .D(n2162), .CK(wb_clk_o), .Q(rstkram[84]) );
  DFFQ_X1M_A12TR rstkram_reg_23__4_ ( .D(n2166), .CK(wb_clk_o), .Q(
        rstkram[164]) );
  DFFQ_X1M_A12TR rstkram_reg_19__4_ ( .D(n2170), .CK(wb_clk_o), .Q(
        rstkram[244]) );
  DFFQ_X1M_A12TR rstkram_reg_15__4_ ( .D(n2174), .CK(wb_clk_o), .Q(
        rstkram[324]) );
  DFFQ_X1M_A12TR rstkram_reg_11__4_ ( .D(n2178), .CK(wb_clk_o), .Q(
        rstkram[404]) );
  DFFQ_X1M_A12TR rstkram_reg_7__4_ ( .D(n2182), .CK(wb_clk_o), .Q(rstkram[484]) );
  DFFQ_X1M_A12TR rstkram_reg_3__4_ ( .D(n2186), .CK(wb_clk_o), .Q(rstkram[564]) );
  DFFQ_X1M_A12TR rstkram_reg_31__13_ ( .D(n2382), .CK(wb_clk_o), .Q(
        rstkram[13]) );
  DFFQ_X1M_A12TR rstkram_reg_27__13_ ( .D(n2386), .CK(wb_clk_o), .Q(
        rstkram[93]) );
  DFFQ_X1M_A12TR rstkram_reg_23__13_ ( .D(n2390), .CK(wb_clk_o), .Q(
        rstkram[173]) );
  DFFQ_X1M_A12TR rstkram_reg_19__13_ ( .D(n2394), .CK(wb_clk_o), .Q(
        rstkram[253]) );
  DFFQ_X1M_A12TR rstkram_reg_15__13_ ( .D(n2398), .CK(wb_clk_o), .Q(
        rstkram[333]) );
  DFFQ_X1M_A12TR rstkram_reg_11__13_ ( .D(n2402), .CK(wb_clk_o), .Q(
        rstkram[413]) );
  DFFQ_X1M_A12TR rstkram_reg_7__13_ ( .D(n2406), .CK(wb_clk_o), .Q(
        rstkram[493]) );
  DFFQ_X1M_A12TR rstkram_reg_3__13_ ( .D(n2410), .CK(wb_clk_o), .Q(
        rstkram[573]) );
  DFFQ_X1M_A12TR rstkram_reg_31__12_ ( .D(n2414), .CK(wb_clk_o), .Q(
        rstkram[12]) );
  DFFQ_X1M_A12TR rstkram_reg_27__12_ ( .D(n2418), .CK(wb_clk_o), .Q(
        rstkram[92]) );
  DFFQ_X1M_A12TR rstkram_reg_23__12_ ( .D(n2422), .CK(wb_clk_o), .Q(
        rstkram[172]) );
  DFFQ_X1M_A12TR rstkram_reg_19__12_ ( .D(n2426), .CK(wb_clk_o), .Q(
        rstkram[252]) );
  DFFQ_X1M_A12TR rstkram_reg_15__12_ ( .D(n2430), .CK(wb_clk_o), .Q(
        rstkram[332]) );
  DFFQ_X1M_A12TR rstkram_reg_11__12_ ( .D(n2434), .CK(wb_clk_o), .Q(
        rstkram[412]) );
  DFFQ_X1M_A12TR rstkram_reg_7__12_ ( .D(n2438), .CK(wb_clk_o), .Q(
        rstkram[492]) );
  DFFQ_X1M_A12TR rstkram_reg_3__12_ ( .D(n2442), .CK(wb_clk_o), .Q(
        rstkram[572]) );
  DFFQ_X1M_A12TR rstkram_reg_31__11_ ( .D(n2446), .CK(wb_clk_o), .Q(
        rstkram[11]) );
  DFFQ_X1M_A12TR rstkram_reg_27__11_ ( .D(n2450), .CK(wb_clk_o), .Q(
        rstkram[91]) );
  DFFQ_X1M_A12TR rstkram_reg_23__11_ ( .D(n2454), .CK(wb_clk_o), .Q(
        rstkram[171]) );
  DFFQ_X1M_A12TR rstkram_reg_19__11_ ( .D(n2458), .CK(wb_clk_o), .Q(
        rstkram[251]) );
  DFFQ_X1M_A12TR rstkram_reg_15__11_ ( .D(n2462), .CK(wb_clk_o), .Q(
        rstkram[331]) );
  DFFQ_X1M_A12TR rstkram_reg_11__11_ ( .D(n2466), .CK(wb_clk_o), .Q(
        rstkram[411]) );
  DFFQ_X1M_A12TR rstkram_reg_7__11_ ( .D(n2470), .CK(wb_clk_o), .Q(
        rstkram[491]) );
  DFFQ_X1M_A12TR rstkram_reg_3__11_ ( .D(n2474), .CK(wb_clk_o), .Q(
        rstkram[571]) );
  DFFQ_X1M_A12TR rstkram_reg_31__10_ ( .D(n2478), .CK(wb_clk_o), .Q(
        rstkram[10]) );
  DFFQ_X1M_A12TR rstkram_reg_27__10_ ( .D(n2482), .CK(wb_clk_o), .Q(
        rstkram[90]) );
  DFFQ_X1M_A12TR rstkram_reg_23__10_ ( .D(n2486), .CK(wb_clk_o), .Q(
        rstkram[170]) );
  DFFQ_X1M_A12TR rstkram_reg_19__10_ ( .D(n2490), .CK(wb_clk_o), .Q(
        rstkram[250]) );
  DFFQ_X1M_A12TR rstkram_reg_15__10_ ( .D(n2494), .CK(wb_clk_o), .Q(
        rstkram[330]) );
  DFFQ_X1M_A12TR rstkram_reg_11__10_ ( .D(n2498), .CK(wb_clk_o), .Q(
        rstkram[410]) );
  DFFQ_X1M_A12TR rstkram_reg_7__10_ ( .D(n2502), .CK(wb_clk_o), .Q(
        rstkram[490]) );
  DFFQ_X1M_A12TR rstkram_reg_3__10_ ( .D(n2506), .CK(wb_clk_o), .Q(
        rstkram[570]) );
  DFFQ_X1M_A12TR rstkram_reg_31__9_ ( .D(n2510), .CK(wb_clk_o), .Q(rstkram[9])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__9_ ( .D(n2514), .CK(wb_clk_o), .Q(rstkram[89]) );
  DFFQ_X1M_A12TR rstkram_reg_23__9_ ( .D(n2518), .CK(wb_clk_o), .Q(
        rstkram[169]) );
  DFFQ_X1M_A12TR rstkram_reg_19__9_ ( .D(n2522), .CK(wb_clk_o), .Q(
        rstkram[249]) );
  DFFQ_X1M_A12TR rstkram_reg_15__9_ ( .D(n2526), .CK(wb_clk_o), .Q(
        rstkram[329]) );
  DFFQ_X1M_A12TR rstkram_reg_11__9_ ( .D(n2530), .CK(wb_clk_o), .Q(
        rstkram[409]) );
  DFFQ_X1M_A12TR rstkram_reg_7__9_ ( .D(n2534), .CK(wb_clk_o), .Q(rstkram[489]) );
  DFFQ_X1M_A12TR rstkram_reg_3__9_ ( .D(n2538), .CK(wb_clk_o), .Q(rstkram[569]) );
  DFFQ_X1M_A12TR rstkram_reg_31__8_ ( .D(n2542), .CK(wb_clk_o), .Q(rstkram[8])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__8_ ( .D(n2546), .CK(wb_clk_o), .Q(rstkram[88]) );
  DFFQ_X1M_A12TR rstkram_reg_23__8_ ( .D(n2550), .CK(wb_clk_o), .Q(
        rstkram[168]) );
  DFFQ_X1M_A12TR rstkram_reg_19__8_ ( .D(n2554), .CK(wb_clk_o), .Q(
        rstkram[248]) );
  DFFQ_X1M_A12TR rstkram_reg_15__8_ ( .D(n2558), .CK(wb_clk_o), .Q(
        rstkram[328]) );
  DFFQ_X1M_A12TR rstkram_reg_11__8_ ( .D(n2562), .CK(wb_clk_o), .Q(
        rstkram[408]) );
  DFFQ_X1M_A12TR rstkram_reg_7__8_ ( .D(n2566), .CK(wb_clk_o), .Q(rstkram[488]) );
  DFFQ_X1M_A12TR rstkram_reg_3__8_ ( .D(n2570), .CK(wb_clk_o), .Q(rstkram[568]) );
  DFFQ_X1M_A12TR rstkram_reg_31__6_ ( .D(n2094), .CK(wb_clk_o), .Q(rstkram[6])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__6_ ( .D(n2098), .CK(wb_clk_o), .Q(rstkram[86]) );
  DFFQ_X1M_A12TR rstkram_reg_23__6_ ( .D(n2102), .CK(wb_clk_o), .Q(
        rstkram[166]) );
  DFFQ_X1M_A12TR rstkram_reg_19__6_ ( .D(n2106), .CK(wb_clk_o), .Q(
        rstkram[246]) );
  DFFQ_X1M_A12TR rstkram_reg_15__6_ ( .D(n2110), .CK(wb_clk_o), .Q(
        rstkram[326]) );
  DFFQ_X1M_A12TR rstkram_reg_11__6_ ( .D(n2114), .CK(wb_clk_o), .Q(
        rstkram[406]) );
  DFFQ_X1M_A12TR rstkram_reg_7__6_ ( .D(n2118), .CK(wb_clk_o), .Q(rstkram[486]) );
  DFFQ_X1M_A12TR rstkram_reg_3__6_ ( .D(n2122), .CK(wb_clk_o), .Q(rstkram[566]) );
  DFFQ_X1M_A12TR rstkram_reg_31__15_ ( .D(n2318), .CK(wb_clk_o), .Q(
        rstkram[15]) );
  DFFQ_X1M_A12TR rstkram_reg_27__15_ ( .D(n2322), .CK(wb_clk_o), .Q(
        rstkram[95]) );
  DFFQ_X1M_A12TR rstkram_reg_23__15_ ( .D(n2326), .CK(wb_clk_o), .Q(
        rstkram[175]) );
  DFFQ_X1M_A12TR rstkram_reg_19__15_ ( .D(n2330), .CK(wb_clk_o), .Q(
        rstkram[255]) );
  DFFQ_X1M_A12TR rstkram_reg_15__15_ ( .D(n2334), .CK(wb_clk_o), .Q(
        rstkram[335]) );
  DFFQ_X1M_A12TR rstkram_reg_11__15_ ( .D(n2338), .CK(wb_clk_o), .Q(
        rstkram[415]) );
  DFFQ_X1M_A12TR rstkram_reg_7__15_ ( .D(n2342), .CK(wb_clk_o), .Q(
        rstkram[495]) );
  DFFQ_X1M_A12TR rstkram_reg_3__15_ ( .D(n2346), .CK(wb_clk_o), .Q(
        rstkram[575]) );
  DFFQ_X1M_A12TR rstkram_reg_31__16_ ( .D(n2670), .CK(wb_clk_o), .Q(
        rstkram[16]) );
  DFFQ_X1M_A12TR rstkram_reg_27__16_ ( .D(n2674), .CK(wb_clk_o), .Q(
        rstkram[96]) );
  DFFQ_X1M_A12TR rstkram_reg_23__16_ ( .D(n2678), .CK(wb_clk_o), .Q(
        rstkram[176]) );
  DFFQ_X1M_A12TR rstkram_reg_19__16_ ( .D(n2682), .CK(wb_clk_o), .Q(
        rstkram[256]) );
  DFFQ_X1M_A12TR rstkram_reg_15__16_ ( .D(n2686), .CK(wb_clk_o), .Q(
        rstkram[336]) );
  DFFQ_X1M_A12TR rstkram_reg_11__16_ ( .D(n2690), .CK(wb_clk_o), .Q(
        rstkram[416]) );
  DFFQ_X1M_A12TR rstkram_reg_7__16_ ( .D(n2694), .CK(wb_clk_o), .Q(
        rstkram[496]) );
  DFFQ_X1M_A12TR rstkram_reg_3__16_ ( .D(n2698), .CK(wb_clk_o), .Q(
        rstkram[576]) );
  DFFQ_X1M_A12TR rstkram_reg_31__17_ ( .D(n2638), .CK(wb_clk_o), .Q(
        rstkram[17]) );
  DFFQ_X1M_A12TR rstkram_reg_27__17_ ( .D(n2642), .CK(wb_clk_o), .Q(
        rstkram[97]) );
  DFFQ_X1M_A12TR rstkram_reg_23__17_ ( .D(n2646), .CK(wb_clk_o), .Q(
        rstkram[177]) );
  DFFQ_X1M_A12TR rstkram_reg_19__17_ ( .D(n2650), .CK(wb_clk_o), .Q(
        rstkram[257]) );
  DFFQ_X1M_A12TR rstkram_reg_15__17_ ( .D(n2654), .CK(wb_clk_o), .Q(
        rstkram[337]) );
  DFFQ_X1M_A12TR rstkram_reg_11__17_ ( .D(n2658), .CK(wb_clk_o), .Q(
        rstkram[417]) );
  DFFQ_X1M_A12TR rstkram_reg_7__17_ ( .D(n2662), .CK(wb_clk_o), .Q(
        rstkram[497]) );
  DFFQ_X1M_A12TR rstkram_reg_3__17_ ( .D(n2666), .CK(wb_clk_o), .Q(
        rstkram[577]) );
  DFFQ_X1M_A12TR rstkram_reg_31__18_ ( .D(n2606), .CK(wb_clk_o), .Q(
        rstkram[18]) );
  DFFQ_X1M_A12TR rstkram_reg_27__18_ ( .D(n2610), .CK(wb_clk_o), .Q(
        rstkram[98]) );
  DFFQ_X1M_A12TR rstkram_reg_23__18_ ( .D(n2614), .CK(wb_clk_o), .Q(
        rstkram[178]) );
  DFFQ_X1M_A12TR rstkram_reg_19__18_ ( .D(n2618), .CK(wb_clk_o), .Q(
        rstkram[258]) );
  DFFQ_X1M_A12TR rstkram_reg_15__18_ ( .D(n2622), .CK(wb_clk_o), .Q(
        rstkram[338]) );
  DFFQ_X1M_A12TR rstkram_reg_11__18_ ( .D(n2626), .CK(wb_clk_o), .Q(
        rstkram[418]) );
  DFFQ_X1M_A12TR rstkram_reg_7__18_ ( .D(n2630), .CK(wb_clk_o), .Q(
        rstkram[498]) );
  DFFQ_X1M_A12TR rstkram_reg_3__18_ ( .D(n2634), .CK(wb_clk_o), .Q(
        rstkram[578]) );
  DFFQ_X1M_A12TR rstkram_reg_31__0_ ( .D(n2286), .CK(wb_clk_o), .Q(rstkram[0])
         );
  DFFQ_X1M_A12TR rstkram_reg_27__0_ ( .D(n2290), .CK(wb_clk_o), .Q(rstkram[80]) );
  DFFQ_X1M_A12TR rstkram_reg_23__0_ ( .D(n2294), .CK(wb_clk_o), .Q(
        rstkram[160]) );
  DFFQ_X1M_A12TR rstkram_reg_19__0_ ( .D(n2298), .CK(wb_clk_o), .Q(
        rstkram[240]) );
  DFFQ_X1M_A12TR rstkram_reg_15__0_ ( .D(n2302), .CK(wb_clk_o), .Q(
        rstkram[320]) );
  DFFQ_X1M_A12TR rstkram_reg_11__0_ ( .D(n2306), .CK(wb_clk_o), .Q(
        rstkram[400]) );
  DFFQ_X1M_A12TR rstkram_reg_7__0_ ( .D(n2310), .CK(wb_clk_o), .Q(rstkram[480]) );
  DFFQ_X1M_A12TR rstkram_reg_3__0_ ( .D(n2314), .CK(wb_clk_o), .Q(rstkram[560]) );
  DFFQ_X1M_A12TR rstkram_reg_29__3_ ( .D(n2192), .CK(wb_clk_o), .Q(rstkram[43]) );
  DFFQ_X1M_A12TR rstkram_reg_29__2_ ( .D(n2224), .CK(wb_clk_o), .Q(rstkram[42]) );
  DFFQ_X1M_A12TR rstkram_reg_29__14_ ( .D(n2352), .CK(wb_clk_o), .Q(
        rstkram[54]) );
  DFFQ_X1M_A12TR rstkram_reg_29__19_ ( .D(n2576), .CK(wb_clk_o), .Q(
        rstkram[59]) );
  DFFQ_X1M_A12TR rstkram_reg_25__3_ ( .D(n2196), .CK(wb_clk_o), .Q(
        rstkram[123]) );
  DFFQ_X1M_A12TR rstkram_reg_25__2_ ( .D(n2228), .CK(wb_clk_o), .Q(
        rstkram[122]) );
  DFFQ_X1M_A12TR rstkram_reg_25__14_ ( .D(n2356), .CK(wb_clk_o), .Q(
        rstkram[134]) );
  DFFQ_X1M_A12TR rstkram_reg_25__19_ ( .D(n2580), .CK(wb_clk_o), .Q(
        rstkram[139]) );
  DFFQ_X1M_A12TR rstkram_reg_21__3_ ( .D(n2200), .CK(wb_clk_o), .Q(
        rstkram[203]) );
  DFFQ_X1M_A12TR rstkram_reg_21__2_ ( .D(n2232), .CK(wb_clk_o), .Q(
        rstkram[202]) );
  DFFQ_X1M_A12TR rstkram_reg_21__14_ ( .D(n2360), .CK(wb_clk_o), .Q(
        rstkram[214]) );
  DFFQ_X1M_A12TR rstkram_reg_21__19_ ( .D(n2584), .CK(wb_clk_o), .Q(
        rstkram[219]) );
  DFFQ_X1M_A12TR rstkram_reg_17__3_ ( .D(n2204), .CK(wb_clk_o), .Q(
        rstkram[283]) );
  DFFQ_X1M_A12TR rstkram_reg_17__2_ ( .D(n2236), .CK(wb_clk_o), .Q(
        rstkram[282]) );
  DFFQ_X1M_A12TR rstkram_reg_17__14_ ( .D(n2364), .CK(wb_clk_o), .Q(
        rstkram[294]) );
  DFFQ_X1M_A12TR rstkram_reg_17__19_ ( .D(n2588), .CK(wb_clk_o), .Q(
        rstkram[299]) );
  DFFQ_X1M_A12TR rstkram_reg_13__3_ ( .D(n2208), .CK(wb_clk_o), .Q(
        rstkram[363]) );
  DFFQ_X1M_A12TR rstkram_reg_13__2_ ( .D(n2240), .CK(wb_clk_o), .Q(
        rstkram[362]) );
  DFFQ_X1M_A12TR rstkram_reg_13__14_ ( .D(n2368), .CK(wb_clk_o), .Q(
        rstkram[374]) );
  DFFQ_X1M_A12TR rstkram_reg_13__19_ ( .D(n2592), .CK(wb_clk_o), .Q(
        rstkram[379]) );
  DFFQ_X1M_A12TR rstkram_reg_9__3_ ( .D(n2212), .CK(wb_clk_o), .Q(rstkram[443]) );
  DFFQ_X1M_A12TR rstkram_reg_9__2_ ( .D(n2244), .CK(wb_clk_o), .Q(rstkram[442]) );
  DFFQ_X1M_A12TR rstkram_reg_9__14_ ( .D(n2372), .CK(wb_clk_o), .Q(
        rstkram[454]) );
  DFFQ_X1M_A12TR rstkram_reg_9__19_ ( .D(n2596), .CK(wb_clk_o), .Q(
        rstkram[459]) );
  DFFQ_X1M_A12TR rstkram_reg_5__3_ ( .D(n2216), .CK(wb_clk_o), .Q(rstkram[523]) );
  DFFQ_X1M_A12TR rstkram_reg_5__2_ ( .D(n2248), .CK(wb_clk_o), .Q(rstkram[522]) );
  DFFQ_X1M_A12TR rstkram_reg_5__14_ ( .D(n2376), .CK(wb_clk_o), .Q(
        rstkram[534]) );
  DFFQ_X1M_A12TR rstkram_reg_5__19_ ( .D(n2600), .CK(wb_clk_o), .Q(
        rstkram[539]) );
  DFFQ_X1M_A12TR rstkram_reg_1__3_ ( .D(n2220), .CK(wb_clk_o), .Q(rstkram[603]) );
  DFFQ_X1M_A12TR rstkram_reg_1__2_ ( .D(n2252), .CK(wb_clk_o), .Q(rstkram[602]) );
  DFFQ_X1M_A12TR rstkram_reg_1__14_ ( .D(n2380), .CK(wb_clk_o), .Q(
        rstkram[614]) );
  DFFQ_X1M_A12TR rstkram_reg_1__19_ ( .D(n2604), .CK(wb_clk_o), .Q(
        rstkram[619]) );
  DFFQ_X1M_A12TR rstkram_reg_29__7_ ( .D(n2064), .CK(wb_clk_o), .Q(rstkram[47]) );
  DFFQ_X1M_A12TR rstkram_reg_25__7_ ( .D(n2068), .CK(wb_clk_o), .Q(
        rstkram[127]) );
  DFFQ_X1M_A12TR rstkram_reg_21__7_ ( .D(n2072), .CK(wb_clk_o), .Q(
        rstkram[207]) );
  DFFQ_X1M_A12TR rstkram_reg_17__7_ ( .D(n2076), .CK(wb_clk_o), .Q(
        rstkram[287]) );
  DFFQ_X1M_A12TR rstkram_reg_13__7_ ( .D(n2080), .CK(wb_clk_o), .Q(
        rstkram[367]) );
  DFFQ_X1M_A12TR rstkram_reg_9__7_ ( .D(n2084), .CK(wb_clk_o), .Q(rstkram[447]) );
  DFFQ_X1M_A12TR rstkram_reg_5__7_ ( .D(n2088), .CK(wb_clk_o), .Q(rstkram[527]) );
  DFFQ_X1M_A12TR rstkram_reg_1__7_ ( .D(n2092), .CK(wb_clk_o), .Q(rstkram[607]) );
  DFFQ_X1M_A12TR rstkram_reg_29__5_ ( .D(n2128), .CK(wb_clk_o), .Q(rstkram[45]) );
  DFFQ_X1M_A12TR rstkram_reg_25__5_ ( .D(n2132), .CK(wb_clk_o), .Q(
        rstkram[125]) );
  DFFQ_X1M_A12TR rstkram_reg_21__5_ ( .D(n2136), .CK(wb_clk_o), .Q(
        rstkram[205]) );
  DFFQ_X1M_A12TR rstkram_reg_17__5_ ( .D(n2140), .CK(wb_clk_o), .Q(
        rstkram[285]) );
  DFFQ_X1M_A12TR rstkram_reg_13__5_ ( .D(n2144), .CK(wb_clk_o), .Q(
        rstkram[365]) );
  DFFQ_X1M_A12TR rstkram_reg_9__5_ ( .D(n2148), .CK(wb_clk_o), .Q(rstkram[445]) );
  DFFQ_X1M_A12TR rstkram_reg_5__5_ ( .D(n2152), .CK(wb_clk_o), .Q(rstkram[525]) );
  DFFQ_X1M_A12TR rstkram_reg_1__5_ ( .D(n2156), .CK(wb_clk_o), .Q(rstkram[605]) );
  DFFQ_X1M_A12TR rstkram_reg_29__1_ ( .D(n2256), .CK(wb_clk_o), .Q(rstkram[41]) );
  DFFQ_X1M_A12TR rstkram_reg_25__1_ ( .D(n2260), .CK(wb_clk_o), .Q(
        rstkram[121]) );
  DFFQ_X1M_A12TR rstkram_reg_21__1_ ( .D(n2264), .CK(wb_clk_o), .Q(
        rstkram[201]) );
  DFFQ_X1M_A12TR rstkram_reg_17__1_ ( .D(n2268), .CK(wb_clk_o), .Q(
        rstkram[281]) );
  DFFQ_X1M_A12TR rstkram_reg_13__1_ ( .D(n2272), .CK(wb_clk_o), .Q(
        rstkram[361]) );
  DFFQ_X1M_A12TR rstkram_reg_9__1_ ( .D(n2276), .CK(wb_clk_o), .Q(rstkram[441]) );
  DFFQ_X1M_A12TR rstkram_reg_5__1_ ( .D(n2280), .CK(wb_clk_o), .Q(rstkram[521]) );
  DFFQ_X1M_A12TR rstkram_reg_1__1_ ( .D(n2284), .CK(wb_clk_o), .Q(rstkram[601]) );
  DFFQ_X1M_A12TR rstkram_reg_29__4_ ( .D(n2160), .CK(wb_clk_o), .Q(rstkram[44]) );
  DFFQ_X1M_A12TR rstkram_reg_25__4_ ( .D(n2164), .CK(wb_clk_o), .Q(
        rstkram[124]) );
  DFFQ_X1M_A12TR rstkram_reg_21__4_ ( .D(n2168), .CK(wb_clk_o), .Q(
        rstkram[204]) );
  DFFQ_X1M_A12TR rstkram_reg_17__4_ ( .D(n2172), .CK(wb_clk_o), .Q(
        rstkram[284]) );
  DFFQ_X1M_A12TR rstkram_reg_13__4_ ( .D(n2176), .CK(wb_clk_o), .Q(
        rstkram[364]) );
  DFFQ_X1M_A12TR rstkram_reg_9__4_ ( .D(n2180), .CK(wb_clk_o), .Q(rstkram[444]) );
  DFFQ_X1M_A12TR rstkram_reg_5__4_ ( .D(n2184), .CK(wb_clk_o), .Q(rstkram[524]) );
  DFFQ_X1M_A12TR rstkram_reg_1__4_ ( .D(n2188), .CK(wb_clk_o), .Q(rstkram[604]) );
  DFFQ_X1M_A12TR rstkram_reg_29__13_ ( .D(n2384), .CK(wb_clk_o), .Q(
        rstkram[53]) );
  DFFQ_X1M_A12TR rstkram_reg_25__13_ ( .D(n2388), .CK(wb_clk_o), .Q(
        rstkram[133]) );
  DFFQ_X1M_A12TR rstkram_reg_21__13_ ( .D(n2392), .CK(wb_clk_o), .Q(
        rstkram[213]) );
  DFFQ_X1M_A12TR rstkram_reg_17__13_ ( .D(n2396), .CK(wb_clk_o), .Q(
        rstkram[293]) );
  DFFQ_X1M_A12TR rstkram_reg_13__13_ ( .D(n2400), .CK(wb_clk_o), .Q(
        rstkram[373]) );
  DFFQ_X1M_A12TR rstkram_reg_9__13_ ( .D(n2404), .CK(wb_clk_o), .Q(
        rstkram[453]) );
  DFFQ_X1M_A12TR rstkram_reg_5__13_ ( .D(n2408), .CK(wb_clk_o), .Q(
        rstkram[533]) );
  DFFQ_X1M_A12TR rstkram_reg_1__13_ ( .D(n2412), .CK(wb_clk_o), .Q(
        rstkram[613]) );
  DFFQ_X1M_A12TR rstkram_reg_29__12_ ( .D(n2416), .CK(wb_clk_o), .Q(
        rstkram[52]) );
  DFFQ_X1M_A12TR rstkram_reg_25__12_ ( .D(n2420), .CK(wb_clk_o), .Q(
        rstkram[132]) );
  DFFQ_X1M_A12TR rstkram_reg_21__12_ ( .D(n2424), .CK(wb_clk_o), .Q(
        rstkram[212]) );
  DFFQ_X1M_A12TR rstkram_reg_17__12_ ( .D(n2428), .CK(wb_clk_o), .Q(
        rstkram[292]) );
  DFFQ_X1M_A12TR rstkram_reg_13__12_ ( .D(n2432), .CK(wb_clk_o), .Q(
        rstkram[372]) );
  DFFQ_X1M_A12TR rstkram_reg_9__12_ ( .D(n2436), .CK(wb_clk_o), .Q(
        rstkram[452]) );
  DFFQ_X1M_A12TR rstkram_reg_5__12_ ( .D(n2440), .CK(wb_clk_o), .Q(
        rstkram[532]) );
  DFFQ_X1M_A12TR rstkram_reg_1__12_ ( .D(n2444), .CK(wb_clk_o), .Q(
        rstkram[612]) );
  DFFQ_X1M_A12TR rstkram_reg_29__11_ ( .D(n2448), .CK(wb_clk_o), .Q(
        rstkram[51]) );
  DFFQ_X1M_A12TR rstkram_reg_25__11_ ( .D(n2452), .CK(wb_clk_o), .Q(
        rstkram[131]) );
  DFFQ_X1M_A12TR rstkram_reg_21__11_ ( .D(n2456), .CK(wb_clk_o), .Q(
        rstkram[211]) );
  DFFQ_X1M_A12TR rstkram_reg_17__11_ ( .D(n2460), .CK(wb_clk_o), .Q(
        rstkram[291]) );
  DFFQ_X1M_A12TR rstkram_reg_13__11_ ( .D(n2464), .CK(wb_clk_o), .Q(
        rstkram[371]) );
  DFFQ_X1M_A12TR rstkram_reg_9__11_ ( .D(n2468), .CK(wb_clk_o), .Q(
        rstkram[451]) );
  DFFQ_X1M_A12TR rstkram_reg_5__11_ ( .D(n2472), .CK(wb_clk_o), .Q(
        rstkram[531]) );
  DFFQ_X1M_A12TR rstkram_reg_1__11_ ( .D(n2476), .CK(wb_clk_o), .Q(
        rstkram[611]) );
  DFFQ_X1M_A12TR rstkram_reg_29__10_ ( .D(n2480), .CK(wb_clk_o), .Q(
        rstkram[50]) );
  DFFQ_X1M_A12TR rstkram_reg_25__10_ ( .D(n2484), .CK(wb_clk_o), .Q(
        rstkram[130]) );
  DFFQ_X1M_A12TR rstkram_reg_21__10_ ( .D(n2488), .CK(wb_clk_o), .Q(
        rstkram[210]) );
  DFFQ_X1M_A12TR rstkram_reg_17__10_ ( .D(n2492), .CK(wb_clk_o), .Q(
        rstkram[290]) );
  DFFQ_X1M_A12TR rstkram_reg_13__10_ ( .D(n2496), .CK(wb_clk_o), .Q(
        rstkram[370]) );
  DFFQ_X1M_A12TR rstkram_reg_9__10_ ( .D(n2500), .CK(wb_clk_o), .Q(
        rstkram[450]) );
  DFFQ_X1M_A12TR rstkram_reg_5__10_ ( .D(n2504), .CK(wb_clk_o), .Q(
        rstkram[530]) );
  DFFQ_X1M_A12TR rstkram_reg_1__10_ ( .D(n2508), .CK(wb_clk_o), .Q(
        rstkram[610]) );
  DFFQ_X1M_A12TR rstkram_reg_29__9_ ( .D(n2512), .CK(wb_clk_o), .Q(rstkram[49]) );
  DFFQ_X1M_A12TR rstkram_reg_25__9_ ( .D(n2516), .CK(wb_clk_o), .Q(
        rstkram[129]) );
  DFFQ_X1M_A12TR rstkram_reg_21__9_ ( .D(n2520), .CK(wb_clk_o), .Q(
        rstkram[209]) );
  DFFQ_X1M_A12TR rstkram_reg_17__9_ ( .D(n2524), .CK(wb_clk_o), .Q(
        rstkram[289]) );
  DFFQ_X1M_A12TR rstkram_reg_13__9_ ( .D(n2528), .CK(wb_clk_o), .Q(
        rstkram[369]) );
  DFFQ_X1M_A12TR rstkram_reg_9__9_ ( .D(n2532), .CK(wb_clk_o), .Q(rstkram[449]) );
  DFFQ_X1M_A12TR rstkram_reg_5__9_ ( .D(n2536), .CK(wb_clk_o), .Q(rstkram[529]) );
  DFFQ_X1M_A12TR rstkram_reg_1__9_ ( .D(n2540), .CK(wb_clk_o), .Q(rstkram[609]) );
  DFFQ_X1M_A12TR rstkram_reg_29__8_ ( .D(n2544), .CK(wb_clk_o), .Q(rstkram[48]) );
  DFFQ_X1M_A12TR rstkram_reg_25__8_ ( .D(n2548), .CK(wb_clk_o), .Q(
        rstkram[128]) );
  DFFQ_X1M_A12TR rstkram_reg_21__8_ ( .D(n2552), .CK(wb_clk_o), .Q(
        rstkram[208]) );
  DFFQ_X1M_A12TR rstkram_reg_17__8_ ( .D(n2556), .CK(wb_clk_o), .Q(
        rstkram[288]) );
  DFFQ_X1M_A12TR rstkram_reg_13__8_ ( .D(n2560), .CK(wb_clk_o), .Q(
        rstkram[368]) );
  DFFQ_X1M_A12TR rstkram_reg_9__8_ ( .D(n2564), .CK(wb_clk_o), .Q(rstkram[448]) );
  DFFQ_X1M_A12TR rstkram_reg_5__8_ ( .D(n2568), .CK(wb_clk_o), .Q(rstkram[528]) );
  DFFQ_X1M_A12TR rstkram_reg_1__8_ ( .D(n2572), .CK(wb_clk_o), .Q(rstkram[608]) );
  DFFQ_X1M_A12TR rstkram_reg_29__6_ ( .D(n2096), .CK(wb_clk_o), .Q(rstkram[46]) );
  DFFQ_X1M_A12TR rstkram_reg_25__6_ ( .D(n2100), .CK(wb_clk_o), .Q(
        rstkram[126]) );
  DFFQ_X1M_A12TR rstkram_reg_21__6_ ( .D(n2104), .CK(wb_clk_o), .Q(
        rstkram[206]) );
  DFFQ_X1M_A12TR rstkram_reg_17__6_ ( .D(n2108), .CK(wb_clk_o), .Q(
        rstkram[286]) );
  DFFQ_X1M_A12TR rstkram_reg_13__6_ ( .D(n2112), .CK(wb_clk_o), .Q(
        rstkram[366]) );
  DFFQ_X1M_A12TR rstkram_reg_9__6_ ( .D(n2116), .CK(wb_clk_o), .Q(rstkram[446]) );
  DFFQ_X1M_A12TR rstkram_reg_5__6_ ( .D(n2120), .CK(wb_clk_o), .Q(rstkram[526]) );
  DFFQ_X1M_A12TR rstkram_reg_1__6_ ( .D(n2124), .CK(wb_clk_o), .Q(rstkram[606]) );
  DFFQ_X1M_A12TR rstkram_reg_29__15_ ( .D(n2320), .CK(wb_clk_o), .Q(
        rstkram[55]) );
  DFFQ_X1M_A12TR rstkram_reg_25__15_ ( .D(n2324), .CK(wb_clk_o), .Q(
        rstkram[135]) );
  DFFQ_X1M_A12TR rstkram_reg_21__15_ ( .D(n2328), .CK(wb_clk_o), .Q(
        rstkram[215]) );
  DFFQ_X1M_A12TR rstkram_reg_17__15_ ( .D(n2332), .CK(wb_clk_o), .Q(
        rstkram[295]) );
  DFFQ_X1M_A12TR rstkram_reg_13__15_ ( .D(n2336), .CK(wb_clk_o), .Q(
        rstkram[375]) );
  DFFQ_X1M_A12TR rstkram_reg_9__15_ ( .D(n2340), .CK(wb_clk_o), .Q(
        rstkram[455]) );
  DFFQ_X1M_A12TR rstkram_reg_5__15_ ( .D(n2344), .CK(wb_clk_o), .Q(
        rstkram[535]) );
  DFFQ_X1M_A12TR rstkram_reg_1__15_ ( .D(n2348), .CK(wb_clk_o), .Q(
        rstkram[615]) );
  DFFQ_X1M_A12TR rstkram_reg_29__16_ ( .D(n2672), .CK(wb_clk_o), .Q(
        rstkram[56]) );
  DFFQ_X1M_A12TR rstkram_reg_25__16_ ( .D(n2676), .CK(wb_clk_o), .Q(
        rstkram[136]) );
  DFFQ_X1M_A12TR rstkram_reg_21__16_ ( .D(n2680), .CK(wb_clk_o), .Q(
        rstkram[216]) );
  DFFQ_X1M_A12TR rstkram_reg_17__16_ ( .D(n2684), .CK(wb_clk_o), .Q(
        rstkram[296]) );
  DFFQ_X1M_A12TR rstkram_reg_13__16_ ( .D(n2688), .CK(wb_clk_o), .Q(
        rstkram[376]) );
  DFFQ_X1M_A12TR rstkram_reg_9__16_ ( .D(n2692), .CK(wb_clk_o), .Q(
        rstkram[456]) );
  DFFQ_X1M_A12TR rstkram_reg_5__16_ ( .D(n2696), .CK(wb_clk_o), .Q(
        rstkram[536]) );
  DFFQ_X1M_A12TR rstkram_reg_1__16_ ( .D(n2700), .CK(wb_clk_o), .Q(
        rstkram[616]) );
  DFFQ_X1M_A12TR rstkram_reg_29__17_ ( .D(n2640), .CK(wb_clk_o), .Q(
        rstkram[57]) );
  DFFQ_X1M_A12TR rstkram_reg_25__17_ ( .D(n2644), .CK(wb_clk_o), .Q(
        rstkram[137]) );
  DFFQ_X1M_A12TR rstkram_reg_21__17_ ( .D(n2648), .CK(wb_clk_o), .Q(
        rstkram[217]) );
  DFFQ_X1M_A12TR rstkram_reg_17__17_ ( .D(n2652), .CK(wb_clk_o), .Q(
        rstkram[297]) );
  DFFQ_X1M_A12TR rstkram_reg_13__17_ ( .D(n2656), .CK(wb_clk_o), .Q(
        rstkram[377]) );
  DFFQ_X1M_A12TR rstkram_reg_9__17_ ( .D(n2660), .CK(wb_clk_o), .Q(
        rstkram[457]) );
  DFFQ_X1M_A12TR rstkram_reg_5__17_ ( .D(n2664), .CK(wb_clk_o), .Q(
        rstkram[537]) );
  DFFQ_X1M_A12TR rstkram_reg_1__17_ ( .D(n2668), .CK(wb_clk_o), .Q(
        rstkram[617]) );
  DFFQ_X1M_A12TR rstkram_reg_29__18_ ( .D(n2608), .CK(wb_clk_o), .Q(
        rstkram[58]) );
  DFFQ_X1M_A12TR rstkram_reg_25__18_ ( .D(n2612), .CK(wb_clk_o), .Q(
        rstkram[138]) );
  DFFQ_X1M_A12TR rstkram_reg_21__18_ ( .D(n2616), .CK(wb_clk_o), .Q(
        rstkram[218]) );
  DFFQ_X1M_A12TR rstkram_reg_17__18_ ( .D(n2620), .CK(wb_clk_o), .Q(
        rstkram[298]) );
  DFFQ_X1M_A12TR rstkram_reg_13__18_ ( .D(n2624), .CK(wb_clk_o), .Q(
        rstkram[378]) );
  DFFQ_X1M_A12TR rstkram_reg_9__18_ ( .D(n2628), .CK(wb_clk_o), .Q(
        rstkram[458]) );
  DFFQ_X1M_A12TR rstkram_reg_5__18_ ( .D(n2632), .CK(wb_clk_o), .Q(
        rstkram[538]) );
  DFFQ_X1M_A12TR rstkram_reg_1__18_ ( .D(n2636), .CK(wb_clk_o), .Q(
        rstkram[618]) );
  DFFQ_X1M_A12TR rstkram_reg_29__0_ ( .D(n2288), .CK(wb_clk_o), .Q(rstkram[40]) );
  DFFQ_X1M_A12TR rstkram_reg_25__0_ ( .D(n2292), .CK(wb_clk_o), .Q(
        rstkram[120]) );
  DFFQ_X1M_A12TR rstkram_reg_21__0_ ( .D(n2296), .CK(wb_clk_o), .Q(
        rstkram[200]) );
  DFFQ_X1M_A12TR rstkram_reg_17__0_ ( .D(n2300), .CK(wb_clk_o), .Q(
        rstkram[280]) );
  DFFQ_X1M_A12TR rstkram_reg_13__0_ ( .D(n2304), .CK(wb_clk_o), .Q(
        rstkram[360]) );
  DFFQ_X1M_A12TR rstkram_reg_9__0_ ( .D(n2308), .CK(wb_clk_o), .Q(rstkram[440]) );
  DFFQ_X1M_A12TR rstkram_reg_5__0_ ( .D(n2312), .CK(wb_clk_o), .Q(rstkram[520]) );
  DFFQ_X1M_A12TR rstkram_reg_1__0_ ( .D(n2316), .CK(wb_clk_o), .Q(rstkram[600]) );
  DFFQ_X1M_A12TR rstkram_reg_28__3_ ( .D(n2193), .CK(wb_clk_o), .Q(rstkram[63]) );
  DFFQ_X1M_A12TR rstkram_reg_28__2_ ( .D(n2225), .CK(wb_clk_o), .Q(rstkram[62]) );
  DFFQ_X1M_A12TR rstkram_reg_28__14_ ( .D(n2353), .CK(wb_clk_o), .Q(
        rstkram[74]) );
  DFFQ_X1M_A12TR rstkram_reg_28__19_ ( .D(n2577), .CK(wb_clk_o), .Q(
        rstkram[79]) );
  DFFQ_X1M_A12TR rstkram_reg_24__3_ ( .D(n2197), .CK(wb_clk_o), .Q(
        rstkram[143]) );
  DFFQ_X1M_A12TR rstkram_reg_24__2_ ( .D(n2229), .CK(wb_clk_o), .Q(
        rstkram[142]) );
  DFFQ_X1M_A12TR rstkram_reg_24__14_ ( .D(n2357), .CK(wb_clk_o), .Q(
        rstkram[154]) );
  DFFQ_X1M_A12TR rstkram_reg_24__19_ ( .D(n2581), .CK(wb_clk_o), .Q(
        rstkram[159]) );
  DFFQ_X1M_A12TR rstkram_reg_20__3_ ( .D(n2201), .CK(wb_clk_o), .Q(
        rstkram[223]) );
  DFFQ_X1M_A12TR rstkram_reg_20__2_ ( .D(n2233), .CK(wb_clk_o), .Q(
        rstkram[222]) );
  DFFQ_X1M_A12TR rstkram_reg_20__14_ ( .D(n2361), .CK(wb_clk_o), .Q(
        rstkram[234]) );
  DFFQ_X1M_A12TR rstkram_reg_20__19_ ( .D(n2585), .CK(wb_clk_o), .Q(
        rstkram[239]) );
  DFFQ_X1M_A12TR rstkram_reg_16__3_ ( .D(n2205), .CK(wb_clk_o), .Q(
        rstkram[303]) );
  DFFQ_X1M_A12TR rstkram_reg_16__2_ ( .D(n2237), .CK(wb_clk_o), .Q(
        rstkram[302]) );
  DFFQ_X1M_A12TR rstkram_reg_16__14_ ( .D(n2365), .CK(wb_clk_o), .Q(
        rstkram[314]) );
  DFFQ_X1M_A12TR rstkram_reg_16__19_ ( .D(n2589), .CK(wb_clk_o), .Q(
        rstkram[319]) );
  DFFQ_X1M_A12TR rstkram_reg_12__3_ ( .D(n2209), .CK(wb_clk_o), .Q(
        rstkram[383]) );
  DFFQ_X1M_A12TR rstkram_reg_12__2_ ( .D(n2241), .CK(wb_clk_o), .Q(
        rstkram[382]) );
  DFFQ_X1M_A12TR rstkram_reg_12__14_ ( .D(n2369), .CK(wb_clk_o), .Q(
        rstkram[394]) );
  DFFQ_X1M_A12TR rstkram_reg_12__19_ ( .D(n2593), .CK(wb_clk_o), .Q(
        rstkram[399]) );
  DFFQ_X1M_A12TR rstkram_reg_8__3_ ( .D(n2213), .CK(wb_clk_o), .Q(rstkram[463]) );
  DFFQ_X1M_A12TR rstkram_reg_8__2_ ( .D(n2245), .CK(wb_clk_o), .Q(rstkram[462]) );
  DFFQ_X1M_A12TR rstkram_reg_8__14_ ( .D(n2373), .CK(wb_clk_o), .Q(
        rstkram[474]) );
  DFFQ_X1M_A12TR rstkram_reg_8__19_ ( .D(n2597), .CK(wb_clk_o), .Q(
        rstkram[479]) );
  DFFQ_X1M_A12TR rstkram_reg_4__3_ ( .D(n2217), .CK(wb_clk_o), .Q(rstkram[543]) );
  DFFQ_X1M_A12TR rstkram_reg_4__2_ ( .D(n2249), .CK(wb_clk_o), .Q(rstkram[542]) );
  DFFQ_X1M_A12TR rstkram_reg_4__14_ ( .D(n2377), .CK(wb_clk_o), .Q(
        rstkram[554]) );
  DFFQ_X1M_A12TR rstkram_reg_4__19_ ( .D(n2601), .CK(wb_clk_o), .Q(
        rstkram[559]) );
  DFFQ_X1M_A12TR rstkram_reg_0__3_ ( .D(n2221), .CK(wb_clk_o), .Q(rstkram[623]) );
  DFFQ_X1M_A12TR rstkram_reg_0__2_ ( .D(n2253), .CK(wb_clk_o), .Q(rstkram[622]) );
  DFFQ_X1M_A12TR rstkram_reg_0__14_ ( .D(n2381), .CK(wb_clk_o), .Q(
        rstkram[634]) );
  DFFQ_X1M_A12TR rstkram_reg_0__19_ ( .D(n2605), .CK(wb_clk_o), .Q(
        rstkram[639]) );
  DFFQ_X1M_A12TR rstkram_reg_28__7_ ( .D(n2065), .CK(wb_clk_o), .Q(rstkram[67]) );
  DFFQ_X1M_A12TR rstkram_reg_24__7_ ( .D(n2069), .CK(wb_clk_o), .Q(
        rstkram[147]) );
  DFFQ_X1M_A12TR rstkram_reg_20__7_ ( .D(n2073), .CK(wb_clk_o), .Q(
        rstkram[227]) );
  DFFQ_X1M_A12TR rstkram_reg_16__7_ ( .D(n2077), .CK(wb_clk_o), .Q(
        rstkram[307]) );
  DFFQ_X1M_A12TR rstkram_reg_12__7_ ( .D(n2081), .CK(wb_clk_o), .Q(
        rstkram[387]) );
  DFFQ_X1M_A12TR rstkram_reg_8__7_ ( .D(n2085), .CK(wb_clk_o), .Q(rstkram[467]) );
  DFFQ_X1M_A12TR rstkram_reg_4__7_ ( .D(n2089), .CK(wb_clk_o), .Q(rstkram[547]) );
  DFFQ_X1M_A12TR rstkram_reg_0__7_ ( .D(n2093), .CK(wb_clk_o), .Q(rstkram[627]) );
  DFFQ_X1M_A12TR rstkram_reg_28__5_ ( .D(n2129), .CK(wb_clk_o), .Q(rstkram[65]) );
  DFFQ_X1M_A12TR rstkram_reg_24__5_ ( .D(n2133), .CK(wb_clk_o), .Q(
        rstkram[145]) );
  DFFQ_X1M_A12TR rstkram_reg_20__5_ ( .D(n2137), .CK(wb_clk_o), .Q(
        rstkram[225]) );
  DFFQ_X1M_A12TR rstkram_reg_16__5_ ( .D(n2141), .CK(wb_clk_o), .Q(
        rstkram[305]) );
  DFFQ_X1M_A12TR rstkram_reg_12__5_ ( .D(n2145), .CK(wb_clk_o), .Q(
        rstkram[385]) );
  DFFQ_X1M_A12TR rstkram_reg_8__5_ ( .D(n2149), .CK(wb_clk_o), .Q(rstkram[465]) );
  DFFQ_X1M_A12TR rstkram_reg_4__5_ ( .D(n2153), .CK(wb_clk_o), .Q(rstkram[545]) );
  DFFQ_X1M_A12TR rstkram_reg_0__5_ ( .D(n2157), .CK(wb_clk_o), .Q(rstkram[625]) );
  DFFQ_X1M_A12TR rstkram_reg_28__1_ ( .D(n2257), .CK(wb_clk_o), .Q(rstkram[61]) );
  DFFQ_X1M_A12TR rstkram_reg_24__1_ ( .D(n2261), .CK(wb_clk_o), .Q(
        rstkram[141]) );
  DFFQ_X1M_A12TR rstkram_reg_20__1_ ( .D(n2265), .CK(wb_clk_o), .Q(
        rstkram[221]) );
  DFFQ_X1M_A12TR rstkram_reg_16__1_ ( .D(n2269), .CK(wb_clk_o), .Q(
        rstkram[301]) );
  DFFQ_X1M_A12TR rstkram_reg_12__1_ ( .D(n2273), .CK(wb_clk_o), .Q(
        rstkram[381]) );
  DFFQ_X1M_A12TR rstkram_reg_8__1_ ( .D(n2277), .CK(wb_clk_o), .Q(rstkram[461]) );
  DFFQ_X1M_A12TR rstkram_reg_4__1_ ( .D(n2281), .CK(wb_clk_o), .Q(rstkram[541]) );
  DFFQ_X1M_A12TR rstkram_reg_0__1_ ( .D(n2285), .CK(wb_clk_o), .Q(rstkram[621]) );
  DFFQ_X1M_A12TR rstkram_reg_28__4_ ( .D(n2161), .CK(wb_clk_o), .Q(rstkram[64]) );
  DFFQ_X1M_A12TR rstkram_reg_24__4_ ( .D(n2165), .CK(wb_clk_o), .Q(
        rstkram[144]) );
  DFFQ_X1M_A12TR rstkram_reg_20__4_ ( .D(n2169), .CK(wb_clk_o), .Q(
        rstkram[224]) );
  DFFQ_X1M_A12TR rstkram_reg_16__4_ ( .D(n2173), .CK(wb_clk_o), .Q(
        rstkram[304]) );
  DFFQ_X1M_A12TR rstkram_reg_12__4_ ( .D(n2177), .CK(wb_clk_o), .Q(
        rstkram[384]) );
  DFFQ_X1M_A12TR rstkram_reg_8__4_ ( .D(n2181), .CK(wb_clk_o), .Q(rstkram[464]) );
  DFFQ_X1M_A12TR rstkram_reg_4__4_ ( .D(n2185), .CK(wb_clk_o), .Q(rstkram[544]) );
  DFFQ_X1M_A12TR rstkram_reg_0__4_ ( .D(n2189), .CK(wb_clk_o), .Q(rstkram[624]) );
  DFFQ_X1M_A12TR rstkram_reg_28__13_ ( .D(n2385), .CK(wb_clk_o), .Q(
        rstkram[73]) );
  DFFQ_X1M_A12TR rstkram_reg_24__13_ ( .D(n2389), .CK(wb_clk_o), .Q(
        rstkram[153]) );
  DFFQ_X1M_A12TR rstkram_reg_20__13_ ( .D(n2393), .CK(wb_clk_o), .Q(
        rstkram[233]) );
  DFFQ_X1M_A12TR rstkram_reg_16__13_ ( .D(n2397), .CK(wb_clk_o), .Q(
        rstkram[313]) );
  DFFQ_X1M_A12TR rstkram_reg_12__13_ ( .D(n2401), .CK(wb_clk_o), .Q(
        rstkram[393]) );
  DFFQ_X1M_A12TR rstkram_reg_8__13_ ( .D(n2405), .CK(wb_clk_o), .Q(
        rstkram[473]) );
  DFFQ_X1M_A12TR rstkram_reg_4__13_ ( .D(n2409), .CK(wb_clk_o), .Q(
        rstkram[553]) );
  DFFQ_X1M_A12TR rstkram_reg_0__13_ ( .D(n2413), .CK(wb_clk_o), .Q(
        rstkram[633]) );
  DFFQ_X1M_A12TR rstkram_reg_28__12_ ( .D(n2417), .CK(wb_clk_o), .Q(
        rstkram[72]) );
  DFFQ_X1M_A12TR rstkram_reg_24__12_ ( .D(n2421), .CK(wb_clk_o), .Q(
        rstkram[152]) );
  DFFQ_X1M_A12TR rstkram_reg_20__12_ ( .D(n2425), .CK(wb_clk_o), .Q(
        rstkram[232]) );
  DFFQ_X1M_A12TR rstkram_reg_16__12_ ( .D(n2429), .CK(wb_clk_o), .Q(
        rstkram[312]) );
  DFFQ_X1M_A12TR rstkram_reg_12__12_ ( .D(n2433), .CK(wb_clk_o), .Q(
        rstkram[392]) );
  DFFQ_X1M_A12TR rstkram_reg_8__12_ ( .D(n2437), .CK(wb_clk_o), .Q(
        rstkram[472]) );
  DFFQ_X1M_A12TR rstkram_reg_4__12_ ( .D(n2441), .CK(wb_clk_o), .Q(
        rstkram[552]) );
  DFFQ_X1M_A12TR rstkram_reg_0__12_ ( .D(n2445), .CK(wb_clk_o), .Q(
        rstkram[632]) );
  DFFQ_X1M_A12TR rstkram_reg_28__11_ ( .D(n2449), .CK(wb_clk_o), .Q(
        rstkram[71]) );
  DFFQ_X1M_A12TR rstkram_reg_24__11_ ( .D(n2453), .CK(wb_clk_o), .Q(
        rstkram[151]) );
  DFFQ_X1M_A12TR rstkram_reg_20__11_ ( .D(n2457), .CK(wb_clk_o), .Q(
        rstkram[231]) );
  DFFQ_X1M_A12TR rstkram_reg_16__11_ ( .D(n2461), .CK(wb_clk_o), .Q(
        rstkram[311]) );
  DFFQ_X1M_A12TR rstkram_reg_12__11_ ( .D(n2465), .CK(wb_clk_o), .Q(
        rstkram[391]) );
  DFFQ_X1M_A12TR rstkram_reg_8__11_ ( .D(n2469), .CK(wb_clk_o), .Q(
        rstkram[471]) );
  DFFQ_X1M_A12TR rstkram_reg_4__11_ ( .D(n2473), .CK(wb_clk_o), .Q(
        rstkram[551]) );
  DFFQ_X1M_A12TR rstkram_reg_0__11_ ( .D(n2477), .CK(wb_clk_o), .Q(
        rstkram[631]) );
  DFFQ_X1M_A12TR rstkram_reg_28__10_ ( .D(n2481), .CK(wb_clk_o), .Q(
        rstkram[70]) );
  DFFQ_X1M_A12TR rstkram_reg_24__10_ ( .D(n2485), .CK(wb_clk_o), .Q(
        rstkram[150]) );
  DFFQ_X1M_A12TR rstkram_reg_20__10_ ( .D(n2489), .CK(wb_clk_o), .Q(
        rstkram[230]) );
  DFFQ_X1M_A12TR rstkram_reg_16__10_ ( .D(n2493), .CK(wb_clk_o), .Q(
        rstkram[310]) );
  DFFQ_X1M_A12TR rstkram_reg_12__10_ ( .D(n2497), .CK(wb_clk_o), .Q(
        rstkram[390]) );
  DFFQ_X1M_A12TR rstkram_reg_8__10_ ( .D(n2501), .CK(wb_clk_o), .Q(
        rstkram[470]) );
  DFFQ_X1M_A12TR rstkram_reg_4__10_ ( .D(n2505), .CK(wb_clk_o), .Q(
        rstkram[550]) );
  DFFQ_X1M_A12TR rstkram_reg_0__10_ ( .D(n2509), .CK(wb_clk_o), .Q(
        rstkram[630]) );
  DFFQ_X1M_A12TR rstkram_reg_28__9_ ( .D(n2513), .CK(wb_clk_o), .Q(rstkram[69]) );
  DFFQ_X1M_A12TR rstkram_reg_24__9_ ( .D(n2517), .CK(wb_clk_o), .Q(
        rstkram[149]) );
  DFFQ_X1M_A12TR rstkram_reg_20__9_ ( .D(n2521), .CK(wb_clk_o), .Q(
        rstkram[229]) );
  DFFQ_X1M_A12TR rstkram_reg_16__9_ ( .D(n2525), .CK(wb_clk_o), .Q(
        rstkram[309]) );
  DFFQ_X1M_A12TR rstkram_reg_12__9_ ( .D(n2529), .CK(wb_clk_o), .Q(
        rstkram[389]) );
  DFFQ_X1M_A12TR rstkram_reg_8__9_ ( .D(n2533), .CK(wb_clk_o), .Q(rstkram[469]) );
  DFFQ_X1M_A12TR rstkram_reg_4__9_ ( .D(n2537), .CK(wb_clk_o), .Q(rstkram[549]) );
  DFFQ_X1M_A12TR rstkram_reg_0__9_ ( .D(n2541), .CK(wb_clk_o), .Q(rstkram[629]) );
  DFFQ_X1M_A12TR rstkram_reg_28__8_ ( .D(n2545), .CK(wb_clk_o), .Q(rstkram[68]) );
  DFFQ_X1M_A12TR rstkram_reg_24__8_ ( .D(n2549), .CK(wb_clk_o), .Q(
        rstkram[148]) );
  DFFQ_X1M_A12TR rstkram_reg_20__8_ ( .D(n2553), .CK(wb_clk_o), .Q(
        rstkram[228]) );
  DFFQ_X1M_A12TR rstkram_reg_16__8_ ( .D(n2557), .CK(wb_clk_o), .Q(
        rstkram[308]) );
  DFFQ_X1M_A12TR rstkram_reg_12__8_ ( .D(n2561), .CK(wb_clk_o), .Q(
        rstkram[388]) );
  DFFQ_X1M_A12TR rstkram_reg_8__8_ ( .D(n2565), .CK(wb_clk_o), .Q(rstkram[468]) );
  DFFQ_X1M_A12TR rstkram_reg_4__8_ ( .D(n2569), .CK(wb_clk_o), .Q(rstkram[548]) );
  DFFQ_X1M_A12TR rstkram_reg_0__8_ ( .D(n2573), .CK(wb_clk_o), .Q(rstkram[628]) );
  DFFQ_X1M_A12TR rstkram_reg_28__6_ ( .D(n2097), .CK(wb_clk_o), .Q(rstkram[66]) );
  DFFQ_X1M_A12TR rstkram_reg_24__6_ ( .D(n2101), .CK(wb_clk_o), .Q(
        rstkram[146]) );
  DFFQ_X1M_A12TR rstkram_reg_20__6_ ( .D(n2105), .CK(wb_clk_o), .Q(
        rstkram[226]) );
  DFFQ_X1M_A12TR rstkram_reg_16__6_ ( .D(n2109), .CK(wb_clk_o), .Q(
        rstkram[306]) );
  DFFQ_X1M_A12TR rstkram_reg_12__6_ ( .D(n2113), .CK(wb_clk_o), .Q(
        rstkram[386]) );
  DFFQ_X1M_A12TR rstkram_reg_8__6_ ( .D(n2117), .CK(wb_clk_o), .Q(rstkram[466]) );
  DFFQ_X1M_A12TR rstkram_reg_4__6_ ( .D(n2121), .CK(wb_clk_o), .Q(rstkram[546]) );
  DFFQ_X1M_A12TR rstkram_reg_0__6_ ( .D(n2125), .CK(wb_clk_o), .Q(rstkram[626]) );
  DFFQ_X1M_A12TR rstkram_reg_28__15_ ( .D(n2321), .CK(wb_clk_o), .Q(
        rstkram[75]) );
  DFFQ_X1M_A12TR rstkram_reg_24__15_ ( .D(n2325), .CK(wb_clk_o), .Q(
        rstkram[155]) );
  DFFQ_X1M_A12TR rstkram_reg_20__15_ ( .D(n2329), .CK(wb_clk_o), .Q(
        rstkram[235]) );
  DFFQ_X1M_A12TR rstkram_reg_16__15_ ( .D(n2333), .CK(wb_clk_o), .Q(
        rstkram[315]) );
  DFFQ_X1M_A12TR rstkram_reg_12__15_ ( .D(n2337), .CK(wb_clk_o), .Q(
        rstkram[395]) );
  DFFQ_X1M_A12TR rstkram_reg_8__15_ ( .D(n2341), .CK(wb_clk_o), .Q(
        rstkram[475]) );
  DFFQ_X1M_A12TR rstkram_reg_4__15_ ( .D(n2345), .CK(wb_clk_o), .Q(
        rstkram[555]) );
  DFFQ_X1M_A12TR rstkram_reg_0__15_ ( .D(n2349), .CK(wb_clk_o), .Q(
        rstkram[635]) );
  DFFQ_X1M_A12TR rstkram_reg_28__16_ ( .D(n2673), .CK(wb_clk_o), .Q(
        rstkram[76]) );
  DFFQ_X1M_A12TR rstkram_reg_24__16_ ( .D(n2677), .CK(wb_clk_o), .Q(
        rstkram[156]) );
  DFFQ_X1M_A12TR rstkram_reg_20__16_ ( .D(n2681), .CK(wb_clk_o), .Q(
        rstkram[236]) );
  DFFQ_X1M_A12TR rstkram_reg_16__16_ ( .D(n2685), .CK(wb_clk_o), .Q(
        rstkram[316]) );
  DFFQ_X1M_A12TR rstkram_reg_12__16_ ( .D(n2689), .CK(wb_clk_o), .Q(
        rstkram[396]) );
  DFFQ_X1M_A12TR rstkram_reg_8__16_ ( .D(n2693), .CK(wb_clk_o), .Q(
        rstkram[476]) );
  DFFQ_X1M_A12TR rstkram_reg_4__16_ ( .D(n2697), .CK(wb_clk_o), .Q(
        rstkram[556]) );
  DFFQ_X1M_A12TR rstkram_reg_0__16_ ( .D(n2701), .CK(wb_clk_o), .Q(
        rstkram[636]) );
  DFFQ_X1M_A12TR rstkram_reg_28__17_ ( .D(n2641), .CK(wb_clk_o), .Q(
        rstkram[77]) );
  DFFQ_X1M_A12TR rstkram_reg_24__17_ ( .D(n2645), .CK(wb_clk_o), .Q(
        rstkram[157]) );
  DFFQ_X1M_A12TR rstkram_reg_20__17_ ( .D(n2649), .CK(wb_clk_o), .Q(
        rstkram[237]) );
  DFFQ_X1M_A12TR rstkram_reg_16__17_ ( .D(n2653), .CK(wb_clk_o), .Q(
        rstkram[317]) );
  DFFQ_X1M_A12TR rstkram_reg_12__17_ ( .D(n2657), .CK(wb_clk_o), .Q(
        rstkram[397]) );
  DFFQ_X1M_A12TR rstkram_reg_8__17_ ( .D(n2661), .CK(wb_clk_o), .Q(
        rstkram[477]) );
  DFFQ_X1M_A12TR rstkram_reg_4__17_ ( .D(n2665), .CK(wb_clk_o), .Q(
        rstkram[557]) );
  DFFQ_X1M_A12TR rstkram_reg_0__17_ ( .D(n2669), .CK(wb_clk_o), .Q(
        rstkram[637]) );
  DFFQ_X1M_A12TR rstkram_reg_28__18_ ( .D(n2609), .CK(wb_clk_o), .Q(
        rstkram[78]) );
  DFFQ_X1M_A12TR rstkram_reg_24__18_ ( .D(n2613), .CK(wb_clk_o), .Q(
        rstkram[158]) );
  DFFQ_X1M_A12TR rstkram_reg_20__18_ ( .D(n2617), .CK(wb_clk_o), .Q(
        rstkram[238]) );
  DFFQ_X1M_A12TR rstkram_reg_16__18_ ( .D(n2621), .CK(wb_clk_o), .Q(
        rstkram[318]) );
  DFFQ_X1M_A12TR rstkram_reg_12__18_ ( .D(n2625), .CK(wb_clk_o), .Q(
        rstkram[398]) );
  DFFQ_X1M_A12TR rstkram_reg_8__18_ ( .D(n2629), .CK(wb_clk_o), .Q(
        rstkram[478]) );
  DFFQ_X1M_A12TR rstkram_reg_4__18_ ( .D(n2633), .CK(wb_clk_o), .Q(
        rstkram[558]) );
  DFFQ_X1M_A12TR rstkram_reg_0__18_ ( .D(n2637), .CK(wb_clk_o), .Q(
        rstkram[638]) );
  DFFQ_X1M_A12TR rstkram_reg_28__0_ ( .D(n2289), .CK(wb_clk_o), .Q(rstkram[60]) );
  DFFQ_X1M_A12TR rstkram_reg_24__0_ ( .D(n2293), .CK(wb_clk_o), .Q(
        rstkram[140]) );
  DFFQ_X1M_A12TR rstkram_reg_20__0_ ( .D(n2297), .CK(wb_clk_o), .Q(
        rstkram[220]) );
  DFFQ_X1M_A12TR rstkram_reg_16__0_ ( .D(n2301), .CK(wb_clk_o), .Q(
        rstkram[300]) );
  DFFQ_X1M_A12TR rstkram_reg_12__0_ ( .D(n2305), .CK(wb_clk_o), .Q(
        rstkram[380]) );
  DFFQ_X1M_A12TR rstkram_reg_8__0_ ( .D(n2309), .CK(wb_clk_o), .Q(rstkram[460]) );
  DFFQ_X1M_A12TR rstkram_reg_4__0_ ( .D(n2313), .CK(wb_clk_o), .Q(rstkram[540]) );
  DFFQ_X1M_A12TR rstkram_reg_0__0_ ( .D(n2317), .CK(wb_clk_o), .Q(rstkram[620]) );
  DFFQ_X1M_A12TR rstkram_reg_30__3_ ( .D(n2191), .CK(wb_clk_o), .Q(rstkram[23]) );
  DFFQ_X1M_A12TR rstkram_reg_30__2_ ( .D(n2223), .CK(wb_clk_o), .Q(rstkram[22]) );
  DFFQ_X1M_A12TR rstkram_reg_30__14_ ( .D(n2351), .CK(wb_clk_o), .Q(
        rstkram[34]) );
  DFFQ_X1M_A12TR rstkram_reg_30__19_ ( .D(n2575), .CK(wb_clk_o), .Q(
        rstkram[39]) );
  DFFQ_X1M_A12TR rstkram_reg_26__3_ ( .D(n2195), .CK(wb_clk_o), .Q(
        rstkram[103]) );
  DFFQ_X1M_A12TR rstkram_reg_26__2_ ( .D(n2227), .CK(wb_clk_o), .Q(
        rstkram[102]) );
  DFFQ_X1M_A12TR rstkram_reg_26__14_ ( .D(n2355), .CK(wb_clk_o), .Q(
        rstkram[114]) );
  DFFQ_X1M_A12TR rstkram_reg_26__19_ ( .D(n2579), .CK(wb_clk_o), .Q(
        rstkram[119]) );
  DFFQ_X1M_A12TR rstkram_reg_22__3_ ( .D(n2199), .CK(wb_clk_o), .Q(
        rstkram[183]) );
  DFFQ_X1M_A12TR rstkram_reg_22__2_ ( .D(n2231), .CK(wb_clk_o), .Q(
        rstkram[182]) );
  DFFQ_X1M_A12TR rstkram_reg_22__14_ ( .D(n2359), .CK(wb_clk_o), .Q(
        rstkram[194]) );
  DFFQ_X1M_A12TR rstkram_reg_22__19_ ( .D(n2583), .CK(wb_clk_o), .Q(
        rstkram[199]) );
  DFFQ_X1M_A12TR rstkram_reg_18__3_ ( .D(n2203), .CK(wb_clk_o), .Q(
        rstkram[263]) );
  DFFQ_X1M_A12TR rstkram_reg_18__2_ ( .D(n2235), .CK(wb_clk_o), .Q(
        rstkram[262]) );
  DFFQ_X1M_A12TR rstkram_reg_18__14_ ( .D(n2363), .CK(wb_clk_o), .Q(
        rstkram[274]) );
  DFFQ_X1M_A12TR rstkram_reg_18__19_ ( .D(n2587), .CK(wb_clk_o), .Q(
        rstkram[279]) );
  DFFQ_X1M_A12TR rstkram_reg_14__3_ ( .D(n2207), .CK(wb_clk_o), .Q(
        rstkram[343]) );
  DFFQ_X1M_A12TR rstkram_reg_14__2_ ( .D(n2239), .CK(wb_clk_o), .Q(
        rstkram[342]) );
  DFFQ_X1M_A12TR rstkram_reg_14__14_ ( .D(n2367), .CK(wb_clk_o), .Q(
        rstkram[354]) );
  DFFQ_X1M_A12TR rstkram_reg_14__19_ ( .D(n2591), .CK(wb_clk_o), .Q(
        rstkram[359]) );
  DFFQ_X1M_A12TR rstkram_reg_10__3_ ( .D(n2211), .CK(wb_clk_o), .Q(
        rstkram[423]) );
  DFFQ_X1M_A12TR rstkram_reg_10__2_ ( .D(n2243), .CK(wb_clk_o), .Q(
        rstkram[422]) );
  DFFQ_X1M_A12TR rstkram_reg_10__14_ ( .D(n2371), .CK(wb_clk_o), .Q(
        rstkram[434]) );
  DFFQ_X1M_A12TR rstkram_reg_10__19_ ( .D(n2595), .CK(wb_clk_o), .Q(
        rstkram[439]) );
  DFFQ_X1M_A12TR rstkram_reg_6__3_ ( .D(n2215), .CK(wb_clk_o), .Q(rstkram[503]) );
  DFFQ_X1M_A12TR rstkram_reg_6__2_ ( .D(n2247), .CK(wb_clk_o), .Q(rstkram[502]) );
  DFFQ_X1M_A12TR rstkram_reg_6__14_ ( .D(n2375), .CK(wb_clk_o), .Q(
        rstkram[514]) );
  DFFQ_X1M_A12TR rstkram_reg_6__19_ ( .D(n2599), .CK(wb_clk_o), .Q(
        rstkram[519]) );
  DFFQ_X1M_A12TR rstkram_reg_2__3_ ( .D(n2219), .CK(wb_clk_o), .Q(rstkram[583]) );
  DFFQ_X1M_A12TR rstkram_reg_2__2_ ( .D(n2251), .CK(wb_clk_o), .Q(rstkram[582]) );
  DFFQ_X1M_A12TR rstkram_reg_2__14_ ( .D(n2379), .CK(wb_clk_o), .Q(
        rstkram[594]) );
  DFFQ_X1M_A12TR rstkram_reg_2__19_ ( .D(n2603), .CK(wb_clk_o), .Q(
        rstkram[599]) );
  DFFQ_X1M_A12TR rstkram_reg_30__7_ ( .D(n2063), .CK(wb_clk_o), .Q(rstkram[27]) );
  DFFQ_X1M_A12TR rstkram_reg_26__7_ ( .D(n2067), .CK(wb_clk_o), .Q(
        rstkram[107]) );
  DFFQ_X1M_A12TR rstkram_reg_22__7_ ( .D(n2071), .CK(wb_clk_o), .Q(
        rstkram[187]) );
  DFFQ_X1M_A12TR rstkram_reg_18__7_ ( .D(n2075), .CK(wb_clk_o), .Q(
        rstkram[267]) );
  DFFQ_X1M_A12TR rstkram_reg_14__7_ ( .D(n2079), .CK(wb_clk_o), .Q(
        rstkram[347]) );
  DFFQ_X1M_A12TR rstkram_reg_10__7_ ( .D(n2083), .CK(wb_clk_o), .Q(
        rstkram[427]) );
  DFFQ_X1M_A12TR rstkram_reg_6__7_ ( .D(n2087), .CK(wb_clk_o), .Q(rstkram[507]) );
  DFFQ_X1M_A12TR rstkram_reg_2__7_ ( .D(n2091), .CK(wb_clk_o), .Q(rstkram[587]) );
  DFFQ_X1M_A12TR rstkram_reg_30__5_ ( .D(n2127), .CK(wb_clk_o), .Q(rstkram[25]) );
  DFFQ_X1M_A12TR rstkram_reg_26__5_ ( .D(n2131), .CK(wb_clk_o), .Q(
        rstkram[105]) );
  DFFQ_X1M_A12TR rstkram_reg_22__5_ ( .D(n2135), .CK(wb_clk_o), .Q(
        rstkram[185]) );
  DFFQ_X1M_A12TR rstkram_reg_18__5_ ( .D(n2139), .CK(wb_clk_o), .Q(
        rstkram[265]) );
  DFFQ_X1M_A12TR rstkram_reg_14__5_ ( .D(n2143), .CK(wb_clk_o), .Q(
        rstkram[345]) );
  DFFQ_X1M_A12TR rstkram_reg_10__5_ ( .D(n2147), .CK(wb_clk_o), .Q(
        rstkram[425]) );
  DFFQ_X1M_A12TR rstkram_reg_6__5_ ( .D(n2151), .CK(wb_clk_o), .Q(rstkram[505]) );
  DFFQ_X1M_A12TR rstkram_reg_2__5_ ( .D(n2155), .CK(wb_clk_o), .Q(rstkram[585]) );
  DFFQ_X1M_A12TR rstkram_reg_30__1_ ( .D(n2255), .CK(wb_clk_o), .Q(rstkram[21]) );
  DFFQ_X1M_A12TR rstkram_reg_26__1_ ( .D(n2259), .CK(wb_clk_o), .Q(
        rstkram[101]) );
  DFFQ_X1M_A12TR rstkram_reg_22__1_ ( .D(n2263), .CK(wb_clk_o), .Q(
        rstkram[181]) );
  DFFQ_X1M_A12TR rstkram_reg_18__1_ ( .D(n2267), .CK(wb_clk_o), .Q(
        rstkram[261]) );
  DFFQ_X1M_A12TR rstkram_reg_14__1_ ( .D(n2271), .CK(wb_clk_o), .Q(
        rstkram[341]) );
  DFFQ_X1M_A12TR rstkram_reg_10__1_ ( .D(n2275), .CK(wb_clk_o), .Q(
        rstkram[421]) );
  DFFQ_X1M_A12TR rstkram_reg_6__1_ ( .D(n2279), .CK(wb_clk_o), .Q(rstkram[501]) );
  DFFQ_X1M_A12TR rstkram_reg_2__1_ ( .D(n2283), .CK(wb_clk_o), .Q(rstkram[581]) );
  DFFQ_X1M_A12TR rstkram_reg_30__4_ ( .D(n2159), .CK(wb_clk_o), .Q(rstkram[24]) );
  DFFQ_X1M_A12TR rstkram_reg_26__4_ ( .D(n2163), .CK(wb_clk_o), .Q(
        rstkram[104]) );
  DFFQ_X1M_A12TR rstkram_reg_22__4_ ( .D(n2167), .CK(wb_clk_o), .Q(
        rstkram[184]) );
  DFFQ_X1M_A12TR rstkram_reg_18__4_ ( .D(n2171), .CK(wb_clk_o), .Q(
        rstkram[264]) );
  DFFQ_X1M_A12TR rstkram_reg_14__4_ ( .D(n2175), .CK(wb_clk_o), .Q(
        rstkram[344]) );
  DFFQ_X1M_A12TR rstkram_reg_10__4_ ( .D(n2179), .CK(wb_clk_o), .Q(
        rstkram[424]) );
  DFFQ_X1M_A12TR rstkram_reg_6__4_ ( .D(n2183), .CK(wb_clk_o), .Q(rstkram[504]) );
  DFFQ_X1M_A12TR rstkram_reg_2__4_ ( .D(n2187), .CK(wb_clk_o), .Q(rstkram[584]) );
  DFFQ_X1M_A12TR rstkram_reg_30__13_ ( .D(n2383), .CK(wb_clk_o), .Q(
        rstkram[33]) );
  DFFQ_X1M_A12TR rstkram_reg_26__13_ ( .D(n2387), .CK(wb_clk_o), .Q(
        rstkram[113]) );
  DFFQ_X1M_A12TR rstkram_reg_22__13_ ( .D(n2391), .CK(wb_clk_o), .Q(
        rstkram[193]) );
  DFFQ_X1M_A12TR rstkram_reg_18__13_ ( .D(n2395), .CK(wb_clk_o), .Q(
        rstkram[273]) );
  DFFQ_X1M_A12TR rstkram_reg_14__13_ ( .D(n2399), .CK(wb_clk_o), .Q(
        rstkram[353]) );
  DFFQ_X1M_A12TR rstkram_reg_10__13_ ( .D(n2403), .CK(wb_clk_o), .Q(
        rstkram[433]) );
  DFFQ_X1M_A12TR rstkram_reg_6__13_ ( .D(n2407), .CK(wb_clk_o), .Q(
        rstkram[513]) );
  DFFQ_X1M_A12TR rstkram_reg_2__13_ ( .D(n2411), .CK(wb_clk_o), .Q(
        rstkram[593]) );
  DFFQ_X1M_A12TR rstkram_reg_30__12_ ( .D(n2415), .CK(wb_clk_o), .Q(
        rstkram[32]) );
  DFFQ_X1M_A12TR rstkram_reg_26__12_ ( .D(n2419), .CK(wb_clk_o), .Q(
        rstkram[112]) );
  DFFQ_X1M_A12TR rstkram_reg_22__12_ ( .D(n2423), .CK(wb_clk_o), .Q(
        rstkram[192]) );
  DFFQ_X1M_A12TR rstkram_reg_18__12_ ( .D(n2427), .CK(wb_clk_o), .Q(
        rstkram[272]) );
  DFFQ_X1M_A12TR rstkram_reg_14__12_ ( .D(n2431), .CK(wb_clk_o), .Q(
        rstkram[352]) );
  DFFQ_X1M_A12TR rstkram_reg_10__12_ ( .D(n2435), .CK(wb_clk_o), .Q(
        rstkram[432]) );
  DFFQ_X1M_A12TR rstkram_reg_6__12_ ( .D(n2439), .CK(wb_clk_o), .Q(
        rstkram[512]) );
  DFFQ_X1M_A12TR rstkram_reg_2__12_ ( .D(n2443), .CK(wb_clk_o), .Q(
        rstkram[592]) );
  DFFQ_X1M_A12TR rstkram_reg_30__11_ ( .D(n2447), .CK(wb_clk_o), .Q(
        rstkram[31]) );
  DFFQ_X1M_A12TR rstkram_reg_26__11_ ( .D(n2451), .CK(wb_clk_o), .Q(
        rstkram[111]) );
  DFFQ_X1M_A12TR rstkram_reg_22__11_ ( .D(n2455), .CK(wb_clk_o), .Q(
        rstkram[191]) );
  DFFQ_X1M_A12TR rstkram_reg_18__11_ ( .D(n2459), .CK(wb_clk_o), .Q(
        rstkram[271]) );
  DFFQ_X1M_A12TR rstkram_reg_14__11_ ( .D(n2463), .CK(wb_clk_o), .Q(
        rstkram[351]) );
  DFFQ_X1M_A12TR rstkram_reg_10__11_ ( .D(n2467), .CK(wb_clk_o), .Q(
        rstkram[431]) );
  DFFQ_X1M_A12TR rstkram_reg_6__11_ ( .D(n2471), .CK(wb_clk_o), .Q(
        rstkram[511]) );
  DFFQ_X1M_A12TR rstkram_reg_2__11_ ( .D(n2475), .CK(wb_clk_o), .Q(
        rstkram[591]) );
  DFFQ_X1M_A12TR rstkram_reg_30__10_ ( .D(n2479), .CK(wb_clk_o), .Q(
        rstkram[30]) );
  DFFQ_X1M_A12TR rstkram_reg_26__10_ ( .D(n2483), .CK(wb_clk_o), .Q(
        rstkram[110]) );
  DFFQ_X1M_A12TR rstkram_reg_22__10_ ( .D(n2487), .CK(wb_clk_o), .Q(
        rstkram[190]) );
  DFFQ_X1M_A12TR rstkram_reg_18__10_ ( .D(n2491), .CK(wb_clk_o), .Q(
        rstkram[270]) );
  DFFQ_X1M_A12TR rstkram_reg_14__10_ ( .D(n2495), .CK(wb_clk_o), .Q(
        rstkram[350]) );
  DFFQ_X1M_A12TR rstkram_reg_10__10_ ( .D(n2499), .CK(wb_clk_o), .Q(
        rstkram[430]) );
  DFFQ_X1M_A12TR rstkram_reg_6__10_ ( .D(n2503), .CK(wb_clk_o), .Q(
        rstkram[510]) );
  DFFQ_X1M_A12TR rstkram_reg_2__10_ ( .D(n2507), .CK(wb_clk_o), .Q(
        rstkram[590]) );
  DFFQ_X1M_A12TR rstkram_reg_30__9_ ( .D(n2511), .CK(wb_clk_o), .Q(rstkram[29]) );
  DFFQ_X1M_A12TR rstkram_reg_26__9_ ( .D(n2515), .CK(wb_clk_o), .Q(
        rstkram[109]) );
  DFFQ_X1M_A12TR rstkram_reg_22__9_ ( .D(n2519), .CK(wb_clk_o), .Q(
        rstkram[189]) );
  DFFQ_X1M_A12TR rstkram_reg_18__9_ ( .D(n2523), .CK(wb_clk_o), .Q(
        rstkram[269]) );
  DFFQ_X1M_A12TR rstkram_reg_14__9_ ( .D(n2527), .CK(wb_clk_o), .Q(
        rstkram[349]) );
  DFFQ_X1M_A12TR rstkram_reg_10__9_ ( .D(n2531), .CK(wb_clk_o), .Q(
        rstkram[429]) );
  DFFQ_X1M_A12TR rstkram_reg_6__9_ ( .D(n2535), .CK(wb_clk_o), .Q(rstkram[509]) );
  DFFQ_X1M_A12TR rstkram_reg_2__9_ ( .D(n2539), .CK(wb_clk_o), .Q(rstkram[589]) );
  DFFQ_X1M_A12TR rstkram_reg_30__8_ ( .D(n2543), .CK(wb_clk_o), .Q(rstkram[28]) );
  DFFQ_X1M_A12TR rstkram_reg_26__8_ ( .D(n2547), .CK(wb_clk_o), .Q(
        rstkram[108]) );
  DFFQ_X1M_A12TR rstkram_reg_22__8_ ( .D(n2551), .CK(wb_clk_o), .Q(
        rstkram[188]) );
  DFFQ_X1M_A12TR rstkram_reg_18__8_ ( .D(n2555), .CK(wb_clk_o), .Q(
        rstkram[268]) );
  DFFQ_X1M_A12TR rstkram_reg_14__8_ ( .D(n2559), .CK(wb_clk_o), .Q(
        rstkram[348]) );
  DFFQ_X1M_A12TR rstkram_reg_10__8_ ( .D(n2563), .CK(wb_clk_o), .Q(
        rstkram[428]) );
  DFFQ_X1M_A12TR rstkram_reg_6__8_ ( .D(n2567), .CK(wb_clk_o), .Q(rstkram[508]) );
  DFFQ_X1M_A12TR rstkram_reg_2__8_ ( .D(n2571), .CK(wb_clk_o), .Q(rstkram[588]) );
  DFFQ_X1M_A12TR rstkram_reg_30__6_ ( .D(n2095), .CK(wb_clk_o), .Q(rstkram[26]) );
  DFFQ_X1M_A12TR rstkram_reg_26__6_ ( .D(n2099), .CK(wb_clk_o), .Q(
        rstkram[106]) );
  DFFQ_X1M_A12TR rstkram_reg_22__6_ ( .D(n2103), .CK(wb_clk_o), .Q(
        rstkram[186]) );
  DFFQ_X1M_A12TR rstkram_reg_18__6_ ( .D(n2107), .CK(wb_clk_o), .Q(
        rstkram[266]) );
  DFFQ_X1M_A12TR rstkram_reg_14__6_ ( .D(n2111), .CK(wb_clk_o), .Q(
        rstkram[346]) );
  DFFQ_X1M_A12TR rstkram_reg_10__6_ ( .D(n2115), .CK(wb_clk_o), .Q(
        rstkram[426]) );
  DFFQ_X1M_A12TR rstkram_reg_6__6_ ( .D(n2119), .CK(wb_clk_o), .Q(rstkram[506]) );
  DFFQ_X1M_A12TR rstkram_reg_2__6_ ( .D(n2123), .CK(wb_clk_o), .Q(rstkram[586]) );
  DFFQ_X1M_A12TR rstkram_reg_30__15_ ( .D(n2319), .CK(wb_clk_o), .Q(
        rstkram[35]) );
  DFFQ_X1M_A12TR rstkram_reg_26__15_ ( .D(n2323), .CK(wb_clk_o), .Q(
        rstkram[115]) );
  DFFQ_X1M_A12TR rstkram_reg_22__15_ ( .D(n2327), .CK(wb_clk_o), .Q(
        rstkram[195]) );
  DFFQ_X1M_A12TR rstkram_reg_18__15_ ( .D(n2331), .CK(wb_clk_o), .Q(
        rstkram[275]) );
  DFFQ_X1M_A12TR rstkram_reg_14__15_ ( .D(n2335), .CK(wb_clk_o), .Q(
        rstkram[355]) );
  DFFQ_X1M_A12TR rstkram_reg_10__15_ ( .D(n2339), .CK(wb_clk_o), .Q(
        rstkram[435]) );
  DFFQ_X1M_A12TR rstkram_reg_6__15_ ( .D(n2343), .CK(wb_clk_o), .Q(
        rstkram[515]) );
  DFFQ_X1M_A12TR rstkram_reg_2__15_ ( .D(n2347), .CK(wb_clk_o), .Q(
        rstkram[595]) );
  DFFQ_X1M_A12TR rstkram_reg_30__16_ ( .D(n2671), .CK(wb_clk_o), .Q(
        rstkram[36]) );
  DFFQ_X1M_A12TR rstkram_reg_26__16_ ( .D(n2675), .CK(wb_clk_o), .Q(
        rstkram[116]) );
  DFFQ_X1M_A12TR rstkram_reg_22__16_ ( .D(n2679), .CK(wb_clk_o), .Q(
        rstkram[196]) );
  DFFQ_X1M_A12TR rstkram_reg_18__16_ ( .D(n2683), .CK(wb_clk_o), .Q(
        rstkram[276]) );
  DFFQ_X1M_A12TR rstkram_reg_14__16_ ( .D(n2687), .CK(wb_clk_o), .Q(
        rstkram[356]) );
  DFFQ_X1M_A12TR rstkram_reg_10__16_ ( .D(n2691), .CK(wb_clk_o), .Q(
        rstkram[436]) );
  DFFQ_X1M_A12TR rstkram_reg_6__16_ ( .D(n2695), .CK(wb_clk_o), .Q(
        rstkram[516]) );
  DFFQ_X1M_A12TR rstkram_reg_2__16_ ( .D(n2699), .CK(wb_clk_o), .Q(
        rstkram[596]) );
  DFFQ_X1M_A12TR rstkram_reg_30__17_ ( .D(n2639), .CK(wb_clk_o), .Q(
        rstkram[37]) );
  DFFQ_X1M_A12TR rstkram_reg_26__17_ ( .D(n2643), .CK(wb_clk_o), .Q(
        rstkram[117]) );
  DFFQ_X1M_A12TR rstkram_reg_22__17_ ( .D(n2647), .CK(wb_clk_o), .Q(
        rstkram[197]) );
  DFFQ_X1M_A12TR rstkram_reg_18__17_ ( .D(n2651), .CK(wb_clk_o), .Q(
        rstkram[277]) );
  DFFQ_X1M_A12TR rstkram_reg_14__17_ ( .D(n2655), .CK(wb_clk_o), .Q(
        rstkram[357]) );
  DFFQ_X1M_A12TR rstkram_reg_10__17_ ( .D(n2659), .CK(wb_clk_o), .Q(
        rstkram[437]) );
  DFFQ_X1M_A12TR rstkram_reg_6__17_ ( .D(n2663), .CK(wb_clk_o), .Q(
        rstkram[517]) );
  DFFQ_X1M_A12TR rstkram_reg_2__17_ ( .D(n2667), .CK(wb_clk_o), .Q(
        rstkram[597]) );
  DFFQ_X1M_A12TR rstkram_reg_30__18_ ( .D(n2607), .CK(wb_clk_o), .Q(
        rstkram[38]) );
  DFFQ_X1M_A12TR rstkram_reg_26__18_ ( .D(n2611), .CK(wb_clk_o), .Q(
        rstkram[118]) );
  DFFQ_X1M_A12TR rstkram_reg_22__18_ ( .D(n2615), .CK(wb_clk_o), .Q(
        rstkram[198]) );
  DFFQ_X1M_A12TR rstkram_reg_18__18_ ( .D(n2619), .CK(wb_clk_o), .Q(
        rstkram[278]) );
  DFFQ_X1M_A12TR rstkram_reg_14__18_ ( .D(n2623), .CK(wb_clk_o), .Q(
        rstkram[358]) );
  DFFQ_X1M_A12TR rstkram_reg_10__18_ ( .D(n2627), .CK(wb_clk_o), .Q(
        rstkram[438]) );
  DFFQ_X1M_A12TR rstkram_reg_6__18_ ( .D(n2631), .CK(wb_clk_o), .Q(
        rstkram[518]) );
  DFFQ_X1M_A12TR rstkram_reg_2__18_ ( .D(n2635), .CK(wb_clk_o), .Q(
        rstkram[598]) );
  DFFQ_X1M_A12TR rstkram_reg_30__0_ ( .D(n2287), .CK(wb_clk_o), .Q(rstkram[20]) );
  DFFQ_X1M_A12TR rstkram_reg_26__0_ ( .D(n2291), .CK(wb_clk_o), .Q(
        rstkram[100]) );
  DFFQ_X1M_A12TR rstkram_reg_22__0_ ( .D(n2295), .CK(wb_clk_o), .Q(
        rstkram[180]) );
  DFFQ_X1M_A12TR rstkram_reg_18__0_ ( .D(n2299), .CK(wb_clk_o), .Q(
        rstkram[260]) );
  DFFQ_X1M_A12TR rstkram_reg_14__0_ ( .D(n2303), .CK(wb_clk_o), .Q(
        rstkram[340]) );
  DFFQ_X1M_A12TR rstkram_reg_10__0_ ( .D(n2307), .CK(wb_clk_o), .Q(
        rstkram[420]) );
  DFFQ_X1M_A12TR rstkram_reg_6__0_ ( .D(n2311), .CK(wb_clk_o), .Q(rstkram[500]) );
  DFFQ_X1M_A12TR rstkram_reg_2__0_ ( .D(n2315), .CK(wb_clk_o), .Q(rstkram[580]) );
  DFFSQ_X1M_A12TR rswdten_reg ( .D(n1829), .CK(wb_clk_o), .SN(qrst), .Q(
        rswdten) );
  DFFNSRPQ_X1M_A12TR riwbwe_reg ( .D(n1660), .CKN(wb_clk_o), .R(n2807), .SN(n3), .Q(iwb_we_o) );
  DFFRPQ_X1M_A12TR rtosu_reg_4_ ( .D(n1649), .CK(wb_clk_o), .R(n2792), .Q(
        rtosu[4]) );
  DFFRPQ_X1M_A12TR rtosu_reg_6_ ( .D(n1648), .CK(wb_clk_o), .R(n2792), .Q(
        rtosu[6]) );
  DFFRPQ_X1M_A12TR rtosu_reg_7_ ( .D(n1647), .CK(wb_clk_o), .R(n2792), .Q(
        rtosu[7]) );
  DFFRPQ_X1M_A12TR rstatus__reg_0_ ( .D(n1646), .CK(wb_clk_o), .R(n2799), .Q(
        rstatus_[0]) );
  DFFRPQ_X1M_A12TR rtosu_reg_5_ ( .D(n1632), .CK(wb_clk_o), .R(n2792), .Q(
        rtosu[5]) );
  DFFRPQ_X1M_A12TR rwreg__reg_7_ ( .D(n1587), .CK(wb_clk_o), .R(n2798), .Q(
        rwreg_[7]) );
  DFFRPQ_X1M_A12TR rwreg__reg_6_ ( .D(n1583), .CK(wb_clk_o), .R(n2798), .Q(
        rwreg_[6]) );
  DFFRPQ_X1M_A12TR rwreg__reg_5_ ( .D(n1579), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg_[5]) );
  DFFRPQ_X1M_A12TR rwreg__reg_4_ ( .D(n1575), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg_[4]) );
  DFFRPQ_X1M_A12TR rwreg__reg_3_ ( .D(n1571), .CK(wb_clk_o), .R(n2791), .Q(
        rwreg_[3]) );
  DFFRPQ_X1M_A12TR rwreg__reg_2_ ( .D(n1567), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg_[2]) );
  DFFRPQ_X1M_A12TR rwreg__reg_1_ ( .D(n1563), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg_[1]) );
  DFFRPQ_X1M_A12TR rwreg__reg_0_ ( .D(n1559), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg_[0]) );
  DFFRPQ_X1M_A12TR rstatus__reg_2_ ( .D(n1556), .CK(wb_clk_o), .R(n2801), .Q(
        rstatus_[2]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_7_ ( .D(n1507), .CK(wb_clk_o), .R(n2792), .Q(
        rtblptru[7]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_6_ ( .D(n1506), .CK(wb_clk_o), .R(n2793), .Q(
        rtblptru[6]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_4_ ( .D(n1504), .CK(wb_clk_o), .R(n2793), .Q(
        rtblptru[4]) );
  DFFRPQ_X1M_A12TR rtablat_reg_5_ ( .D(n1467), .CK(wb_clk_o), .R(n2795), .Q(
        iwb_dat_o[13]) );
  DFFRPQ_X1M_A12TR rstatus__reg_4_ ( .D(n1414), .CK(wb_clk_o), .R(n2799), .Q(
        rstatus_[4]) );
  DFFNSRPQ_X1M_A12TR rinth_reg_2_ ( .D(rinth[1]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rinth[2]) );
  DFFNSRPQ_X1M_A12TR rintl_reg_2_ ( .D(rintl[1]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rintl[2]) );
  DFFNSRPQ_X1M_A12TR rqclk_reg_0_ ( .D(n1805), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(qena[0]) );
  DFFNSRPQ_X1M_A12TR rmxskp_reg_2_ ( .D(n1715), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rmxskp[2]) );
  DFFNSRPQ_X1M_A12TR rclrwdt__reg ( .D(n1676), .CKN(wb_clk_o), .R(n2807), .SN(
        n3), .Q(rclrwdt_) );
  DFFNSRPQ_X1M_A12TR rdwbwe_reg ( .D(n1662), .CKN(wb_clk_o), .R(n2807), .SN(n3), .Q(dwb_we_o) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_12_ ( .D(n2057), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[12]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_3_ ( .D(n1552), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(rpcnxt[3]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_7_ ( .D(n1982), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[7]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_6_ ( .D(n1983), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[6]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_5_ ( .D(n1984), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[5]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_4_ ( .D(n1985), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[4]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_3_ ( .D(n1986), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[3]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_2_ ( .D(n1987), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[2]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_1_ ( .D(n1988), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[1]) );
  DFFNSRPQ_X1M_A12TR rilat_reg_0_ ( .D(n1989), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rilat[0]) );
  DFFNSRPQ_X1M_A12TR rpcu_reg_4_ ( .D(n1461), .CKN(wb_clk_o), .R(n2818), .SN(
        n3), .Q(rpcu_4_) );
  DFFNSRPQ_X1M_A12TR riwbsel_reg_1_ ( .D(n1481), .CKN(wb_clk_o), .R(n2818), 
        .SN(n3), .Q(iwb_sel_o[1]) );
  DFFNSRPQ_X1M_A12TR riwbsel_reg_0_ ( .D(n1471), .CKN(wb_clk_o), .R(n2818), 
        .SN(n3), .Q(iwb_sel_o[0]) );
  DFFRPQ_X1M_A12TR rprodl_reg_0_ ( .D(n1952), .CK(wb_clk_o), .R(n2796), .Q(
        rprodl[0]) );
  DFFRPQ_X1M_A12TR rprodh_reg_1_ ( .D(n1959), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[1]) );
  DFFRPQ_X1M_A12TR rprodh_reg_2_ ( .D(n1958), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[2]) );
  DFFRPQ_X1M_A12TR rprodh_reg_3_ ( .D(n1957), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[3]) );
  DFFRPQ_X1M_A12TR rprodh_reg_4_ ( .D(n1956), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[4]) );
  DFFRPQ_X1M_A12TR rprodh_reg_0_ ( .D(n1960), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[0]) );
  DFFRPQ_X1M_A12TR rprodl_reg_1_ ( .D(n1951), .CK(wb_clk_o), .R(n2796), .Q(
        rprodl[1]) );
  DFFRPQ_X1M_A12TR rprodl_reg_2_ ( .D(n1950), .CK(wb_clk_o), .R(n2796), .Q(
        rprodl[2]) );
  DFFRPQ_X1M_A12TR rprodl_reg_3_ ( .D(n1949), .CK(wb_clk_o), .R(n2791), .Q(
        rprodl[3]) );
  DFFRPQ_X1M_A12TR rprodl_reg_4_ ( .D(n1948), .CK(wb_clk_o), .R(n2791), .Q(
        rprodl[4]) );
  DFFRPQ_X1M_A12TR rprodh_reg_6_ ( .D(n1954), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[6]) );
  DFFRPQ_X1M_A12TR rprodh_reg_7_ ( .D(n1953), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[7]) );
  DFFRPQ_X1M_A12TR rprodl_reg_6_ ( .D(n1945), .CK(wb_clk_o), .R(n2791), .Q(
        rprodl[6]) );
  DFFRPQ_X1M_A12TR rprodl_reg_7_ ( .D(n1944), .CK(wb_clk_o), .R(n2791), .Q(
        rprodl[7]) );
  DFFRPQ_X1M_A12TR rprodh_reg_5_ ( .D(n1955), .CK(wb_clk_o), .R(n2792), .Q(
        rprodh[5]) );
  DFFRPQ_X1M_A12TR rprodl_reg_5_ ( .D(n1947), .CK(wb_clk_o), .R(n2791), .Q(
        rprodl[5]) );
  DFFRPQ_X1M_A12TR rstatus__reg_1_ ( .D(n1413), .CK(wb_clk_o), .R(n2794), .Q(
        rstatus_[1]) );
  DFFRPQ_X1M_A12TR rstatus__reg_3_ ( .D(n1645), .CK(wb_clk_o), .R(n2794), .Q(
        rstatus_[3]) );
  DFFRPQ_X1M_A12TR rbsr__reg_7_ ( .D(n1628), .CK(wb_clk_o), .R(n2794), .Q(
        rbsr_[7]) );
  DFFRPQ_X1M_A12TR rbsr__reg_6_ ( .D(n1625), .CK(wb_clk_o), .R(n2797), .Q(
        rbsr_[6]) );
  DFFRPQ_X1M_A12TR rbsr__reg_5_ ( .D(n1622), .CK(wb_clk_o), .R(n2797), .Q(
        rbsr_[5]) );
  DFFRPQ_X1M_A12TR rbsr__reg_4_ ( .D(n1619), .CK(wb_clk_o), .R(n2797), .Q(
        rbsr_[4]) );
  DFFRPQ_X1M_A12TR rbsr__reg_3_ ( .D(n1616), .CK(wb_clk_o), .R(n2798), .Q(
        rbsr_[3]) );
  DFFRPQ_X1M_A12TR rbsr__reg_2_ ( .D(n1613), .CK(wb_clk_o), .R(n2798), .Q(
        rbsr_[2]) );
  DFFRPQ_X1M_A12TR rbsr__reg_1_ ( .D(n1610), .CK(wb_clk_o), .R(n2798), .Q(
        rbsr_[1]) );
  DFFRPQ_X1M_A12TR rbsr__reg_0_ ( .D(n1607), .CK(wb_clk_o), .R(n2798), .Q(
        rbsr_[0]) );
  DFFRPQ_X1M_A12TR rpclath_reg_5_ ( .D(n1547), .CK(wb_clk_o), .R(n2802), .Q(
        rpclath[5]) );
  DFFRPQ_X1M_A12TR rpclath_reg_0_ ( .D(n1517), .CK(wb_clk_o), .R(n2801), .Q(
        rpclath[0]) );
  DFFRPQ_X1M_A12TR rtablat_reg_7_ ( .D(n1469), .CK(wb_clk_o), .R(n2795), .Q(
        iwb_dat_o[15]) );
  DFFRPQ_X1M_A12TR rtablat_reg_6_ ( .D(n1468), .CK(wb_clk_o), .R(n2795), .Q(
        iwb_dat_o[14]) );
  DFFRPQ_X1M_A12TR rtablat_reg_4_ ( .D(n1466), .CK(wb_clk_o), .R(n2794), .Q(
        iwb_dat_o[12]) );
  DFFRPQ_X1M_A12TR rtablat_reg_3_ ( .D(n1465), .CK(wb_clk_o), .R(n2794), .Q(
        iwb_dat_o[11]) );
  DFFRPQ_X1M_A12TR rtablat_reg_2_ ( .D(n1464), .CK(wb_clk_o), .R(n2794), .Q(
        iwb_dat_o[10]) );
  DFFRPQ_X1M_A12TR rtablat_reg_1_ ( .D(n1463), .CK(wb_clk_o), .R(n2794), .Q(
        iwb_dat_o[9]) );
  DFFRPQ_X1M_A12TR rstkunf_reg ( .D(n1872), .CK(wb_clk_o), .R(n2791), .Q(
        rstkunf) );
  DFFRPQ_X1M_A12TR rpclatu_reg_7_ ( .D(n1511), .CK(wb_clk_o), .R(n2793), .Q(
        rpclatu[7]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_6_ ( .D(n1510), .CK(wb_clk_o), .R(n2793), .Q(
        rpclatu[6]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_3_ ( .D(n1508), .CK(wb_clk_o), .R(n2803), .Q(
        rpclatu[3]) );
  DFFRPQ_X1M_A12TR rtablat_reg_0_ ( .D(n1462), .CK(wb_clk_o), .R(n2794), .Q(
        iwb_dat_o[8]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_4_ ( .D(n1459), .CK(wb_clk_o), .R(n2793), .Q(
        rpclatu[4]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_1_ ( .D(n1421), .CK(wb_clk_o), .R(n2803), .Q(
        rpclatu[1]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_2_ ( .D(n1417), .CK(wb_clk_o), .R(n2803), .Q(
        rpclatu[2]) );
  DFFRPQ_X1M_A12TR rpclath_reg_6_ ( .D(n1548), .CK(wb_clk_o), .R(n2802), .Q(
        rpclath[6]) );
  DFFRPQ_X1M_A12TR rpclath_reg_4_ ( .D(n1541), .CK(wb_clk_o), .R(n2802), .Q(
        rpclath[4]) );
  DFFRPQ_X1M_A12TR rpclath_reg_3_ ( .D(n1535), .CK(wb_clk_o), .R(n2801), .Q(
        rpclath[3]) );
  DFFRPQ_X1M_A12TR rpclath_reg_2_ ( .D(n1529), .CK(wb_clk_o), .R(n2801), .Q(
        rpclath[2]) );
  DFFRPQ_X1M_A12TR rpclath_reg_1_ ( .D(n1523), .CK(wb_clk_o), .R(n2793), .Q(
        rpclath[1]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_5_ ( .D(n1509), .CK(wb_clk_o), .R(n2793), .Q(
        rpclatu[5]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_5_ ( .D(n1505), .CK(wb_clk_o), .R(n2793), .Q(
        rtblptru[5]) );
  DFFRPQ_X1M_A12TR rpclath_reg_7_ ( .D(n1435), .CK(wb_clk_o), .R(n2802), .Q(
        rpclath[7]) );
  DFFRPQ_X1M_A12TR rpclatu_reg_0_ ( .D(n1428), .CK(wb_clk_o), .R(n2802), .Q(
        rpclatu[0]) );
  DFFRPQ_X1M_A12TR rstkful_reg ( .D(n1870), .CK(wb_clk_o), .R(n2791), .Q(
        rstkful) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_7_ ( .D(n2744), .CK(wb_clk_o), .R(n2800), .Q(
        rsfrdat[7]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_1_ ( .D(n2705), .CK(wb_clk_o), .R(n2805), .Q(
        rsfrdat[1]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_4_ ( .D(n2740), .CK(wb_clk_o), .R(n2801), .Q(
        rsfrdat[4]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_2_ ( .D(n2704), .CK(wb_clk_o), .R(n2805), .Q(
        rsfrdat[2]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_3_ ( .D(n2703), .CK(wb_clk_o), .R(n2804), .Q(
        rsfrdat[3]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_6_ ( .D(n2702), .CK(wb_clk_o), .R(n2803), .Q(
        rsfrdat[6]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_5_ ( .D(n1946), .CK(wb_clk_o), .R(n2802), .Q(
        rsfrdat[5]) );
  DFFRPQ_X1M_A12TR rsfrdat_reg_0_ ( .D(n2706), .CK(wb_clk_o), .R(n2791), .Q(
        rsfrdat[0]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_0_ ( .D(n1550), .CKN(wb_clk_o), .R(n2817), .SN(
        n3), .Q(rpcl_0_) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_9_ ( .D(n1454), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(dwb_adr_o[9]) );
  DFFNSRPQ_X1M_A12TR rsleep__reg ( .D(n1691), .CKN(wb_clk_o), .R(n2807), .SN(
        n3), .Q(rsleep_) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_13_ ( .D(n1501), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(rdwbadr[13]) );
  DFFNSRPQ_X1M_A12TR rmxstal_reg_2_ ( .D(n1644), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxstal[2]) );
  DFFNSRPQ_X1M_A12TR rintl_reg_0_ ( .D(int_i[0]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rintl[0]) );
  DFFNSRPQ_X1M_A12TR rmxskp_reg_0_ ( .D(n1766), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rmxskp[0]) );
  DFFNSRPQ_X1M_A12TR rqclk_reg_2_ ( .D(n1801), .CKN(wb_clk_o), .R(n2821), .SN(
        n3), .Q(qena[2]) );
  DFFNSRPQ_X1M_A12TR rmxsta_reg_1_ ( .D(n1747), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxsta[1]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_7_ ( .D(n1458), .CKN(wb_clk_o), .R(n2818), 
        .SN(n3), .Q(dwb_adr_o[7]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_10_ ( .D(n1452), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(dwb_adr_o[10]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_12_ ( .D(n1499), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rdwbadr[12]) );
  DFFNSRPQ_X1M_A12TR rclrwdt_reg ( .D(n845), .CKN(wb_clk_o), .R(n2807), .SN(n3), .Q(rclrwdt) );
  DFFNSRPQ_X1M_A12TR rmxsta_reg_0_ ( .D(n1749), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxsta[0]) );
  DFFNSRPQ_X1M_A12TR rintl_reg_1_ ( .D(rintl[0]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rintl[1]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_6_ ( .D(n1448), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(dwb_adr_o[6]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_11_ ( .D(n1450), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(dwb_adr_o[11]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_8_ ( .D(n1456), .CKN(wb_clk_o), .R(n2818), 
        .SN(n3), .Q(dwb_adr_o[8]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_15_ ( .D(n1503), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(rdwbadr[15]) );
  DFFNSRPQ_X1M_A12TR rpcu_reg_3_ ( .D(n1856), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[18]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_6_ ( .D(n1838), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[13]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_5_ ( .D(n1546), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[12]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_4_ ( .D(n1540), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[11]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_3_ ( .D(n1534), .CKN(wb_clk_o), .R(n2814), .SN(
        n3), .Q(wpclat[10]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_2_ ( .D(n1528), .CKN(wb_clk_o), .R(n2814), .SN(
        n3), .Q(wpclat[9]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_1_ ( .D(n1522), .CKN(wb_clk_o), .R(n2812), .SN(
        n3), .Q(wpclat[8]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_0_ ( .D(n1516), .CKN(wb_clk_o), .R(n2814), .SN(
        n3), .Q(wpclat[7]) );
  DFFNSRPQ_X1M_A12TR rpch_reg_7_ ( .D(n1437), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[14]) );
  DFFNSRPQ_X1M_A12TR rpcu_reg_0_ ( .D(n1430), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[15]) );
  DFFNSRPQ_X1M_A12TR rpcu_reg_1_ ( .D(n1423), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[16]) );
  DFFNSRPQ_X1M_A12TR rpcu_reg_2_ ( .D(n1419), .CKN(wb_clk_o), .R(n2815), .SN(
        n3), .Q(wpclat[17]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_2_ ( .D(n1846), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(rpcnxt[2]) );
  DFFNSRPQ_X1M_A12TR rmxsta_reg_2_ ( .D(n1701), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxsta[2]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_6_ ( .D(rprng[5]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[6]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_1_ ( .D(rprng[0]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[1]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_2_ ( .D(rprng[1]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[2]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_13_ ( .D(n2056), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[13]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_0_ ( .D(n1889), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(rpcnxt[0]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_1_ ( .D(n1861), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(rpcnxt[1]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_18_ ( .D(n1858), .CKN(wb_clk_o), .R(n2815), 
        .SN(n3), .Q(rpcnxt[18]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_17_ ( .D(n1843), .CKN(wb_clk_o), .R(n2815), 
        .SN(n3), .Q(rpcnxt[17]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_13_ ( .D(n1840), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[13]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_6_ ( .D(n1594), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rpcnxt[6]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_12_ ( .D(n1543), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[12]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_11_ ( .D(n1537), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[11]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_10_ ( .D(n1531), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[10]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_9_ ( .D(n1525), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(rpcnxt[9]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_8_ ( .D(n1519), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rpcnxt[8]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_7_ ( .D(n1513), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rpcnxt[7]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_5_ ( .D(n1443), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(rpcnxt[5]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_14_ ( .D(n1440), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[14]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_15_ ( .D(n1433), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[15]) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_16_ ( .D(n1426), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(rpcnxt[16]) );
  DFFNSRPQ_X1M_A12TR rinth_reg_0_ ( .D(int_i[1]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rinth[0]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_14_ ( .D(n1904), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(rdwbadr[14]) );
  DFFNSRPQ_X1M_A12TR rc__reg ( .D(n1495), .CKN(wb_clk_o), .R(n2817), .SN(n3), 
        .Q(rc_) );
  DFFNSRPQ_X1M_A12TR rfsm_reg_0_ ( .D(rnxt[0]), .CKN(wb_clk_o), .R(n2807), 
        .SN(n3), .Q(rfsm[0]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_2_ ( .D(n1780), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rmask[2]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_6_ ( .D(n1778), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rmask[6]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_3_ ( .D(n1770), .CKN(wb_clk_o), .R(n2821), .SN(
        n3), .Q(rmask[3]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_1_ ( .D(n1768), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rmask[1]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_7_ ( .D(n1762), .CKN(wb_clk_o), .R(n2821), .SN(
        n3), .Q(rmask[7]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_0_ ( .D(n262), .CKN(wb_clk_o), .R(n4431), .SN(
        n3), .Q(rprng[0]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_15_ ( .D(n2054), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(reaptr[15]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_4_ ( .D(n2018), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr1h[4]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_14_ ( .D(n2055), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[14]) );
  DFFNSRPQ_X1M_A12TR rfsm_reg_1_ ( .D(rnxt[1]), .CKN(wb_clk_o), .R(n2807), 
        .SN(n3), .Q(rfsm[1]) );
  DFFRPQ_X1M_A12TR rstkptr__reg_4_ ( .D(n1652), .CK(wb_clk_o), .R(n2803), .Q(
        rstkptr_[4]) );
  DFFRPQ_X1M_A12TR rbsr_reg_5_ ( .D(n1623), .CK(wb_clk_o), .R(n2797), .Q(
        wfilebsr[13]) );
  DFFRPQ_X1M_A12TR rdc_reg ( .D(n2707), .CK(wb_clk_o), .R(n2794), .Q(rdc) );
  DFFNSRPQ_X1M_A12TR rmxtbl_reg_2_ ( .D(n1717), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rmxtbl[2]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_5_ ( .D(n1638), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(wpclat[4]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_7_ ( .D(n2015), .CK(wb_clk_o), .R(n2793), .Q(
        rfsr1h[7]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_6_ ( .D(n2016), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr1h[6]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_5_ ( .D(n2017), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr1h[5]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_4_ ( .D(n2034), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr0h[4]) );
  DFFRPQ_X1M_A12TR rbsr_reg_0_ ( .D(n1608), .CK(wb_clk_o), .R(n2798), .Q(
        wfilebsr[8]) );
  DFFRPQ_X1M_A12TR rstkptr__reg_3_ ( .D(n1653), .CK(wb_clk_o), .R(n2804), .Q(
        rstkptr_[3]) );
  DFFNSRPQ_X1M_A12TR rinth_reg_1_ ( .D(rinth[0]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rinth[1]) );
  DFFNSRPQ_X1M_A12TR rmxnpc_reg_0_ ( .D(n1713), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rmxnpc[0]) );
  DFFNSRPQ_X1M_A12TR rmxsha_reg_0_ ( .D(n1682), .CKN(wb_clk_o), .R(n2807), 
        .SN(n3), .Q(rmxsha[0]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_7_ ( .D(n2031), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr0h[7]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_6_ ( .D(n2032), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr0h[6]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_5_ ( .D(n2033), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr0h[5]) );
  DFFRPQ_X1M_A12TR rbsr_reg_7_ ( .D(n1629), .CK(wb_clk_o), .R(n2793), .Q(
        wfilebsr[15]) );
  DFFRPQ_X1M_A12TR rbsr_reg_6_ ( .D(n1626), .CK(wb_clk_o), .R(n2797), .Q(
        wfilebsr[14]) );
  DFFRPQ_X1M_A12TR rbsr_reg_4_ ( .D(n1620), .CK(wb_clk_o), .R(n2798), .Q(
        wfilebsr[12]) );
  DFFRPQ_X1M_A12TR rbsr_reg_3_ ( .D(n1617), .CK(wb_clk_o), .R(n2798), .Q(
        wfilebsr[11]) );
  DFFRPQ_X1M_A12TR rbsr_reg_2_ ( .D(n1614), .CK(wb_clk_o), .R(n2798), .Q(
        wfilebsr[10]) );
  DFFRPQ_X1M_A12TR rbsr_reg_1_ ( .D(n1611), .CK(wb_clk_o), .R(n2798), .Q(
        wfilebsr[9]) );
  DFFRPQ_X1M_A12TR rfsr2h_reg_4_ ( .D(n2010), .CK(wb_clk_o), .R(n2800), .Q(
        rfsr2h[4]) );
  DFFRPQ_X1M_A12TR rz_reg ( .D(n2741), .CK(wb_clk_o), .R(n2801), .Q(rz) );
  DFFRPQ_X1M_A12TR rn_reg ( .D(n2742), .CK(wb_clk_o), .R(n2800), .Q(rn) );
  DFFNSRPQ_X1M_A12TR rmxbcc_reg_1_ ( .D(n17841), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(rmxbcc[1]) );
  DFFNSRPQ_X1M_A12TR rmxskp_reg_1_ ( .D(n1774), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(rmxskp[1]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_7_ ( .D(rprng[6]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[7]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_6_ ( .D(n1733), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[6]) );
  DFFNSRPQ_X1M_A12TR rmxstk_reg_0_ ( .D(n1680), .CKN(wb_clk_o), .R(n2814), 
        .SN(n3), .Q(rmxstk[0]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_7_ ( .D(n1736), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[7]) );
  DFFNSRPQ_X1M_A12TR rdwbstb_reg ( .D(n1809), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(dwb_stb_o) );
  DFFNSRPQ_X1M_A12TR rmxtbl_reg_1_ ( .D(n1708), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rmxtbl[1]) );
  DFFNSRPQ_X1M_A12TR riwbstb_reg ( .D(n1658), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(iwb_stb_o) );
  DFFRPQ_X1M_A12TR rov_reg ( .D(n2743), .CK(wb_clk_o), .R(n2794), .Q(rov) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_11_ ( .D(n2058), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[11]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_10_ ( .D(n2059), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[10]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_8_ ( .D(n2061), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[8]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_9_ ( .D(n2060), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(reaptr[9]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_16_ ( .D(n2737), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(rwdt[16]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_4_ ( .D(n17821), .CKN(wb_clk_o), .R(n2820), 
        .SN(n3), .Q(rmask[4]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_0_ ( .D(n1776), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rmask[0]) );
  DFFNSRPQ_X1M_A12TR rmask_reg_5_ ( .D(n1772), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rmask[5]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_3_ ( .D(rprng[2]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[3]) );
  DFFNSRPQ_X1M_A12TR rmxstk_reg_1_ ( .D(n1678), .CKN(wb_clk_o), .R(n2807), 
        .SN(n3), .Q(rmxstk[1]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_4_ ( .D(n1727), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[4]) );
  DFFNSRPQ_X1M_A12TR rnskp_reg ( .D(n1906), .CKN(wb_clk_o), .R(iwb_adr_o[0]), 
        .SN(qrst), .Q(rnskp) );
  DFFNSRPQ_X1M_A12TR rpcnxt_reg_4_ ( .D(n1591), .CKN(wb_clk_o), .R(n2813), 
        .SN(n3), .Q(rpcnxt[4]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_0_ ( .D(n1705), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[0]) );
  DFFNSRPQ_X1M_A12TR rintf_reg_1_ ( .D(n2720), .CKN(wb_clk_o), .R(n4431), .SN(
        n3), .Q(rintf[1]) );
  DFFNSRPQ_X1M_A12TR rbcc_reg ( .D(n1891), .CKN(wb_clk_o), .R(n2812), .SN(n3), 
        .Q(rbcc) );
  DFFNSRPQ_X1M_A12TR rmxtbl_reg_0_ ( .D(n1703), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxtbl[0]) );
  DFFNSRPQ_X1M_A12TR rmxsha_reg_1_ ( .D(n1684), .CKN(wb_clk_o), .R(n2807), 
        .SN(n3), .Q(rmxsha[1]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_7_ ( .D(n1895), .CKN(wb_clk_o), .R(n2814), .SN(
        n3), .Q(wpclat[6]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_1_ ( .D(n1887), .CKN(wb_clk_o), .R(n2817), .SN(
        n3), .Q(wpclat[0]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_2_ ( .D(n1864), .CKN(wb_clk_o), .R(n2817), .SN(
        n3), .Q(wpclat[1]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_3_ ( .D(n1849), .CKN(wb_clk_o), .R(n2814), .SN(
        n3), .Q(wpclat[2]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_4_ ( .D(n1555), .CKN(wb_clk_o), .R(n2819), .SN(
        n3), .Q(wpclat[3]) );
  DFFNSRPQ_X1M_A12TR rpcl_reg_6_ ( .D(n1446), .CKN(wb_clk_o), .R(n2809), .SN(
        n3), .Q(wpclat[5]) );
  DFFNSRPQ_X1M_A12TR rmxtbl_reg_3_ ( .D(n1722), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rmxtbl[3]) );
  DFFNSRPQ_X1M_A12TR rmxbcc_reg_2_ ( .D(n17871), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rmxbcc[2]) );
  DFFNSRPQ_X1M_A12TR rmxdst_reg_1_ ( .D(n4434), .CKN(wb_clk_o), .R(n2806), 
        .SN(n3), .Q(rmxdst[1]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_5_ ( .D(rprng[4]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[5]) );
  DFFNSRPQ_X1M_A12TR rmxfsr_reg_1_ ( .D(n1605), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxfsr[1]) );
  DFFRPQ_X1M_A12TR rstkptr__reg_2_ ( .D(n1654), .CK(wb_clk_o), .R(n2803), .Q(
        rstkptr_[2]) );
  DFFRPQ_X1M_A12TR rstkptr__reg_1_ ( .D(n1655), .CK(wb_clk_o), .R(n2804), .Q(
        rstkptr_[1]) );
  DFFRPQ_X1M_A12TR rstkptr__reg_0_ ( .D(n1656), .CK(wb_clk_o), .R(n2795), .Q(
        rstkptr_[0]) );
  DFFNSRPQ_X1M_A12TR rprng_reg_4_ ( .D(rprng[3]), .CKN(wb_clk_o), .R(n4431), 
        .SN(n3), .Q(rprng[4]) );
  DFFNSRPQ_X1M_A12TR rmxfsr_reg_3_ ( .D(n1603), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(rmxfsr[3]) );
  DFFNSRPQ_X1M_A12TR rmxsrc_reg_0_ ( .D(n1755), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxsrc[0]) );
  DFFNSRPQ_X1M_A12TR rintf_reg_0_ ( .D(n2719), .CKN(wb_clk_o), .R(n4431), .SN(
        n3), .Q(rintf[0]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_5_ ( .D(n1730), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[5]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_4_ ( .D(n1875), .CKN(wb_clk_o), .R(n2813), 
        .SN(n3), .Q(dwb_adr_o[4]) );
  DFFNSRPQ_X1M_A12TR rmxsrc_reg_1_ ( .D(n1757), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxsrc[1]) );
  DFFNSRPQ_X1M_A12TR rsleep_reg ( .D(n846), .CKN(wb_clk_o), .R(n2807), .SN(n3), 
        .Q(rsleep) );
  DFFNSRPQ_X1M_A12TR rmxtgt_reg_1_ ( .D(n1743), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rmxtgt[1]) );
  DFFNSRPQ_X1M_A12TR rmxbsr_reg_0_ ( .D(n1751), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(rmxbsr[0]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_3_ ( .D(n1971), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[19]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_2_ ( .D(n1719), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[2]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_2_ ( .D(n2734), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[2]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_6_ ( .D(n2730), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[6]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_1_ ( .D(n1881), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(dwb_adr_o[1]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_0_ ( .D(n1597), .CKN(wb_clk_o), .R(n2813), 
        .SN(n3), .Q(dwb_adr_o[0]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_5_ ( .D(n2731), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[5]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_1_ ( .D(n2735), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[1]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_15_ ( .D(n2006), .CKN(wb_clk_o), .R(n2823), .SN(
        n3), .Q(rwdt[15]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_1_ ( .D(n1992), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[1]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_2_ ( .D(n1993), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[2]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_3_ ( .D(n1994), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[3]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_4_ ( .D(n1995), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[4]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_5_ ( .D(n1996), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[5]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_6_ ( .D(n1997), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[6]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_7_ ( .D(n1998), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[7]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_8_ ( .D(n1999), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[8]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_9_ ( .D(n2000), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[9]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_10_ ( .D(n2001), .CKN(wb_clk_o), .R(n2806), .SN(
        n3), .Q(rwdt[10]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_11_ ( .D(n2002), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(rwdt[11]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_12_ ( .D(n2003), .CKN(wb_clk_o), .R(n2823), .SN(
        n3), .Q(rwdt[12]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_13_ ( .D(n2004), .CKN(wb_clk_o), .R(n2823), .SN(
        n3), .Q(rwdt[13]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_14_ ( .D(n2005), .CKN(wb_clk_o), .R(n2823), .SN(
        n3), .Q(rwdt[14]) );
  DFFRPQ_X1M_A12TR rstkptr_reg_5_ ( .D(n1873), .CK(wb_clk_o), .R(n2791), .Q(
        rstkptr_5_) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_1_ ( .D(n1710), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[1]) );
  DFFNSRPQ_X1M_A12TR rmxtgt_reg_0_ ( .D(n1741), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(rmxtgt[0]) );
  DFFNSRPQ_X1M_A12TR rmxfsr_reg_2_ ( .D(n1601), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(rmxfsr[2]) );
  DFFNSRPQ_X1M_A12TR rmxstal_reg_1_ ( .D(n1640), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxstal[1]) );
  DFFNSRPQ_X1M_A12TR rmxnpc_reg_2_ ( .D(n17901), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rmxnpc[2]) );
  DFFNSRPQ_X1M_A12TR rmxdst_reg_0_ ( .D(n1699), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxdst[0]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_3_ ( .D(n2733), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[3]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_5_ ( .D(n1831), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(dwb_adr_o[5]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_4_ ( .D(n2732), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[4]) );
  DFFNSRPQ_X1M_A12TR reaptr_reg_3_ ( .D(n1724), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(reaptr[3]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_7_ ( .D(n2729), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[7]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_0_ ( .D(n2736), .CKN(wb_clk_o), .R(n2808), 
        .SN(n3), .Q(rromlat[0]) );
  DFFNSRPQ_X1M_A12TR rmxstal_reg_0_ ( .D(n1642), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxstal[0]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_9_ ( .D(n2709), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[9]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_8_ ( .D(n2710), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[8]) );
  DFFNSRPQ_X1M_A12TR rmxfsr_reg_0_ ( .D(n1599), .CKN(wb_clk_o), .R(n2819), 
        .SN(n3), .Q(rmxfsr[0]) );
  DFFNSRPQ_X1M_A12TR rmxalu_reg_3_ ( .D(n1697), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxalu[3]) );
  DFFNSRPQ_X1M_A12TR rmxbsr_reg_1_ ( .D(n1764), .CKN(wb_clk_o), .R(n2821), 
        .SN(n3), .Q(rmxbsr[1]) );
  DFFNSRPQ_X1M_A12TR rmxnpc_reg_1_ ( .D(n1753), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxnpc[1]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_15_ ( .D(n2721), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rromlat[15]) );
  DFFNSRPQ_X1M_A12TR rqcnt_reg_1_ ( .D(n17971), .CKN(wb_clk_o), .R(
        iwb_adr_o[0]), .SN(qrst), .Q(qfsm[1]) );
  DFFNSRPQ_X1M_A12TR rmxalu_reg_2_ ( .D(n1695), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxalu[2]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_12_ ( .D(n2724), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rromlat[12]) );
  DFFNSRPQ_X1M_A12TR rmxalu_reg_1_ ( .D(n1739), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxalu[1]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_3_ ( .D(n2019), .CK(wb_clk_o), .R(n2804), .Q(
        rfsr1h[3]) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_2_ ( .D(n1558), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(dwb_adr_o[2]) );
  DFFRPQ_X1M_A12TR rfsr2h_reg_3_ ( .D(n2011), .CK(wb_clk_o), .R(n2801), .Q(
        rfsr2h[3]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_3_ ( .D(n2035), .CK(wb_clk_o), .R(n2801), .Q(
        rfsr0h[3]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_0_ ( .D(n1970), .CK(wb_clk_o), .R(n2804), .Q(
        wtblat[8]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_1_ ( .D(n1973), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[17]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_2_ ( .D(n1972), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[18]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_8_ ( .D(n2728), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(rromlat[8]) );
  DFFNSRPQ_X1M_A12TR rmxbcc_reg_0_ ( .D(n1759), .CKN(wb_clk_o), .R(n2809), 
        .SN(n3), .Q(rmxbcc[0]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_11_ ( .D(n2725), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rromlat[11]) );
  DFFNSRPQ_X1M_A12TR rwdt_reg_0_ ( .D(n1991), .CKN(wb_clk_o), .R(n2807), .SN(
        n3), .Q(rwdt[0]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_10_ ( .D(n2726), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rromlat[10]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_13_ ( .D(n2723), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rromlat[13]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_2_ ( .D(n1866), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(dwb_dat_o[2]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_6_ ( .D(n1833), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(dwb_dat_o[6]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_5_ ( .D(n1634), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(dwb_dat_o[5]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_5_ ( .D(n1965), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[13]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_6_ ( .D(n1964), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[14]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_7_ ( .D(n1963), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[15]) );
  DFFRPQ_X1M_A12TR rtblptru_reg_0_ ( .D(n1974), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[16]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_5_ ( .D(n1977), .CK(wb_clk_o), .R(n2803), .Q(
        wtblat[5]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_6_ ( .D(n1976), .CK(wb_clk_o), .R(n2806), .Q(
        wtblat[6]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_7_ ( .D(n1975), .CK(wb_clk_o), .R(n2804), .Q(
        wtblat[7]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_1_ ( .D(n1969), .CK(wb_clk_o), .R(n2804), .Q(
        wtblat[9]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_2_ ( .D(n1968), .CK(wb_clk_o), .R(n2804), .Q(
        wtblat[10]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_3_ ( .D(n1967), .CK(wb_clk_o), .R(n2804), .Q(
        wtblat[11]) );
  DFFRPQ_X1M_A12TR rtblptrh_reg_4_ ( .D(n1966), .CK(wb_clk_o), .R(n2805), .Q(
        wtblat[12]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_1_ ( .D(n1981), .CK(wb_clk_o), .R(n2795), .Q(
        wtblat[1]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_2_ ( .D(n1980), .CK(wb_clk_o), .R(n2795), .Q(
        wtblat[2]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_3_ ( .D(n1979), .CK(wb_clk_o), .R(n2804), .Q(
        wtblat[3]) );
  DFFRPQ_X1M_A12TR rsfrstb_reg ( .D(n1902), .CK(wb_clk_o), .R(n2800), .Q(
        rsfrstb) );
  DFFNSRPQ_X1M_A12TR rdwbadr_reg_3_ ( .D(n1631), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(dwb_adr_o[3]) );
  DFFNSRPQ_X1M_A12TR rmxalu_reg_0_ ( .D(n1693), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rmxalu[0]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_0_ ( .D(n1899), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(dwb_dat_o[0]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_14_ ( .D(n2722), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(rromlat[14]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_1_ ( .D(n1883), .CKN(wb_clk_o), .R(n2813), 
        .SN(n3), .Q(dwb_dat_o[1]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_3_ ( .D(n1851), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(dwb_dat_o[3]) );
  DFFNSRPQ_X1M_A12TR rresult_reg_4_ ( .D(n1877), .CKN(wb_clk_o), .R(n2813), 
        .SN(n3), .Q(dwb_dat_o[4]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_4_ ( .D(n1978), .CK(wb_clk_o), .R(n2801), .Q(
        wtblat[4]) );
  DFFRPQN_X1M_A12TR rfsr2h_reg_7_ ( .D(n2007), .CK(wb_clk_o), .R(wb_rst_o), 
        .QN(n1940) );
  DFFRPQN_X1M_A12TR rfsr2h_reg_6_ ( .D(n2008), .CK(wb_clk_o), .R(n2823), .QN(
        n1941) );
  DFFRPQN_X1M_A12TR rfsr2h_reg_5_ ( .D(n2009), .CK(wb_clk_o), .R(wb_rst_o), 
        .QN(n1942) );
  DFFNSRPQ_X1M_A12TR rresult_reg_7_ ( .D(n1897), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(dwb_dat_o[7]) );
  DFFNSRPQ_X1M_A12TR rromlat_reg_9_ ( .D(n2727), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(rromlat[9]) );
  DFFRPQ_X1M_A12TR rwreg_reg_5_ ( .D(n1580), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg[5]) );
  DFFRPQ_X1M_A12TR rwreg_reg_7_ ( .D(n1588), .CK(wb_clk_o), .R(n2798), .Q(
        rwreg[7]) );
  DFFRPQ_X1M_A12TR rwreg_reg_6_ ( .D(n1584), .CK(wb_clk_o), .R(n2798), .Q(
        rwreg[6]) );
  DFFRPQ_X1M_A12TR rwreg_reg_4_ ( .D(n1576), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg[4]) );
  DFFRPQ_X1M_A12TR rwreg_reg_3_ ( .D(n1572), .CK(wb_clk_o), .R(n2791), .Q(
        rwreg[3]) );
  DFFRPQ_X1M_A12TR rwreg_reg_2_ ( .D(n1568), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg[2]) );
  DFFRPQ_X1M_A12TR rwreg_reg_1_ ( .D(n1564), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg[1]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_18_ ( .D(n1937), .CKN(wb_clk_o), .R(n2815), 
        .SN(n3), .Q(iwb_adr_o[19]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_6_ ( .D(n2712), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[6]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_5_ ( .D(n2713), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[5]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_5_ ( .D(n2025), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr1l[5]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_6_ ( .D(n2024), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr1l[6]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_7_ ( .D(n2023), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr1l[7]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_1_ ( .D(n2029), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr1l[1]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_2_ ( .D(n2028), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr1l[2]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_3_ ( .D(n2027), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr1l[3]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_4_ ( .D(n2026), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr1l[4]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_1_ ( .D(n2045), .CK(wb_clk_o), .R(n2795), .Q(
        rfsr0l[1]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_2_ ( .D(n2044), .CK(wb_clk_o), .R(n2795), .Q(
        rfsr0l[2]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_3_ ( .D(n2043), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr0l[3]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_4_ ( .D(n2042), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr0l[4]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_6_ ( .D(n2047), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr2l[6]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_7_ ( .D(n2738), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr2l[7]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_5_ ( .D(n2048), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr2l[5]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_1_ ( .D(n2052), .CK(wb_clk_o), .R(n2794), .Q(
        rfsr2l[1]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_4_ ( .D(n2049), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr2l[4]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_5_ ( .D(n2041), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr0l[5]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_3_ ( .D(n2050), .CK(wb_clk_o), .R(n2797), .Q(
        rfsr2l[3]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_2_ ( .D(n2051), .CK(wb_clk_o), .R(n2795), .Q(
        rfsr2l[2]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_6_ ( .D(n2040), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr0l[6]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_7_ ( .D(n2039), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr0l[7]) );
  DFFNSRPQ_X1M_A12TR rqcnt_reg_0_ ( .D(n1799), .CKN(wb_clk_o), .R(iwb_adr_o[0]), .SN(qrst), .Q(qfsm[0]) );
  DFFRPQ_X1M_A12TR rc_reg ( .D(n2739), .CK(wb_clk_o), .R(n2801), .Q(wrrc_7_)
         );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_1_ ( .D(n1922), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(iwb_adr_o[2]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_17_ ( .D(n1936), .CKN(wb_clk_o), .R(n2815), 
        .SN(n3), .Q(iwb_adr_o[18]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_4_ ( .D(n1923), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(iwb_adr_o[5]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_6_ ( .D(n1925), .CKN(wb_clk_o), .R(n2811), 
        .SN(n3), .Q(iwb_adr_o[7]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_7_ ( .D(n1926), .CKN(wb_clk_o), .R(n2812), 
        .SN(n3), .Q(iwb_adr_o[8]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_8_ ( .D(n1927), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(iwb_adr_o[9]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_9_ ( .D(n1928), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(iwb_adr_o[10]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_10_ ( .D(n1929), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(iwb_adr_o[11]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_11_ ( .D(n1930), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(iwb_adr_o[12]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_12_ ( .D(n1931), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(iwb_adr_o[13]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_13_ ( .D(n1932), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(iwb_adr_o[14]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_5_ ( .D(n1924), .CKN(wb_clk_o), .R(n2810), 
        .SN(n3), .Q(iwb_adr_o[6]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_14_ ( .D(n1933), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(iwb_adr_o[15]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_15_ ( .D(n1934), .CKN(wb_clk_o), .R(n2816), 
        .SN(n3), .Q(iwb_adr_o[16]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_16_ ( .D(n1935), .CKN(wb_clk_o), .R(n2815), 
        .SN(n3), .Q(iwb_adr_o[17]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_3_ ( .D(n1961), .CKN(wb_clk_o), .R(n2813), 
        .SN(n3), .Q(iwb_adr_o[4]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_2_ ( .D(n1962), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(iwb_adr_o[3]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_0_ ( .D(n2038), .CK(wb_clk_o), .R(n2796), .Q(
        rfsr0h[0]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_4_ ( .D(n2714), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[4]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_1_ ( .D(n2021), .CK(wb_clk_o), .R(n2793), .Q(
        rfsr1h[1]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_2_ ( .D(n2020), .CK(wb_clk_o), .R(n2804), .Q(
        rfsr1h[2]) );
  DFFRPQ_X1M_A12TR rfsr1h_reg_0_ ( .D(n2022), .CK(wb_clk_o), .R(n2793), .Q(
        rfsr1h[0]) );
  DFFRPQ_X1M_A12TR rfsr2h_reg_2_ ( .D(n2012), .CK(wb_clk_o), .R(n2795), .Q(
        rfsr2h[2]) );
  DFFRPQ_X1M_A12TR rfsr2h_reg_1_ ( .D(n2013), .CK(wb_clk_o), .R(n2795), .Q(
        rfsr2h[1]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_1_ ( .D(n2037), .CK(wb_clk_o), .R(n2805), .Q(
        rfsr0h[1]) );
  DFFRPQ_X1M_A12TR rfsr0h_reg_2_ ( .D(n2036), .CK(wb_clk_o), .R(n2805), .Q(
        rfsr0h[2]) );
  DFFRPQ_X1M_A12TR rfsr2h_reg_0_ ( .D(n2014), .CK(wb_clk_o), .R(n2795), .Q(
        rfsr2h[0]) );
  DFFRPQ_X1M_A12TR rtblptrl_reg_0_ ( .D(n1990), .CK(wb_clk_o), .R(n2795), .Q(
        wtblat[0]) );
  DFFNSRPQ_X1M_A12TR rreset_reg ( .D(rreset_), .CKN(wb_clk_o), .R(n4431), .SN(
        n3), .Q(qrst) );
  DFFNSRPQ_X1M_A12TR rireg_reg_3_ ( .D(n2715), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[3]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_2_ ( .D(n2716), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[2]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_1_ ( .D(n2717), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[1]) );
  DFFRPQ_X1M_A12TR rwreg_reg_0_ ( .D(n1560), .CK(wb_clk_o), .R(n2799), .Q(
        rwreg[0]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_1_ ( .D(n1885), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(rsrc[1]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_4_ ( .D(n1879), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(rsrc[4]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_2_ ( .D(n1868), .CKN(wb_clk_o), .R(n2813), .SN(
        n3), .Q(rsrc[2]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_3_ ( .D(n1853), .CKN(wb_clk_o), .R(n2810), .SN(
        n3), .Q(rsrc[3]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_6_ ( .D(n1835), .CKN(wb_clk_o), .R(n2807), .SN(
        n3), .Q(rsrc[6]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_5_ ( .D(n1636), .CKN(wb_clk_o), .R(n2812), .SN(
        n3), .Q(rsrc[5]) );
  DFFRPQ_X1M_A12TR rfsr1l_reg_0_ ( .D(n2030), .CK(wb_clk_o), .R(n2793), .Q(
        rfsr1l[0]) );
  DFFRPQ_X1M_A12TR rfsr2l_reg_0_ ( .D(n2053), .CK(wb_clk_o), .R(n2794), .Q(
        rfsr2l[0]) );
  DFFRPQ_X1M_A12TR rfsr0l_reg_0_ ( .D(n2046), .CK(wb_clk_o), .R(n2794), .Q(
        rfsr0l[0]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_0_ ( .D(n2718), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[0]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_0_ ( .D(n1901), .CKN(wb_clk_o), .R(n2811), .SN(
        n3), .Q(rsrc[0]) );
  DFFNSRPQ_X1M_A12TR rsrc_reg_7_ ( .D(n1893), .CKN(wb_clk_o), .R(n2810), .SN(
        n3), .Q(rsrc[7]) );
  DFFNSRPQ_X1M_A12TR riwbadr_reg_0_ ( .D(n1921), .CKN(wb_clk_o), .R(n2817), 
        .SN(n3), .Q(iwb_adr_o[1]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_6_ ( .D(n1582), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rtgt[6]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_5_ ( .D(n1578), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rtgt[5]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_3_ ( .D(n1570), .CKN(wb_clk_o), .R(n2817), .SN(
        n3), .Q(rtgt[3]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_2_ ( .D(n1566), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rtgt[2]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_1_ ( .D(n1562), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rtgt[1]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_4_ ( .D(n1574), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rtgt[4]) );
  DFFNSRPQ_X1M_A12TR rqclk_reg_1_ ( .D(n1803), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(qena[1]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_7_ ( .D(n1586), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(rtgt[7]) );
  DFFRPQ_X1M_A12TR rtosu_reg_3_ ( .D(n1854), .CK(wb_clk_o), .R(n2803), .Q(
        wstkw[19]) );
  DFFRPQ_X1M_A12TR rtosu_reg_1_ ( .D(n1420), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[17]) );
  DFFRPQ_X1M_A12TR rtosu_reg_2_ ( .D(n1416), .CK(wb_clk_o), .R(n2803), .Q(
        wstkw[18]) );
  DFFRPQ_X1M_A12TR rtosl_reg_4_ ( .D(n1553), .CK(wb_clk_o), .R(n2800), .Q(
        wstkw[4]) );
  DFFRPQ_X1M_A12TR rtosl_reg_0_ ( .D(n4432), .CK(wb_clk_o), .R(n2805), .Q(
        wstkw[0]) );
  DFFRPQ_X1M_A12TR rtosl_reg_5_ ( .D(n1592), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[5]) );
  DFFRPQ_X1M_A12TR rtosh_reg_6_ ( .D(n1836), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[14]) );
  DFFRPQ_X1M_A12TR rtosh_reg_4_ ( .D(n1538), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[12]) );
  DFFRPQ_X1M_A12TR rtosh_reg_3_ ( .D(n1532), .CK(wb_clk_o), .R(n2799), .Q(
        wstkw[11]) );
  DFFRPQ_X1M_A12TR rtosh_reg_2_ ( .D(n1526), .CK(wb_clk_o), .R(n2801), .Q(
        wstkw[10]) );
  DFFRPQ_X1M_A12TR rtosh_reg_1_ ( .D(n1520), .CK(wb_clk_o), .R(n2806), .Q(
        wstkw[9]) );
  DFFRPQ_X1M_A12TR rtosh_reg_7_ ( .D(n1434), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[15]) );
  DFFRPQ_X1M_A12TR rtosl_reg_2_ ( .D(n1862), .CK(wb_clk_o), .R(n2804), .Q(
        wstkw[2]) );
  DFFRPQ_X1M_A12TR rtosl_reg_3_ ( .D(n1847), .CK(wb_clk_o), .R(n2801), .Q(
        wstkw[3]) );
  DFFRPQ_X1M_A12TR rtosl_reg_7_ ( .D(n1595), .CK(wb_clk_o), .R(n2800), .Q(
        wstkw[7]) );
  DFFRPQ_X1M_A12TR rtosl_reg_1_ ( .D(n1589), .CK(wb_clk_o), .R(n2804), .Q(
        wstkw[1]) );
  DFFRPQ_X1M_A12TR rtosh_reg_5_ ( .D(n1544), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[13]) );
  DFFRPQ_X1M_A12TR rtosh_reg_0_ ( .D(n1514), .CK(wb_clk_o), .R(n2801), .Q(
        wstkw[8]) );
  DFFRPQ_X1M_A12TR rtosl_reg_6_ ( .D(n1444), .CK(wb_clk_o), .R(n2803), .Q(
        wstkw[6]) );
  DFFRPQ_X1M_A12TR rtosu_reg_0_ ( .D(n1427), .CK(wb_clk_o), .R(n2802), .Q(
        wstkw[16]) );
  DFFNSRPQ_X1M_A12TR rtgt_reg_0_ ( .D(n1497), .CKN(wb_clk_o), .R(n2820), .SN(
        n3), .Q(wneg[0]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_10_ ( .D(n2708), .CKN(wb_clk_o), .R(n2823), 
        .SN(n3), .Q(rireg[10]) );
  DFFNSRPQ_X1M_A12TR rqclk_reg_3_ ( .D(n1807), .CKN(wb_clk_o), .R(iwb_adr_o[0]), .SN(qrst), .Q(qena[3]) );
  DFFNSRPQ_X1M_A12TR rireg_reg_7_ ( .D(n2711), .CKN(wb_clk_o), .R(n2822), .SN(
        n3), .Q(rireg[7]) );
  DFFRPQ_X1M_A12TR rstkptr_reg_4_ ( .D(n1650), .CK(wb_clk_o), .R(n2803), .Q(
        n218) );
  DFFRPQ_X1M_A12TR rstkptr_reg_2_ ( .D(n1869), .CK(wb_clk_o), .R(n2803), .Q(
        n216) );
  DFFRPQ_X1M_A12TR rstkptr_reg_3_ ( .D(n1651), .CK(wb_clk_o), .R(n2791), .Q(
        n217) );
  ADDH_X1M_A12TR add_1310_u1_1_4 ( .A(n218), .B(add_1310_carry[4]), .CO(
        add_1310_carry[5]), .S(wstkinc[4]) );
  ADDH_X1M_A12TR add_1310_u1_1_2 ( .A(n216), .B(add_1310_carry[2]), .CO(
        add_1310_carry[3]), .S(wstkinc[2]) );
  ADDH_X1M_A12TR add_1310_u1_1_3 ( .A(n217), .B(add_1310_carry[3]), .CO(
        add_1310_carry[4]), .S(wstkinc[3]) );
  ADDH_X1M_A12TR add_1310_u1_1_1 ( .A(n215), .B(n214), .CO(add_1310_carry[2]), 
        .S(wstkinc[1]) );
  DFFNSRPQ_X1M_A12TR rreset__reg ( .D(n2745), .CKN(wb_clk_o), .R(n4431), .SN(
        n3), .Q(rreset_) );
  DFFRPQ_X3M_A12TR rstkptr_reg_0_ ( .D(n1871), .CK(wb_clk_o), .R(n2791), .Q(
        n214) );
  XNOR2_X1M_A12TR u2736 ( .A(rstkptr_5_), .B(n2848), .Y(n2746) );
  MXT2_X1M_A12TR u2737 ( .A(n2876), .B(n2871), .S0(n218), .Y(n2747) );
  MXT2_X1M_A12TR u2738 ( .A(n2886), .B(n2881), .S0(n218), .Y(n2748) );
  MXT2_X1M_A12TR u2739 ( .A(n2996), .B(n2991), .S0(n218), .Y(n2749) );
  MXT2_X1M_A12TR u2740 ( .A(n2926), .B(n2921), .S0(n218), .Y(n2750) );
  MXT2_X1M_A12TR u2741 ( .A(n2866), .B(n2861), .S0(n218), .Y(n2751) );
  MXT2_X1M_A12TR u2742 ( .A(n2986), .B(n2981), .S0(n218), .Y(n2752) );
  MXT2_X1M_A12TR u2743 ( .A(n2976), .B(n2971), .S0(n218), .Y(n2753) );
  MXT2_X1M_A12TR u2744 ( .A(n2966), .B(n2961), .S0(n218), .Y(n2754) );
  MXT2_X1M_A12TR u2745 ( .A(n2956), .B(n2951), .S0(n218), .Y(n2755) );
  MXT2_X1M_A12TR u2746 ( .A(n2946), .B(n2941), .S0(n218), .Y(n2756) );
  MXT2_X1M_A12TR u2747 ( .A(n2936), .B(n2931), .S0(n218), .Y(n2757) );
  MXT2_X1M_A12TR u2748 ( .A(n2916), .B(n2911), .S0(n218), .Y(n2758) );
  MXT2_X1M_A12TR u2749 ( .A(n3006), .B(n3001), .S0(n218), .Y(n2759) );
  MXT2_X1M_A12TR u2750 ( .A(n3016), .B(n3011), .S0(n218), .Y(n2760) );
  BUFH_X1M_A12TR u2751 ( .A(n2838), .Y(n2798) );
  BUFH_X1M_A12TR u2752 ( .A(n2840), .Y(n2793) );
  BUFH_X1M_A12TR u2753 ( .A(n2839), .Y(n2796) );
  BUFH_X1M_A12TR u2754 ( .A(n2837), .Y(n2799) );
  BUFH_X1M_A12TR u2755 ( .A(n2841), .Y(n2792) );
  BUFH_X1M_A12TR u2756 ( .A(n2839), .Y(n2795) );
  BUFH_X1M_A12TR u2757 ( .A(n2836), .Y(n2802) );
  BUFH_X1M_A12TR u2758 ( .A(n2835), .Y(n2804) );
  BUFH_X1M_A12TR u2759 ( .A(n2835), .Y(n2803) );
  BUFH_X1M_A12TR u2760 ( .A(n2841), .Y(n2791) );
  BUFH_X1M_A12TR u2761 ( .A(n2838), .Y(n2797) );
  BUFH_X1M_A12TR u2762 ( .A(n2834), .Y(n2805) );
  BUFH_X1M_A12TR u2763 ( .A(n2840), .Y(n2794) );
  BUFH_X1M_A12TR u2764 ( .A(n2836), .Y(n2801) );
  BUFH_X1M_A12TR u2765 ( .A(n2837), .Y(n2800) );
  BUFH_X1M_A12TR u2766 ( .A(n2834), .Y(n2806) );
  BUFH_X1M_A12TR u2767 ( .A(n2828), .Y(n2818) );
  BUFH_X1M_A12TR u2768 ( .A(n2833), .Y(n2808) );
  BUFH_X1M_A12TR u2769 ( .A(n2827), .Y(n2820) );
  BUFH_X1M_A12TR u2770 ( .A(n2827), .Y(n2819) );
  BUFH_X1M_A12TR u2771 ( .A(n2833), .Y(n2807) );
  BUFH_X1M_A12TR u2772 ( .A(n2829), .Y(n2816) );
  BUFH_X1M_A12TR u2773 ( .A(n2829), .Y(n2815) );
  BUFH_X1M_A12TR u2774 ( .A(n2832), .Y(n2809) );
  BUFH_X1M_A12TR u2775 ( .A(n2830), .Y(n2813) );
  BUFH_X1M_A12TR u2776 ( .A(n2828), .Y(n2817) );
  BUFH_X1M_A12TR u2777 ( .A(n2831), .Y(n2812) );
  BUFH_X1M_A12TR u2778 ( .A(n2832), .Y(n2810) );
  BUFH_X1M_A12TR u2779 ( .A(n2831), .Y(n2811) );
  BUFH_X1M_A12TR u2780 ( .A(n2830), .Y(n2814) );
  BUFH_X1M_A12TR u2781 ( .A(n2826), .Y(n2821) );
  BUFH_X1M_A12TR u2782 ( .A(n2826), .Y(n2822) );
  BUFH_X1M_A12TR u2783 ( .A(n2825), .Y(n2823) );
  BUFH_X1M_A12TR u2784 ( .A(n2825), .Y(wb_rst_o) );
  BUFH_X1M_A12TR u2785 ( .A(n2846), .Y(n2827) );
  BUFH_X1M_A12TR u2786 ( .A(n2842), .Y(n2839) );
  BUFH_X1M_A12TR u2787 ( .A(n2844), .Y(n2833) );
  BUFH_X1M_A12TR u2788 ( .A(n2846), .Y(n2829) );
  BUFH_X1M_A12TR u2789 ( .A(n2844), .Y(n2835) );
  BUFH_X1M_A12TR u2790 ( .A(n2842), .Y(n2841) );
  BUFH_X1M_A12TR u2791 ( .A(n2843), .Y(n2838) );
  BUFH_X1M_A12TR u2792 ( .A(n2844), .Y(n2834) );
  BUFH_X1M_A12TR u2793 ( .A(n2846), .Y(n2828) );
  BUFH_X1M_A12TR u2794 ( .A(n2842), .Y(n2840) );
  BUFH_X1M_A12TR u2795 ( .A(n2845), .Y(n2832) );
  BUFH_X1M_A12TR u2796 ( .A(n2843), .Y(n2836) );
  BUFH_X1M_A12TR u2797 ( .A(n2845), .Y(n2831) );
  BUFH_X1M_A12TR u2798 ( .A(n2843), .Y(n2837) );
  BUFH_X1M_A12TR u2799 ( .A(n2845), .Y(n2830) );
  BUFH_X1M_A12TR u2800 ( .A(n2847), .Y(n2826) );
  BUFH_X1M_A12TR u2801 ( .A(n2847), .Y(n2825) );
  XOR2_X1M_A12TR u2802 ( .A(wsub[5]), .B(n2770), .Y(wsubc[5]) );
  XOR2_X1M_A12TR u2803 ( .A(n4428), .B(n2764), .Y(wneg[5]) );
  XOR2_X1M_A12TR u2804 ( .A(wsub[6]), .B(n2771), .Y(wsubc[6]) );
  XOR2_X1M_A12TR u2805 ( .A(n4429), .B(n2765), .Y(wneg[6]) );
  XOR2_X1M_A12TR u2806 ( .A(wsub[3]), .B(n2768), .Y(wsubc[3]) );
  XOR2_X1M_A12TR u2807 ( .A(n4426), .B(n2762), .Y(wneg[3]) );
  XOR2_X1M_A12TR u2808 ( .A(wsub[2]), .B(n2767), .Y(wsubc[2]) );
  XOR2_X1M_A12TR u2809 ( .A(n4425), .B(n2761), .Y(wneg[2]) );
  XOR2_X1M_A12TR u2810 ( .A(wsub[4]), .B(n2769), .Y(wsubc[4]) );
  XOR2_X1M_A12TR u2811 ( .A(n4427), .B(n2763), .Y(wneg[4]) );
  XOR2_X1M_A12TR u2812 ( .A(wsub[1]), .B(n2790), .Y(wsubc[1]) );
  XOR2_X1M_A12TR u2813 ( .A(n4424), .B(n4423), .Y(wneg[1]) );
  XOR2_X1M_A12TR u2814 ( .A(wsub[7]), .B(n2772), .Y(wsubc[7]) );
  XOR2_X1M_A12TR u2815 ( .A(n4430), .B(n2766), .Y(wneg[7]) );
  BUFH_X1M_A12TR u2816 ( .A(n4433), .Y(n2844) );
  BUFH_X1M_A12TR u2817 ( .A(n4433), .Y(n2846) );
  BUFH_X1M_A12TR u2818 ( .A(n4433), .Y(n2842) );
  BUFH_X1M_A12TR u2819 ( .A(n4433), .Y(n2843) );
  BUFH_X1M_A12TR u2820 ( .A(n4433), .Y(n2845) );
  BUFH_X1M_A12TR u2821 ( .A(n4433), .Y(n2847) );
  XNOR2_X1M_A12TR u2822 ( .A(wadd[8]), .B(n2850), .Y(waddc[8]) );
  NAND2_X1M_A12TR u2823 ( .A(n2778), .B(wadd[7]), .Y(n2850) );
  XOR2_X1M_A12TR u2824 ( .A(wadd[1]), .B(n2789), .Y(waddc[1]) );
  XOR2_X1M_A12TR u2825 ( .A(wadd[5]), .B(n2776), .Y(waddc[5]) );
  XOR2_X1M_A12TR u2826 ( .A(wadd[6]), .B(n2777), .Y(waddc[6]) );
  XOR2_X1M_A12TR u2827 ( .A(wadd[3]), .B(n2774), .Y(waddc[3]) );
  XOR2_X1M_A12TR u2828 ( .A(wadd[2]), .B(n2773), .Y(waddc[2]) );
  XOR2_X1M_A12TR u2829 ( .A(wadd[4]), .B(n2775), .Y(waddc[4]) );
  XOR2_X1M_A12TR u2830 ( .A(wadd[7]), .B(n2778), .Y(waddc[7]) );
  XNOR2_X1M_A12TR u2831 ( .A(wsub[8]), .B(n2849), .Y(wsubc[8]) );
  NAND2_X1M_A12TR u2832 ( .A(n2772), .B(wsub[7]), .Y(n2849) );
  AND2_X1M_A12TR u2833 ( .A(n4423), .B(n4424), .Y(n2761) );
  AND2_X1M_A12TR u2834 ( .A(n2761), .B(n4425), .Y(n2762) );
  AND2_X1M_A12TR u2835 ( .A(n2762), .B(n4426), .Y(n2763) );
  AND2_X1M_A12TR u2836 ( .A(n2763), .B(n4427), .Y(n2764) );
  AND2_X1M_A12TR u2837 ( .A(n2764), .B(n4428), .Y(n2765) );
  AND2_X1M_A12TR u2838 ( .A(n2765), .B(n4429), .Y(n2766) );
  AND2_X1M_A12TR u2839 ( .A(n2790), .B(wsub[1]), .Y(n2767) );
  AND2_X1M_A12TR u2840 ( .A(n2767), .B(wsub[2]), .Y(n2768) );
  AND2_X1M_A12TR u2841 ( .A(n2768), .B(wsub[3]), .Y(n2769) );
  AND2_X1M_A12TR u2842 ( .A(n2769), .B(wsub[4]), .Y(n2770) );
  AND2_X1M_A12TR u2843 ( .A(n2770), .B(wsub[5]), .Y(n2771) );
  AND2_X1M_A12TR u2844 ( .A(n2771), .B(wsub[6]), .Y(n2772) );
  AND2_X1M_A12TR u2845 ( .A(n2789), .B(wadd[1]), .Y(n2773) );
  AND2_X1M_A12TR u2846 ( .A(n2773), .B(wadd[2]), .Y(n2774) );
  AND2_X1M_A12TR u2847 ( .A(n2774), .B(wadd[3]), .Y(n2775) );
  AND2_X1M_A12TR u2848 ( .A(n2775), .B(wadd[4]), .Y(n2776) );
  AND2_X1M_A12TR u2849 ( .A(n2776), .B(wadd[5]), .Y(n2777) );
  AND2_X1M_A12TR u2850 ( .A(n2777), .B(wadd[6]), .Y(n2778) );
  AND2_X1M_A12TR u2851 ( .A(n2766), .B(n4430), .Y(n2779) );
  XNOR2_X1M_A12TR u2852 ( .A(n215), .B(n214), .Y(wstkdec[1]) );
  XNOR2_X1M_A12TR u2853 ( .A(wrrc_7_), .B(wsub[0]), .Y(wsubc[0]) );
  MXT2_X1M_A12TR u2854 ( .A(n3036), .B(n3031), .S0(n218), .Y(n2780) );
  MXT2_X1M_A12TR u2855 ( .A(n3026), .B(n3021), .S0(n218), .Y(n2781) );
  MXT2_X1M_A12TR u2856 ( .A(n3046), .B(n3041), .S0(n218), .Y(n2782) );
  NAND2XB_X1M_A12TR u2857 ( .BN(n3051), .A(n3069), .Y(n3068) );
  MXT2_X1M_A12TR u2858 ( .A(n2896), .B(n2891), .S0(n218), .Y(n2783) );
  MXT2_X1M_A12TR u2859 ( .A(n2906), .B(n2901), .S0(n218), .Y(n2784) );
  XOR2_X1M_A12TR u2860 ( .A(rireg[0]), .B(iwb_adr_o[1]), .Y(n366) );
  XNOR2_X1M_A12TR u2861 ( .A(n217), .B(n2788), .Y(wstkdec[3]) );
  MXIT2_X0P7M_A12TR u2862 ( .A(n2856), .B(n2851), .S0(n218), .Y(n3051) );
  MXIT4_X1M_A12TR u2863 ( .A(n2857), .B(n2858), .C(n2859), .D(n2860), .S0(n217), .S1(n216), .Y(n2856) );
  MXIT4_X1M_A12TR u2864 ( .A(n2852), .B(n2853), .C(n2854), .D(n2855), .S0(n217), .S1(n216), .Y(n2851) );
  MXIT4_X1M_A12TR u2865 ( .A(rstkram[380]), .B(rstkram[340]), .C(rstkram[360]), 
        .D(rstkram[320]), .S0(n215), .S1(n214), .Y(n2860) );
  MXIT4_X1M_A12TR u2866 ( .A(n3017), .B(n3018), .C(n3019), .D(n3020), .S0(n217), .S1(n216), .Y(n3016) );
  MXIT4_X1M_A12TR u2867 ( .A(n3012), .B(n3013), .C(n3014), .D(n3015), .S0(n217), .S1(n216), .Y(n3011) );
  MXIT4_X1M_A12TR u2868 ( .A(rstkram[396]), .B(rstkram[356]), .C(rstkram[376]), 
        .D(rstkram[336]), .S0(n215), .S1(n214), .Y(n3020) );
  MXIT4_X1M_A12TR u2869 ( .A(n3007), .B(n3008), .C(n3009), .D(n3010), .S0(n217), .S1(n216), .Y(n3006) );
  MXIT4_X1M_A12TR u2870 ( .A(n3002), .B(n3003), .C(n3004), .D(n3005), .S0(n217), .S1(n216), .Y(n3001) );
  MXIT4_X1M_A12TR u2871 ( .A(rstkram[395]), .B(rstkram[355]), .C(rstkram[375]), 
        .D(rstkram[335]), .S0(n215), .S1(n214), .Y(n3010) );
  MXIT4_X1M_A12TR u2872 ( .A(n2917), .B(n2918), .C(n2919), .D(n2920), .S0(n217), .S1(n216), .Y(n2916) );
  MXIT4_X1M_A12TR u2873 ( .A(n2912), .B(n2913), .C(n2914), .D(n2915), .S0(n217), .S1(n216), .Y(n2911) );
  MXIT4_X1M_A12TR u2874 ( .A(rstkram[386]), .B(rstkram[346]), .C(rstkram[366]), 
        .D(rstkram[326]), .S0(n215), .S1(n214), .Y(n2920) );
  MXIT4_X1M_A12TR u2875 ( .A(n2937), .B(n2938), .C(n2939), .D(n2940), .S0(n217), .S1(n216), .Y(n2936) );
  MXIT4_X1M_A12TR u2876 ( .A(n2932), .B(n2933), .C(n2934), .D(n2935), .S0(n217), .S1(n216), .Y(n2931) );
  MXIT4_X1M_A12TR u2877 ( .A(rstkram[388]), .B(rstkram[348]), .C(rstkram[368]), 
        .D(rstkram[328]), .S0(n215), .S1(n214), .Y(n2940) );
  MXIT4_X1M_A12TR u2878 ( .A(n2947), .B(n2948), .C(n2949), .D(n2950), .S0(n217), .S1(n216), .Y(n2946) );
  MXIT4_X1M_A12TR u2879 ( .A(n2942), .B(n2943), .C(n2944), .D(n2945), .S0(n217), .S1(n216), .Y(n2941) );
  MXIT4_X1M_A12TR u2880 ( .A(rstkram[389]), .B(rstkram[349]), .C(rstkram[369]), 
        .D(rstkram[329]), .S0(n215), .S1(n214), .Y(n2950) );
  MXIT4_X1M_A12TR u2881 ( .A(n2957), .B(n2958), .C(n2959), .D(n2960), .S0(n217), .S1(n216), .Y(n2956) );
  MXIT4_X1M_A12TR u2882 ( .A(n2952), .B(n2953), .C(n2954), .D(n2955), .S0(n217), .S1(n216), .Y(n2951) );
  MXIT4_X1M_A12TR u2883 ( .A(rstkram[390]), .B(rstkram[350]), .C(rstkram[370]), 
        .D(rstkram[330]), .S0(n215), .S1(n214), .Y(n2960) );
  MXIT4_X1M_A12TR u2884 ( .A(n2967), .B(n2968), .C(n2969), .D(n2970), .S0(n217), .S1(n216), .Y(n2966) );
  MXIT4_X1M_A12TR u2885 ( .A(n2962), .B(n2963), .C(n2964), .D(n2965), .S0(n217), .S1(n216), .Y(n2961) );
  MXIT4_X1M_A12TR u2886 ( .A(rstkram[391]), .B(rstkram[351]), .C(rstkram[371]), 
        .D(rstkram[331]), .S0(n215), .S1(n214), .Y(n2970) );
  MXIT4_X1M_A12TR u2887 ( .A(n2977), .B(n2978), .C(n2979), .D(n2980), .S0(n217), .S1(n216), .Y(n2976) );
  MXIT4_X1M_A12TR u2888 ( .A(n2972), .B(n2973), .C(n2974), .D(n2975), .S0(n217), .S1(n216), .Y(n2971) );
  MXIT4_X1M_A12TR u2889 ( .A(rstkram[392]), .B(rstkram[352]), .C(rstkram[372]), 
        .D(rstkram[332]), .S0(n215), .S1(n214), .Y(n2980) );
  MXIT4_X1M_A12TR u2890 ( .A(n2987), .B(n2988), .C(n2989), .D(n2990), .S0(n217), .S1(n216), .Y(n2986) );
  MXIT4_X1M_A12TR u2891 ( .A(n2982), .B(n2983), .C(n2984), .D(n2985), .S0(n217), .S1(n216), .Y(n2981) );
  MXIT4_X1M_A12TR u2892 ( .A(rstkram[393]), .B(rstkram[353]), .C(rstkram[373]), 
        .D(rstkram[333]), .S0(n215), .S1(n214), .Y(n2990) );
  MXIT4_X1M_A12TR u2893 ( .A(n2867), .B(n2868), .C(n2869), .D(n2870), .S0(n217), .S1(n216), .Y(n2866) );
  MXIT4_X1M_A12TR u2894 ( .A(n2862), .B(n2863), .C(n2864), .D(n2865), .S0(n217), .S1(n216), .Y(n2861) );
  MXIT4_X1M_A12TR u2895 ( .A(rstkram[381]), .B(rstkram[341]), .C(rstkram[361]), 
        .D(rstkram[321]), .S0(n215), .S1(n214), .Y(n2870) );
  MXIT4_X1M_A12TR u2896 ( .A(n2927), .B(n2928), .C(n2929), .D(n2930), .S0(n217), .S1(n216), .Y(n2926) );
  MXIT4_X1M_A12TR u2897 ( .A(n2922), .B(n2923), .C(n2924), .D(n2925), .S0(n217), .S1(n216), .Y(n2921) );
  MXIT4_X1M_A12TR u2898 ( .A(rstkram[387]), .B(rstkram[347]), .C(rstkram[367]), 
        .D(rstkram[327]), .S0(n215), .S1(n214), .Y(n2930) );
  MXIT4_X1M_A12TR u2899 ( .A(n2997), .B(n2998), .C(n2999), .D(n3000), .S0(n217), .S1(n216), .Y(n2996) );
  MXIT4_X1M_A12TR u2900 ( .A(n2992), .B(n2993), .C(n2994), .D(n2995), .S0(n217), .S1(n216), .Y(n2991) );
  MXIT4_X1M_A12TR u2901 ( .A(rstkram[394]), .B(rstkram[354]), .C(rstkram[374]), 
        .D(rstkram[334]), .S0(n215), .S1(n214), .Y(n3000) );
  MXIT4_X1M_A12TR u2902 ( .A(n2887), .B(n2888), .C(n2889), .D(n2890), .S0(n217), .S1(n216), .Y(n2886) );
  MXIT4_X1M_A12TR u2903 ( .A(n2882), .B(n2883), .C(n2884), .D(n2885), .S0(n217), .S1(n216), .Y(n2881) );
  MXIT4_X1M_A12TR u2904 ( .A(rstkram[383]), .B(rstkram[343]), .C(rstkram[363]), 
        .D(rstkram[323]), .S0(n215), .S1(n214), .Y(n2890) );
  MXIT4_X1M_A12TR u2905 ( .A(n2877), .B(n2878), .C(n2879), .D(n2880), .S0(n217), .S1(n216), .Y(n2876) );
  MXIT4_X1M_A12TR u2906 ( .A(n2872), .B(n2873), .C(n2874), .D(n2875), .S0(n217), .S1(n216), .Y(n2871) );
  MXIT4_X1M_A12TR u2907 ( .A(rstkram[382]), .B(rstkram[342]), .C(rstkram[362]), 
        .D(rstkram[322]), .S0(n215), .S1(n214), .Y(n2880) );
  XNOR2_X1M_A12TR u2908 ( .A(n216), .B(n2785), .Y(wstkdec[2]) );
  XOR2_X1M_A12TR u2909 ( .A(wrrc_7_), .B(wadd[0]), .Y(waddc[0]) );
  OR2_X1M_A12TR u2910 ( .A(n214), .B(n215), .Y(n2785) );
  XNOR2_X1M_A12TR u2911 ( .A(n218), .B(n2787), .Y(wstkdec[4]) );
  MXIT4_X1M_A12TR u2912 ( .A(rstkram[140]), .B(rstkram[100]), .C(rstkram[120]), 
        .D(rstkram[80]), .S0(n215), .S1(n214), .Y(n2853) );
  MXIT4_X1M_A12TR u2913 ( .A(rstkram[460]), .B(rstkram[420]), .C(rstkram[440]), 
        .D(rstkram[400]), .S0(n215), .S1(n214), .Y(n2858) );
  MXIT4_X1M_A12TR u2914 ( .A(rstkram[158]), .B(rstkram[118]), .C(rstkram[138]), 
        .D(rstkram[98]), .S0(n215), .S1(n214), .Y(n3033) );
  MXIT4_X1M_A12TR u2915 ( .A(rstkram[478]), .B(rstkram[438]), .C(rstkram[458]), 
        .D(rstkram[418]), .S0(n215), .S1(n214), .Y(n3038) );
  MXIT4_X1M_A12TR u2916 ( .A(rstkram[157]), .B(rstkram[117]), .C(rstkram[137]), 
        .D(rstkram[97]), .S0(n215), .S1(n214), .Y(n3023) );
  MXIT4_X1M_A12TR u2917 ( .A(rstkram[477]), .B(rstkram[437]), .C(rstkram[457]), 
        .D(rstkram[417]), .S0(n215), .S1(n214), .Y(n3028) );
  MXIT4_X1M_A12TR u2918 ( .A(rstkram[156]), .B(rstkram[116]), .C(rstkram[136]), 
        .D(rstkram[96]), .S0(n215), .S1(n214), .Y(n3013) );
  MXIT4_X1M_A12TR u2919 ( .A(rstkram[476]), .B(rstkram[436]), .C(rstkram[456]), 
        .D(rstkram[416]), .S0(n215), .S1(n214), .Y(n3018) );
  MXIT4_X1M_A12TR u2920 ( .A(rstkram[155]), .B(rstkram[115]), .C(rstkram[135]), 
        .D(rstkram[95]), .S0(n215), .S1(n214), .Y(n3003) );
  MXIT4_X1M_A12TR u2921 ( .A(rstkram[475]), .B(rstkram[435]), .C(rstkram[455]), 
        .D(rstkram[415]), .S0(n215), .S1(n214), .Y(n3008) );
  MXIT4_X1M_A12TR u2922 ( .A(rstkram[146]), .B(rstkram[106]), .C(rstkram[126]), 
        .D(rstkram[86]), .S0(n215), .S1(n214), .Y(n2913) );
  MXIT4_X1M_A12TR u2923 ( .A(rstkram[466]), .B(rstkram[426]), .C(rstkram[446]), 
        .D(rstkram[406]), .S0(n215), .S1(n214), .Y(n2918) );
  MXIT4_X1M_A12TR u2924 ( .A(rstkram[148]), .B(rstkram[108]), .C(rstkram[128]), 
        .D(rstkram[88]), .S0(n215), .S1(n214), .Y(n2933) );
  MXIT4_X1M_A12TR u2925 ( .A(rstkram[468]), .B(rstkram[428]), .C(rstkram[448]), 
        .D(rstkram[408]), .S0(n215), .S1(n214), .Y(n2938) );
  MXIT4_X1M_A12TR u2926 ( .A(rstkram[149]), .B(rstkram[109]), .C(rstkram[129]), 
        .D(rstkram[89]), .S0(n215), .S1(n214), .Y(n2943) );
  MXIT4_X1M_A12TR u2927 ( .A(rstkram[469]), .B(rstkram[429]), .C(rstkram[449]), 
        .D(rstkram[409]), .S0(n215), .S1(n214), .Y(n2948) );
  MXIT4_X1M_A12TR u2928 ( .A(rstkram[150]), .B(rstkram[110]), .C(rstkram[130]), 
        .D(rstkram[90]), .S0(n215), .S1(n214), .Y(n2953) );
  MXIT4_X1M_A12TR u2929 ( .A(rstkram[470]), .B(rstkram[430]), .C(rstkram[450]), 
        .D(rstkram[410]), .S0(n215), .S1(n214), .Y(n2958) );
  MXIT4_X1M_A12TR u2930 ( .A(rstkram[151]), .B(rstkram[111]), .C(rstkram[131]), 
        .D(rstkram[91]), .S0(n215), .S1(n214), .Y(n2963) );
  MXIT4_X1M_A12TR u2931 ( .A(rstkram[471]), .B(rstkram[431]), .C(rstkram[451]), 
        .D(rstkram[411]), .S0(n215), .S1(n214), .Y(n2968) );
  MXIT4_X1M_A12TR u2932 ( .A(rstkram[152]), .B(rstkram[112]), .C(rstkram[132]), 
        .D(rstkram[92]), .S0(n215), .S1(n214), .Y(n2973) );
  MXIT4_X1M_A12TR u2933 ( .A(rstkram[472]), .B(rstkram[432]), .C(rstkram[452]), 
        .D(rstkram[412]), .S0(n215), .S1(n214), .Y(n2978) );
  MXIT4_X1M_A12TR u2934 ( .A(rstkram[153]), .B(rstkram[113]), .C(rstkram[133]), 
        .D(rstkram[93]), .S0(n215), .S1(n214), .Y(n2983) );
  MXIT4_X1M_A12TR u2935 ( .A(rstkram[473]), .B(rstkram[433]), .C(rstkram[453]), 
        .D(rstkram[413]), .S0(n215), .S1(n214), .Y(n2988) );
  MXIT4_X1M_A12TR u2936 ( .A(rstkram[144]), .B(rstkram[104]), .C(rstkram[124]), 
        .D(rstkram[84]), .S0(n215), .S1(n214), .Y(n2893) );
  MXIT4_X1M_A12TR u2937 ( .A(rstkram[464]), .B(rstkram[424]), .C(rstkram[444]), 
        .D(rstkram[404]), .S0(n215), .S1(n214), .Y(n2898) );
  MXIT4_X1M_A12TR u2938 ( .A(rstkram[141]), .B(rstkram[101]), .C(rstkram[121]), 
        .D(rstkram[81]), .S0(n215), .S1(n214), .Y(n2863) );
  MXIT4_X1M_A12TR u2939 ( .A(rstkram[461]), .B(rstkram[421]), .C(rstkram[441]), 
        .D(rstkram[401]), .S0(n215), .S1(n214), .Y(n2868) );
  MXIT4_X1M_A12TR u2940 ( .A(rstkram[145]), .B(rstkram[105]), .C(rstkram[125]), 
        .D(rstkram[85]), .S0(n215), .S1(n214), .Y(n2903) );
  MXIT4_X1M_A12TR u2941 ( .A(rstkram[465]), .B(rstkram[425]), .C(rstkram[445]), 
        .D(rstkram[405]), .S0(n215), .S1(n214), .Y(n2908) );
  MXIT4_X1M_A12TR u2942 ( .A(rstkram[147]), .B(rstkram[107]), .C(rstkram[127]), 
        .D(rstkram[87]), .S0(n215), .S1(n214), .Y(n2923) );
  MXIT4_X1M_A12TR u2943 ( .A(rstkram[467]), .B(rstkram[427]), .C(rstkram[447]), 
        .D(rstkram[407]), .S0(n215), .S1(n214), .Y(n2928) );
  MXIT4_X1M_A12TR u2944 ( .A(rstkram[154]), .B(rstkram[114]), .C(rstkram[134]), 
        .D(rstkram[94]), .S0(n215), .S1(n214), .Y(n2993) );
  MXIT4_X1M_A12TR u2945 ( .A(rstkram[474]), .B(rstkram[434]), .C(rstkram[454]), 
        .D(rstkram[414]), .S0(n215), .S1(n214), .Y(n2998) );
  MXIT4_X1M_A12TR u2946 ( .A(rstkram[143]), .B(rstkram[103]), .C(rstkram[123]), 
        .D(rstkram[83]), .S0(n215), .S1(n214), .Y(n2883) );
  MXIT4_X1M_A12TR u2947 ( .A(rstkram[463]), .B(rstkram[423]), .C(rstkram[443]), 
        .D(rstkram[403]), .S0(n215), .S1(n214), .Y(n2888) );
  MXIT4_X1M_A12TR u2948 ( .A(rstkram[159]), .B(rstkram[119]), .C(rstkram[139]), 
        .D(rstkram[99]), .S0(n215), .S1(n214), .Y(n3043) );
  MXIT4_X1M_A12TR u2949 ( .A(rstkram[479]), .B(rstkram[439]), .C(rstkram[459]), 
        .D(rstkram[419]), .S0(n215), .S1(n214), .Y(n3048) );
  MXIT4_X1M_A12TR u2950 ( .A(rstkram[142]), .B(rstkram[102]), .C(rstkram[122]), 
        .D(rstkram[82]), .S0(n215), .S1(n214), .Y(n2873) );
  MXIT4_X1M_A12TR u2951 ( .A(rstkram[462]), .B(rstkram[422]), .C(rstkram[442]), 
        .D(rstkram[402]), .S0(n215), .S1(n214), .Y(n2878) );
  MXIT4_X1M_A12TR u2952 ( .A(rstkram[300]), .B(rstkram[260]), .C(rstkram[280]), 
        .D(rstkram[240]), .S0(n215), .S1(n214), .Y(n2852) );
  MXIT4_X1M_A12TR u2953 ( .A(rstkram[620]), .B(rstkram[580]), .C(rstkram[600]), 
        .D(rstkram[560]), .S0(n215), .S1(n214), .Y(n2857) );
  MXIT4_X1M_A12TR u2954 ( .A(rstkram[316]), .B(rstkram[276]), .C(rstkram[296]), 
        .D(rstkram[256]), .S0(n215), .S1(n214), .Y(n3012) );
  MXIT4_X1M_A12TR u2955 ( .A(rstkram[636]), .B(rstkram[596]), .C(rstkram[616]), 
        .D(rstkram[576]), .S0(n215), .S1(n214), .Y(n3017) );
  MXIT4_X1M_A12TR u2956 ( .A(rstkram[315]), .B(rstkram[275]), .C(rstkram[295]), 
        .D(rstkram[255]), .S0(n215), .S1(n214), .Y(n3002) );
  MXIT4_X1M_A12TR u2957 ( .A(rstkram[635]), .B(rstkram[595]), .C(rstkram[615]), 
        .D(rstkram[575]), .S0(n215), .S1(n214), .Y(n3007) );
  MXIT4_X1M_A12TR u2958 ( .A(rstkram[306]), .B(rstkram[266]), .C(rstkram[286]), 
        .D(rstkram[246]), .S0(n215), .S1(n214), .Y(n2912) );
  MXIT4_X1M_A12TR u2959 ( .A(rstkram[626]), .B(rstkram[586]), .C(rstkram[606]), 
        .D(rstkram[566]), .S0(n215), .S1(n214), .Y(n2917) );
  MXIT4_X1M_A12TR u2960 ( .A(rstkram[308]), .B(rstkram[268]), .C(rstkram[288]), 
        .D(rstkram[248]), .S0(n215), .S1(n214), .Y(n2932) );
  MXIT4_X1M_A12TR u2961 ( .A(rstkram[628]), .B(rstkram[588]), .C(rstkram[608]), 
        .D(rstkram[568]), .S0(n215), .S1(n214), .Y(n2937) );
  MXIT4_X1M_A12TR u2962 ( .A(rstkram[309]), .B(rstkram[269]), .C(rstkram[289]), 
        .D(rstkram[249]), .S0(n215), .S1(n214), .Y(n2942) );
  MXIT4_X1M_A12TR u2963 ( .A(rstkram[629]), .B(rstkram[589]), .C(rstkram[609]), 
        .D(rstkram[569]), .S0(n215), .S1(n214), .Y(n2947) );
  MXIT4_X1M_A12TR u2964 ( .A(rstkram[310]), .B(rstkram[270]), .C(rstkram[290]), 
        .D(rstkram[250]), .S0(n215), .S1(n214), .Y(n2952) );
  MXIT4_X1M_A12TR u2965 ( .A(rstkram[630]), .B(rstkram[590]), .C(rstkram[610]), 
        .D(rstkram[570]), .S0(n215), .S1(n214), .Y(n2957) );
  MXIT4_X1M_A12TR u2966 ( .A(rstkram[311]), .B(rstkram[271]), .C(rstkram[291]), 
        .D(rstkram[251]), .S0(n215), .S1(n214), .Y(n2962) );
  MXIT4_X1M_A12TR u2967 ( .A(rstkram[631]), .B(rstkram[591]), .C(rstkram[611]), 
        .D(rstkram[571]), .S0(n215), .S1(n214), .Y(n2967) );
  MXIT4_X1M_A12TR u2968 ( .A(rstkram[312]), .B(rstkram[272]), .C(rstkram[292]), 
        .D(rstkram[252]), .S0(n215), .S1(n214), .Y(n2972) );
  MXIT4_X1M_A12TR u2969 ( .A(rstkram[632]), .B(rstkram[592]), .C(rstkram[612]), 
        .D(rstkram[572]), .S0(n215), .S1(n214), .Y(n2977) );
  MXIT4_X1M_A12TR u2970 ( .A(rstkram[313]), .B(rstkram[273]), .C(rstkram[293]), 
        .D(rstkram[253]), .S0(n215), .S1(n214), .Y(n2982) );
  MXIT4_X1M_A12TR u2971 ( .A(rstkram[633]), .B(rstkram[593]), .C(rstkram[613]), 
        .D(rstkram[573]), .S0(n215), .S1(n214), .Y(n2987) );
  MXIT4_X1M_A12TR u2972 ( .A(rstkram[301]), .B(rstkram[261]), .C(rstkram[281]), 
        .D(rstkram[241]), .S0(n215), .S1(n214), .Y(n2862) );
  MXIT4_X1M_A12TR u2973 ( .A(rstkram[621]), .B(rstkram[581]), .C(rstkram[601]), 
        .D(rstkram[561]), .S0(n215), .S1(n214), .Y(n2867) );
  MXIT4_X1M_A12TR u2974 ( .A(rstkram[307]), .B(rstkram[267]), .C(rstkram[287]), 
        .D(rstkram[247]), .S0(n215), .S1(n214), .Y(n2922) );
  MXIT4_X1M_A12TR u2975 ( .A(rstkram[627]), .B(rstkram[587]), .C(rstkram[607]), 
        .D(rstkram[567]), .S0(n215), .S1(n214), .Y(n2927) );
  MXIT4_X1M_A12TR u2976 ( .A(rstkram[314]), .B(rstkram[274]), .C(rstkram[294]), 
        .D(rstkram[254]), .S0(n215), .S1(n214), .Y(n2992) );
  MXIT4_X1M_A12TR u2977 ( .A(rstkram[634]), .B(rstkram[594]), .C(rstkram[614]), 
        .D(rstkram[574]), .S0(n215), .S1(n214), .Y(n2997) );
  MXIT4_X1M_A12TR u2978 ( .A(rstkram[303]), .B(rstkram[263]), .C(rstkram[283]), 
        .D(rstkram[243]), .S0(n215), .S1(n214), .Y(n2882) );
  MXIT4_X1M_A12TR u2979 ( .A(rstkram[623]), .B(rstkram[583]), .C(rstkram[603]), 
        .D(rstkram[563]), .S0(n215), .S1(n214), .Y(n2887) );
  MXIT4_X1M_A12TR u2980 ( .A(rstkram[302]), .B(rstkram[262]), .C(rstkram[282]), 
        .D(rstkram[242]), .S0(n215), .S1(n214), .Y(n2872) );
  MXIT4_X1M_A12TR u2981 ( .A(rstkram[622]), .B(rstkram[582]), .C(rstkram[602]), 
        .D(rstkram[562]), .S0(n215), .S1(n214), .Y(n2877) );
  MXIT4_X1M_A12TR u2982 ( .A(rstkram[220]), .B(rstkram[180]), .C(rstkram[200]), 
        .D(rstkram[160]), .S0(n215), .S1(n214), .Y(n2854) );
  MXIT4_X1M_A12TR u2983 ( .A(rstkram[540]), .B(rstkram[500]), .C(rstkram[520]), 
        .D(rstkram[480]), .S0(n215), .S1(n214), .Y(n2859) );
  MXIT4_X1M_A12TR u2984 ( .A(rstkram[236]), .B(rstkram[196]), .C(rstkram[216]), 
        .D(rstkram[176]), .S0(n215), .S1(n214), .Y(n3014) );
  MXIT4_X1M_A12TR u2985 ( .A(rstkram[556]), .B(rstkram[516]), .C(rstkram[536]), 
        .D(rstkram[496]), .S0(n215), .S1(n214), .Y(n3019) );
  MXIT4_X1M_A12TR u2986 ( .A(rstkram[235]), .B(rstkram[195]), .C(rstkram[215]), 
        .D(rstkram[175]), .S0(n215), .S1(n214), .Y(n3004) );
  MXIT4_X1M_A12TR u2987 ( .A(rstkram[555]), .B(rstkram[515]), .C(rstkram[535]), 
        .D(rstkram[495]), .S0(n215), .S1(n214), .Y(n3009) );
  MXIT4_X1M_A12TR u2988 ( .A(rstkram[226]), .B(rstkram[186]), .C(rstkram[206]), 
        .D(rstkram[166]), .S0(n215), .S1(n214), .Y(n2914) );
  MXIT4_X1M_A12TR u2989 ( .A(rstkram[546]), .B(rstkram[506]), .C(rstkram[526]), 
        .D(rstkram[486]), .S0(n215), .S1(n214), .Y(n2919) );
  MXIT4_X1M_A12TR u2990 ( .A(rstkram[228]), .B(rstkram[188]), .C(rstkram[208]), 
        .D(rstkram[168]), .S0(n215), .S1(n214), .Y(n2934) );
  MXIT4_X1M_A12TR u2991 ( .A(rstkram[548]), .B(rstkram[508]), .C(rstkram[528]), 
        .D(rstkram[488]), .S0(n215), .S1(n214), .Y(n2939) );
  MXIT4_X1M_A12TR u2992 ( .A(rstkram[229]), .B(rstkram[189]), .C(rstkram[209]), 
        .D(rstkram[169]), .S0(n215), .S1(n214), .Y(n2944) );
  MXIT4_X1M_A12TR u2993 ( .A(rstkram[549]), .B(rstkram[509]), .C(rstkram[529]), 
        .D(rstkram[489]), .S0(n215), .S1(n214), .Y(n2949) );
  MXIT4_X1M_A12TR u2994 ( .A(rstkram[230]), .B(rstkram[190]), .C(rstkram[210]), 
        .D(rstkram[170]), .S0(n215), .S1(n214), .Y(n2954) );
  MXIT4_X1M_A12TR u2995 ( .A(rstkram[550]), .B(rstkram[510]), .C(rstkram[530]), 
        .D(rstkram[490]), .S0(n215), .S1(n214), .Y(n2959) );
  MXIT4_X1M_A12TR u2996 ( .A(rstkram[231]), .B(rstkram[191]), .C(rstkram[211]), 
        .D(rstkram[171]), .S0(n215), .S1(n214), .Y(n2964) );
  MXIT4_X1M_A12TR u2997 ( .A(rstkram[551]), .B(rstkram[511]), .C(rstkram[531]), 
        .D(rstkram[491]), .S0(n215), .S1(n214), .Y(n2969) );
  MXIT4_X1M_A12TR u2998 ( .A(rstkram[232]), .B(rstkram[192]), .C(rstkram[212]), 
        .D(rstkram[172]), .S0(n215), .S1(n214), .Y(n2974) );
  MXIT4_X1M_A12TR u2999 ( .A(rstkram[552]), .B(rstkram[512]), .C(rstkram[532]), 
        .D(rstkram[492]), .S0(n215), .S1(n214), .Y(n2979) );
  MXIT4_X1M_A12TR u3000 ( .A(rstkram[233]), .B(rstkram[193]), .C(rstkram[213]), 
        .D(rstkram[173]), .S0(n215), .S1(n214), .Y(n2984) );
  MXIT4_X1M_A12TR u3001 ( .A(rstkram[553]), .B(rstkram[513]), .C(rstkram[533]), 
        .D(rstkram[493]), .S0(n215), .S1(n214), .Y(n2989) );
  MXIT4_X1M_A12TR u3002 ( .A(rstkram[221]), .B(rstkram[181]), .C(rstkram[201]), 
        .D(rstkram[161]), .S0(n215), .S1(n214), .Y(n2864) );
  MXIT4_X1M_A12TR u3003 ( .A(rstkram[541]), .B(rstkram[501]), .C(rstkram[521]), 
        .D(rstkram[481]), .S0(n215), .S1(n214), .Y(n2869) );
  MXIT4_X1M_A12TR u3004 ( .A(rstkram[227]), .B(rstkram[187]), .C(rstkram[207]), 
        .D(rstkram[167]), .S0(n215), .S1(n214), .Y(n2924) );
  MXIT4_X1M_A12TR u3005 ( .A(rstkram[547]), .B(rstkram[507]), .C(rstkram[527]), 
        .D(rstkram[487]), .S0(n215), .S1(n214), .Y(n2929) );
  MXIT4_X1M_A12TR u3006 ( .A(rstkram[234]), .B(rstkram[194]), .C(rstkram[214]), 
        .D(rstkram[174]), .S0(n215), .S1(n214), .Y(n2994) );
  MXIT4_X1M_A12TR u3007 ( .A(rstkram[554]), .B(rstkram[514]), .C(rstkram[534]), 
        .D(rstkram[494]), .S0(n215), .S1(n214), .Y(n2999) );
  MXIT4_X1M_A12TR u3008 ( .A(rstkram[223]), .B(rstkram[183]), .C(rstkram[203]), 
        .D(rstkram[163]), .S0(n215), .S1(n214), .Y(n2884) );
  MXIT4_X1M_A12TR u3009 ( .A(rstkram[543]), .B(rstkram[503]), .C(rstkram[523]), 
        .D(rstkram[483]), .S0(n215), .S1(n214), .Y(n2889) );
  MXIT4_X1M_A12TR u3010 ( .A(rstkram[222]), .B(rstkram[182]), .C(rstkram[202]), 
        .D(rstkram[162]), .S0(n215), .S1(n214), .Y(n2874) );
  MXIT4_X1M_A12TR u3011 ( .A(rstkram[542]), .B(rstkram[502]), .C(rstkram[522]), 
        .D(rstkram[482]), .S0(n215), .S1(n214), .Y(n2879) );
  MXIT4_X1M_A12TR u3012 ( .A(rstkram[60]), .B(rstkram[20]), .C(rstkram[40]), 
        .D(rstkram[0]), .S0(n215), .S1(n214), .Y(n2855) );
  MXIT4_X1M_A12TR u3013 ( .A(rstkram[76]), .B(rstkram[36]), .C(rstkram[56]), 
        .D(rstkram[16]), .S0(n215), .S1(n214), .Y(n3015) );
  MXIT4_X1M_A12TR u3014 ( .A(rstkram[75]), .B(rstkram[35]), .C(rstkram[55]), 
        .D(rstkram[15]), .S0(n215), .S1(n214), .Y(n3005) );
  MXIT4_X1M_A12TR u3015 ( .A(rstkram[66]), .B(rstkram[26]), .C(rstkram[46]), 
        .D(rstkram[6]), .S0(n215), .S1(n214), .Y(n2915) );
  MXIT4_X1M_A12TR u3016 ( .A(rstkram[68]), .B(rstkram[28]), .C(rstkram[48]), 
        .D(rstkram[8]), .S0(n215), .S1(n214), .Y(n2935) );
  MXIT4_X1M_A12TR u3017 ( .A(rstkram[69]), .B(rstkram[29]), .C(rstkram[49]), 
        .D(rstkram[9]), .S0(n215), .S1(n214), .Y(n2945) );
  MXIT4_X1M_A12TR u3018 ( .A(rstkram[70]), .B(rstkram[30]), .C(rstkram[50]), 
        .D(rstkram[10]), .S0(n215), .S1(n214), .Y(n2955) );
  MXIT4_X1M_A12TR u3019 ( .A(rstkram[71]), .B(rstkram[31]), .C(rstkram[51]), 
        .D(rstkram[11]), .S0(n215), .S1(n214), .Y(n2965) );
  MXIT4_X1M_A12TR u3020 ( .A(rstkram[72]), .B(rstkram[32]), .C(rstkram[52]), 
        .D(rstkram[12]), .S0(n215), .S1(n214), .Y(n2975) );
  MXIT4_X1M_A12TR u3021 ( .A(rstkram[73]), .B(rstkram[33]), .C(rstkram[53]), 
        .D(rstkram[13]), .S0(n215), .S1(n214), .Y(n2985) );
  MXIT4_X1M_A12TR u3022 ( .A(rstkram[61]), .B(rstkram[21]), .C(rstkram[41]), 
        .D(rstkram[1]), .S0(n215), .S1(n214), .Y(n2865) );
  MXIT4_X1M_A12TR u3023 ( .A(rstkram[67]), .B(rstkram[27]), .C(rstkram[47]), 
        .D(rstkram[7]), .S0(n215), .S1(n214), .Y(n2925) );
  MXIT4_X1M_A12TR u3024 ( .A(rstkram[74]), .B(rstkram[34]), .C(rstkram[54]), 
        .D(rstkram[14]), .S0(n215), .S1(n214), .Y(n2995) );
  MXIT4_X1M_A12TR u3025 ( .A(rstkram[63]), .B(rstkram[23]), .C(rstkram[43]), 
        .D(rstkram[3]), .S0(n215), .S1(n214), .Y(n2885) );
  MXIT4_X1M_A12TR u3026 ( .A(rstkram[62]), .B(rstkram[22]), .C(rstkram[42]), 
        .D(rstkram[2]), .S0(n215), .S1(n214), .Y(n2875) );
  NOR2_X1M_A12TR u3027 ( .A(n2787), .B(n218), .Y(n2848) );
  AND2_X1M_A12TR u3028 ( .A(rireg[0]), .B(iwb_adr_o[1]), .Y(n2786) );
  OR2_X1M_A12TR u3029 ( .A(n2788), .B(n217), .Y(n2787) );
  OR2_X1M_A12TR u3030 ( .A(n2785), .B(n216), .Y(n2788) );
  MXIT4_X1M_A12TR u3031 ( .A(n3032), .B(n3033), .C(n3034), .D(n3035), .S0(n217), .S1(n216), .Y(n3031) );
  MXIT4_X1M_A12TR u3032 ( .A(rstkram[78]), .B(rstkram[38]), .C(rstkram[58]), 
        .D(rstkram[18]), .S0(n215), .S1(n214), .Y(n3035) );
  MXIT4_X1M_A12TR u3033 ( .A(rstkram[238]), .B(rstkram[198]), .C(rstkram[218]), 
        .D(rstkram[178]), .S0(n215), .S1(n214), .Y(n3034) );
  MXIT4_X1M_A12TR u3034 ( .A(rstkram[318]), .B(rstkram[278]), .C(rstkram[298]), 
        .D(rstkram[258]), .S0(n215), .S1(n214), .Y(n3032) );
  MXIT4_X1M_A12TR u3035 ( .A(n3022), .B(n3023), .C(n3024), .D(n3025), .S0(n217), .S1(n216), .Y(n3021) );
  MXIT4_X1M_A12TR u3036 ( .A(rstkram[77]), .B(rstkram[37]), .C(rstkram[57]), 
        .D(rstkram[17]), .S0(n215), .S1(n214), .Y(n3025) );
  MXIT4_X1M_A12TR u3037 ( .A(rstkram[237]), .B(rstkram[197]), .C(rstkram[217]), 
        .D(rstkram[177]), .S0(n215), .S1(n214), .Y(n3024) );
  MXIT4_X1M_A12TR u3038 ( .A(rstkram[317]), .B(rstkram[277]), .C(rstkram[297]), 
        .D(rstkram[257]), .S0(n215), .S1(n214), .Y(n3022) );
  MXIT4_X1M_A12TR u3039 ( .A(n2892), .B(n2893), .C(n2894), .D(n2895), .S0(n217), .S1(n216), .Y(n2891) );
  MXIT4_X1M_A12TR u3040 ( .A(rstkram[64]), .B(rstkram[24]), .C(rstkram[44]), 
        .D(rstkram[4]), .S0(n215), .S1(n214), .Y(n2895) );
  MXIT4_X1M_A12TR u3041 ( .A(rstkram[224]), .B(rstkram[184]), .C(rstkram[204]), 
        .D(rstkram[164]), .S0(n215), .S1(n214), .Y(n2894) );
  MXIT4_X1M_A12TR u3042 ( .A(rstkram[304]), .B(rstkram[264]), .C(rstkram[284]), 
        .D(rstkram[244]), .S0(n215), .S1(n214), .Y(n2892) );
  MXIT4_X1M_A12TR u3043 ( .A(n2902), .B(n2903), .C(n2904), .D(n2905), .S0(n217), .S1(n216), .Y(n2901) );
  MXIT4_X1M_A12TR u3044 ( .A(rstkram[65]), .B(rstkram[25]), .C(rstkram[45]), 
        .D(rstkram[5]), .S0(n215), .S1(n214), .Y(n2905) );
  MXIT4_X1M_A12TR u3045 ( .A(rstkram[225]), .B(rstkram[185]), .C(rstkram[205]), 
        .D(rstkram[165]), .S0(n215), .S1(n214), .Y(n2904) );
  MXIT4_X1M_A12TR u3046 ( .A(rstkram[305]), .B(rstkram[265]), .C(rstkram[285]), 
        .D(rstkram[245]), .S0(n215), .S1(n214), .Y(n2902) );
  MXIT4_X1M_A12TR u3047 ( .A(n3042), .B(n3043), .C(n3044), .D(n3045), .S0(n217), .S1(n216), .Y(n3041) );
  MXIT4_X1M_A12TR u3048 ( .A(rstkram[79]), .B(rstkram[39]), .C(rstkram[59]), 
        .D(rstkram[19]), .S0(n215), .S1(n214), .Y(n3045) );
  MXIT4_X1M_A12TR u3049 ( .A(rstkram[239]), .B(rstkram[199]), .C(rstkram[219]), 
        .D(rstkram[179]), .S0(n215), .S1(n214), .Y(n3044) );
  MXIT4_X1M_A12TR u3050 ( .A(rstkram[319]), .B(rstkram[279]), .C(rstkram[299]), 
        .D(rstkram[259]), .S0(n215), .S1(n214), .Y(n3042) );
  MXIT4_X1M_A12TR u3051 ( .A(n3037), .B(n3038), .C(n3039), .D(n3040), .S0(n217), .S1(n216), .Y(n3036) );
  MXIT4_X1M_A12TR u3052 ( .A(rstkram[398]), .B(rstkram[358]), .C(rstkram[378]), 
        .D(rstkram[338]), .S0(n215), .S1(n214), .Y(n3040) );
  MXIT4_X1M_A12TR u3053 ( .A(rstkram[558]), .B(rstkram[518]), .C(rstkram[538]), 
        .D(rstkram[498]), .S0(n215), .S1(n214), .Y(n3039) );
  MXIT4_X1M_A12TR u3054 ( .A(rstkram[638]), .B(rstkram[598]), .C(rstkram[618]), 
        .D(rstkram[578]), .S0(n215), .S1(n214), .Y(n3037) );
  MXIT4_X1M_A12TR u3055 ( .A(n3027), .B(n3028), .C(n3029), .D(n3030), .S0(n217), .S1(n216), .Y(n3026) );
  MXIT4_X1M_A12TR u3056 ( .A(rstkram[397]), .B(rstkram[357]), .C(rstkram[377]), 
        .D(rstkram[337]), .S0(n215), .S1(n214), .Y(n3030) );
  MXIT4_X1M_A12TR u3057 ( .A(rstkram[557]), .B(rstkram[517]), .C(rstkram[537]), 
        .D(rstkram[497]), .S0(n215), .S1(n214), .Y(n3029) );
  MXIT4_X1M_A12TR u3058 ( .A(rstkram[637]), .B(rstkram[597]), .C(rstkram[617]), 
        .D(rstkram[577]), .S0(n215), .S1(n214), .Y(n3027) );
  MXIT4_X1M_A12TR u3059 ( .A(n2897), .B(n2898), .C(n2899), .D(n2900), .S0(n217), .S1(n216), .Y(n2896) );
  MXIT4_X1M_A12TR u3060 ( .A(rstkram[384]), .B(rstkram[344]), .C(rstkram[364]), 
        .D(rstkram[324]), .S0(n215), .S1(n214), .Y(n2900) );
  MXIT4_X1M_A12TR u3061 ( .A(rstkram[544]), .B(rstkram[504]), .C(rstkram[524]), 
        .D(rstkram[484]), .S0(n215), .S1(n214), .Y(n2899) );
  MXIT4_X1M_A12TR u3062 ( .A(rstkram[624]), .B(rstkram[584]), .C(rstkram[604]), 
        .D(rstkram[564]), .S0(n215), .S1(n214), .Y(n2897) );
  MXIT4_X1M_A12TR u3063 ( .A(n2907), .B(n2908), .C(n2909), .D(n2910), .S0(n217), .S1(n216), .Y(n2906) );
  MXIT4_X1M_A12TR u3064 ( .A(rstkram[385]), .B(rstkram[345]), .C(rstkram[365]), 
        .D(rstkram[325]), .S0(n215), .S1(n214), .Y(n2910) );
  MXIT4_X1M_A12TR u3065 ( .A(rstkram[545]), .B(rstkram[505]), .C(rstkram[525]), 
        .D(rstkram[485]), .S0(n215), .S1(n214), .Y(n2909) );
  MXIT4_X1M_A12TR u3066 ( .A(rstkram[625]), .B(rstkram[585]), .C(rstkram[605]), 
        .D(rstkram[565]), .S0(n215), .S1(n214), .Y(n2907) );
  MXIT4_X1M_A12TR u3067 ( .A(n3047), .B(n3048), .C(n3049), .D(n3050), .S0(n217), .S1(n216), .Y(n3046) );
  MXIT4_X1M_A12TR u3068 ( .A(rstkram[399]), .B(rstkram[359]), .C(rstkram[379]), 
        .D(rstkram[339]), .S0(n215), .S1(n214), .Y(n3050) );
  MXIT4_X1M_A12TR u3069 ( .A(rstkram[559]), .B(rstkram[519]), .C(rstkram[539]), 
        .D(rstkram[499]), .S0(n215), .S1(n214), .Y(n3049) );
  MXIT4_X1M_A12TR u3070 ( .A(rstkram[639]), .B(rstkram[599]), .C(rstkram[619]), 
        .D(rstkram[579]), .S0(n215), .S1(n214), .Y(n3047) );
  AND2_X1M_A12TR u3071 ( .A(wadd[0]), .B(wrrc_7_), .Y(n2789) );
  OR2_X1M_A12TR u3072 ( .A(wsub[0]), .B(wrrc_7_), .Y(n2790) );
  TIEHI_X1M_A12TR u3073 ( .Y(n3) );
  TIELO_X1M_A12TR u3074 ( .Y(iwb_adr_o[0]) );
  AO21A1AI2_X0P5M_A12TR u3075 ( .A0(n3052), .A1(n3053), .B0(n3054), .C0(n3055), 
        .Y(rnxt[1]) );
  AO21A1AI2_X0P5M_A12TR u3076 ( .A0(rsleep), .A1(n3056), .B0(n3057), .C0(n3058), .Y(n3055) );
  INV_X0P5B_A12TR u3077 ( .A(n3059), .Y(n3057) );
  OAI22_X0P5M_A12TR u3078 ( .A0(n3060), .A1(n3054), .B0(n3061), .B1(n3062), 
        .Y(rnxt[0]) );
  OAI2XB1_X0P5M_A12TR u3079 ( .A1N(n3056), .A0(rsleep), .B0(n3059), .Y(n3062)
         );
  NAND2_X0P5A_A12TR u3080 ( .A(inte_i[7]), .B(n3060), .Y(n3059) );
  NAND2_X0P5A_A12TR u3081 ( .A(inte_i[6]), .B(n3052), .Y(n3056) );
  AND3_X0P5M_A12TR u3082 ( .A(n3063), .B(rintl[0]), .C(rintl[1]), .Y(n3052) );
  INV_X0P5B_A12TR u3083 ( .A(rintl[2]), .Y(n3063) );
  INV_X0P5B_A12TR u3084 ( .A(n3058), .Y(n3061) );
  INV_X0P5B_A12TR u3085 ( .A(n3053), .Y(n3060) );
  NAND3B_X0P5M_A12TR u3086 ( .AN(rinth[2]), .B(rinth[0]), .C(rinth[1]), .Y(
        n3053) );
  INV_X0P5B_A12TR u3087 ( .A(rst_i), .Y(n4431) );
  OAI221_X0P5M_A12TR u3088 ( .A0(n3064), .A1(n3065), .B0(n3066), .B1(n3067), 
        .C0(n3068), .Y(n4432) );
  INV_X0P5B_A12TR u3089 ( .A(wstkw[0]), .Y(n3065) );
  INV_X0P5B_A12TR u3090 ( .A(qrst), .Y(n4433) );
  NAND3B_X0P5M_A12TR u3091 ( .AN(n3070), .B(n3071), .C(n3072), .Y(n4434) );
  MXIT2_X0P5M_A12TR u3092 ( .A(n3073), .B(rmxdst[1]), .S0(n3074), .Y(n3071) );
  OAI22_X0P5M_A12TR u3093 ( .A0(n3075), .A1(n3076), .B0(n3077), .B1(n3078), 
        .Y(n3070) );
  INV_X0P5B_A12TR u3094 ( .A(n3079), .Y(n3077) );
  AOI21_X0P5M_A12TR u3095 ( .A0(n3080), .A1(n3081), .B0(rwdt[16]), .Y(n2745)
         );
  NOR3_X0P5A_A12TR u3096 ( .A(n3082), .B(n3083), .C(n3084), .Y(n3081) );
  NAND3_X0P5A_A12TR u3097 ( .A(n3085), .B(n3086), .C(rromlat[0]), .Y(n3082) );
  NOR3_X0P5A_A12TR u3098 ( .A(n3087), .B(n3088), .C(n3089), .Y(n3080) );
  NAND3_X0P5A_A12TR u3099 ( .A(rromlat[4]), .B(rromlat[3]), .C(rromlat[5]), 
        .Y(n3087) );
  MXIT2_X0P5M_A12TR u3100 ( .A(n3090), .B(n3091), .S0(n3092), .Y(n2744) );
  INV_X0P5B_A12TR u3101 ( .A(rsfrdat[7]), .Y(n3091) );
  NOR3_X0P5A_A12TR u3102 ( .A(n3093), .B(n3094), .C(n3095), .Y(n3090) );
  OAI221_X0P5M_A12TR u3103 ( .A0(n3096), .A1(n3097), .B0(n3098), .B1(n3099), 
        .C0(n3100), .Y(n3095) );
  AOI222_X0P5M_A12TR u3104 ( .A0(wpclat[6]), .A1(n3101), .B0(wstkw[15]), .B1(
        n3102), .C0(rpclatu[7]), .C1(n3103), .Y(n3100) );
  OAI211_X0P5M_A12TR u3105 ( .A0(n3104), .A1(n3105), .B0(n3106), .C0(n3107), 
        .Y(n3094) );
  AOI222_X0P5M_A12TR u3106 ( .A0(rpclath[7]), .A1(n3108), .B0(iwb_dat_o[15]), 
        .B1(n3109), .C0(wstkw[7]), .C1(n3110), .Y(n3107) );
  AOI22_X0P5M_A12TR u3107 ( .A0(wfilebsr[15]), .A1(n3111), .B0(rwreg[7]), .B1(
        n3112), .Y(n3106) );
  NAND4_X0P5A_A12TR u3108 ( .A(n3113), .B(n3114), .C(n3115), .D(n3116), .Y(
        n3093) );
  AOI222_X0P5M_A12TR u3109 ( .A0(rfsr1h[7]), .A1(n3117), .B0(wtblat[15]), .B1(
        n3118), .C0(wtblat[7]), .C1(n3119), .Y(n3116) );
  AOI222_X0P5M_A12TR u3110 ( .A0(rprodh[7]), .A1(n3120), .B0(rfsr1l[7]), .B1(
        n3121), .C0(rfsr2l[7]), .C1(n3122), .Y(n3115) );
  AOI222_X0P5M_A12TR u3111 ( .A0(rfsr0l[7]), .A1(n3123), .B0(n3124), .B1(n3125), .C0(rprng[7]), .C1(n3126), .Y(n3114) );
  AOI22_X0P5M_A12TR u3112 ( .A0(rfsr0h[7]), .A1(n3127), .B0(rprodl[7]), .B1(
        n3128), .Y(n3113) );
  OAI22_X0P5M_A12TR u3113 ( .A0(n3129), .A1(n3130), .B0(n3131), .B1(n3132), 
        .Y(n2743) );
  AOI222_X0P5M_A12TR u3114 ( .A0(rstatus_[3]), .A1(n3133), .B0(n3134), .B1(
        n3135), .C0(dwb_dat_o[3]), .C1(n3136), .Y(n3132) );
  XNOR2_X0P5M_A12TR u3115 ( .A(rsrc[7]), .B(rtgt[7]), .Y(n3135) );
  NOR2_X0P5A_A12TR u3116 ( .A(n3137), .B(n3138), .Y(n3134) );
  XNOR2_X0P5M_A12TR u3117 ( .A(rsrc[7]), .B(dwb_dat_o[7]), .Y(n3137) );
  INV_X0P5B_A12TR u3118 ( .A(rov), .Y(n3130) );
  AO21A1AI2_X0P5M_A12TR u3119 ( .A0(n3139), .A1(n3140), .B0(n3141), .C0(n3142), 
        .Y(n2742) );
  AO21A1AI2_X0P5M_A12TR u3120 ( .A0(n3143), .A1(dwb_dat_o[7]), .B0(n3144), 
        .C0(n3139), .Y(n3142) );
  OAI22_X0P5M_A12TR u3121 ( .A0(n3145), .A1(n3146), .B0(n3147), .B1(n3148), 
        .Y(n3144) );
  AND2_X0P5M_A12TR u3122 ( .A(n3149), .B(n3150), .Y(n3139) );
  NAND4_X0P5A_A12TR u3123 ( .A(rmxstal[0]), .B(rmxstal[1]), .C(n3151), .D(
        n3152), .Y(n3150) );
  AO21A1AI2_X0P5M_A12TR u3124 ( .A0(n3140), .A1(n3149), .B0(n3153), .C0(n3154), 
        .Y(n2741) );
  AO21A1AI2_X0P5M_A12TR u3125 ( .A0(n3155), .A1(n3143), .B0(n3156), .C0(n3149), 
        .Y(n3154) );
  OAI22_X0P5M_A12TR u3126 ( .A0(n3145), .A1(n3157), .B0(n3147), .B1(n3158), 
        .Y(n3156) );
  AO21A1AI2_X0P5M_A12TR u3127 ( .A0(n3159), .A1(n3160), .B0(n3161), .C0(n3151), 
        .Y(n3149) );
  MXIT2_X0P5M_A12TR u3128 ( .A(n3162), .B(n3163), .S0(n3092), .Y(n2740) );
  INV_X0P5B_A12TR u3129 ( .A(rsfrdat[4]), .Y(n3163) );
  NOR3_X0P5A_A12TR u3130 ( .A(n3164), .B(n3165), .C(n3166), .Y(n3162) );
  OAI221_X0P5M_A12TR u3131 ( .A0(n3096), .A1(n3167), .B0(n3098), .B1(n3168), 
        .C0(n3169), .Y(n3166) );
  AOI222_X0P5M_A12TR u3132 ( .A0(wpclat[3]), .A1(n3101), .B0(wstkw[12]), .B1(
        n3102), .C0(rpclatu[4]), .C1(n3103), .Y(n3169) );
  INV_X0P5B_A12TR u3133 ( .A(n218), .Y(n3168) );
  OAI211_X0P5M_A12TR u3134 ( .A0(n3104), .A1(n3170), .B0(n3171), .C0(n3172), 
        .Y(n3165) );
  AOI222_X0P5M_A12TR u3135 ( .A0(rpclath[4]), .A1(n3108), .B0(iwb_dat_o[12]), 
        .B1(n3109), .C0(wstkw[4]), .C1(n3110), .Y(n3172) );
  AOI22_X0P5M_A12TR u3136 ( .A0(wfilebsr[12]), .A1(n3111), .B0(rwreg[4]), .B1(
        n3112), .Y(n3171) );
  NAND4_X0P5A_A12TR u3137 ( .A(n3173), .B(n3174), .C(n3175), .D(n3176), .Y(
        n3164) );
  AOI222_X0P5M_A12TR u3138 ( .A0(wtblat[4]), .A1(n3119), .B0(rn), .B1(n3177), 
        .C0(wtblat[12]), .C1(n3118), .Y(n3176) );
  AOI222_X0P5M_A12TR u3139 ( .A0(rfsr2l[4]), .A1(n3122), .B0(rfsr1h[4]), .B1(
        n3117), .C0(rfsr1l[4]), .C1(n3121), .Y(n3175) );
  AOI222_X0P5M_A12TR u3140 ( .A0(rprng[4]), .A1(n3126), .B0(rprodh[4]), .B1(
        n3120), .C0(rfsr2h[4]), .C1(n3124), .Y(n3174) );
  AOI222_X0P5M_A12TR u3141 ( .A0(rprodl[4]), .A1(n3128), .B0(rfsr0l[4]), .B1(
        n3123), .C0(rfsr0h[4]), .C1(n3127), .Y(n3173) );
  AO21A1AI2_X0P5M_A12TR u3142 ( .A0(n3140), .A1(n3178), .B0(n3179), .C0(n3180), 
        .Y(n2739) );
  AO21A1AI2_X0P5M_A12TR u3143 ( .A0(rc_), .A1(n3143), .B0(n3181), .C0(n3178), 
        .Y(n3180) );
  OAI22_X0P5M_A12TR u3144 ( .A0(n3145), .A1(n3182), .B0(n3067), .B1(n3147), 
        .Y(n3181) );
  INV_X0P5B_A12TR u3145 ( .A(n3133), .Y(n3145) );
  OAI21_X0P5M_A12TR u3146 ( .A0(rmxstal[1]), .A1(n3161), .B0(n3131), .Y(n3178)
         );
  OAI221_X0P5M_A12TR u3147 ( .A0(n3089), .A1(n3183), .B0(n3184), .B1(n3185), 
        .C0(n3186), .Y(n2738) );
  AOI222_X0P5M_A12TR u3148 ( .A0(wfsrdec2[7]), .A1(n3187), .B0(rfsr2l[7]), 
        .B1(n3188), .C0(n3189), .C1(dwb_dat_o[7]), .Y(n3186) );
  INV_X0P5B_A12TR u3149 ( .A(wfsrinc2[7]), .Y(n3185) );
  AO22_X0P5M_A12TR u3150 ( .A0(n240), .A1(n3190), .B0(rwdt[16]), .B1(n3191), 
        .Y(n2737) );
  MXIT2_X0P5M_A12TR u3151 ( .A(n3192), .B(n3193), .S0(n3194), .Y(n2736) );
  MXIT2_X0P5M_A12TR u3152 ( .A(n3083), .B(n3195), .S0(n3194), .Y(n2735) );
  MXIT2_X0P5M_A12TR u3153 ( .A(n3084), .B(n3196), .S0(n3194), .Y(n2734) );
  MXIT2_X0P5M_A12TR u3154 ( .A(n3197), .B(n3198), .S0(n3194), .Y(n2733) );
  MXIT2_X0P5M_A12TR u3155 ( .A(n3199), .B(n3200), .S0(n3194), .Y(n2732) );
  MXIT2_X0P5M_A12TR u3156 ( .A(n3201), .B(n3202), .S0(n3194), .Y(n2731) );
  MXIT2_X0P5M_A12TR u3157 ( .A(n3088), .B(n3203), .S0(n3194), .Y(n2730) );
  MXIT2_X0P5M_A12TR u3158 ( .A(n3089), .B(n3204), .S0(n3194), .Y(n2729) );
  MXIT2_X0P5M_A12TR u3159 ( .A(n3205), .B(n3206), .S0(n3194), .Y(n2728) );
  MXIT2_X0P5M_A12TR u3160 ( .A(n3207), .B(n3208), .S0(n3194), .Y(n2727) );
  MXIT2_X0P5M_A12TR u3161 ( .A(n3209), .B(n3210), .S0(n3194), .Y(n2726) );
  MXIT2_X0P5M_A12TR u3162 ( .A(n3211), .B(n3212), .S0(n3194), .Y(n2725) );
  MXIT2_X0P5M_A12TR u3163 ( .A(n3213), .B(n3214), .S0(n3194), .Y(n2724) );
  MXIT2_X0P5M_A12TR u3164 ( .A(n3215), .B(n3216), .S0(n3194), .Y(n2723) );
  MXIT2_X0P5M_A12TR u3165 ( .A(n3217), .B(n3218), .S0(n3194), .Y(n2722) );
  MXIT2_X0P5M_A12TR u3166 ( .A(n3219), .B(n3220), .S0(n3194), .Y(n2721) );
  NOR2_X0P5A_A12TR u3167 ( .A(n3138), .B(n3221), .Y(n3194) );
  MXIT2_X0P5M_A12TR u3168 ( .A(n3222), .B(n3223), .S0(n3224), .Y(n2720) );
  NAND2_X0P5A_A12TR u3169 ( .A(rintf[1]), .B(n3074), .Y(n3222) );
  MXIT2_X0P5M_A12TR u3170 ( .A(n3225), .B(n3226), .S0(n3224), .Y(n2719) );
  NOR2_X0P5A_A12TR u3171 ( .A(n3058), .B(n3221), .Y(n3224) );
  NOR2_X0P5A_A12TR u3172 ( .A(rfsm[1]), .B(rfsm[0]), .Y(n3058) );
  NAND2_X0P5A_A12TR u3173 ( .A(rintf[0]), .B(n3074), .Y(n3225) );
  MXIT2_X0P5M_A12TR u3174 ( .A(n3192), .B(n3227), .S0(n3228), .Y(n2718) );
  MXIT2_X0P5M_A12TR u3175 ( .A(n3083), .B(n3229), .S0(n3228), .Y(n2717) );
  MXIT2_X0P5M_A12TR u3176 ( .A(n3084), .B(n3230), .S0(n3228), .Y(n2716) );
  MXIT2_X0P5M_A12TR u3177 ( .A(n3197), .B(n3231), .S0(n3228), .Y(n2715) );
  MXIT2_X0P5M_A12TR u3178 ( .A(n3199), .B(n3232), .S0(n3228), .Y(n2714) );
  MXIT2_X0P5M_A12TR u3179 ( .A(n3201), .B(n3233), .S0(n3228), .Y(n2713) );
  MXIT2_X0P5M_A12TR u3180 ( .A(n3088), .B(n3234), .S0(n3228), .Y(n2712) );
  MXIT2_X0P5M_A12TR u3181 ( .A(n3089), .B(n3235), .S0(n3228), .Y(n2711) );
  MXT2_X0P5M_A12TR u3182 ( .A(rromlat[8]), .B(rireg[8]), .S0(n3228), .Y(n2710)
         );
  MXT2_X0P5M_A12TR u3183 ( .A(rromlat[9]), .B(rireg[9]), .S0(n3228), .Y(n2709)
         );
  MXT2_X0P5M_A12TR u3184 ( .A(rromlat[10]), .B(rireg[10]), .S0(n3228), .Y(
        n2708) );
  OAI22_X0P5M_A12TR u3185 ( .A0(n3129), .A1(n3236), .B0(n3131), .B1(n3237), 
        .Y(n2707) );
  AOI222_X0P5M_A12TR u3186 ( .A0(dwb_dat_o[4]), .A1(n3143), .B0(dwb_dat_o[1]), 
        .B1(n3136), .C0(rstatus_[1]), .C1(n3133), .Y(n3237) );
  NOR2_X0P5A_A12TR u3187 ( .A(n3238), .B(n3239), .Y(n3133) );
  INV_X0P5B_A12TR u3188 ( .A(n3147), .Y(n3136) );
  NAND2_X0P5A_A12TR u3189 ( .A(n3177), .B(n3240), .Y(n3147) );
  INV_X0P5B_A12TR u3190 ( .A(rdc), .Y(n3236) );
  NOR2B_X0P5M_A12TR u3191 ( .AN(n3140), .B(n3131), .Y(n3129) );
  INV_X0P5B_A12TR u3192 ( .A(n3241), .Y(n3131) );
  OAI31_X0P5M_A12TR u3193 ( .A0(n3161), .A1(n3160), .A2(n3152), .B0(n3151), 
        .Y(n3241) );
  NAND2_X0P5A_A12TR u3194 ( .A(n3242), .B(n3138), .Y(n3151) );
  INV_X0P5B_A12TR u3195 ( .A(rmxstal[0]), .Y(n3160) );
  NAND2_X0P5A_A12TR u3196 ( .A(n3243), .B(n3242), .Y(n3161) );
  MXIT2_X0P5M_A12TR u3197 ( .A(n3244), .B(n3245), .S0(n3152), .Y(n3243) );
  INV_X0P5B_A12TR u3198 ( .A(rmxstal[2]), .Y(n3152) );
  NOR2_X0P5A_A12TR u3199 ( .A(rmxstal[1]), .B(rmxstal[0]), .Y(n3245) );
  XNOR2_X0P5M_A12TR u3200 ( .A(n3159), .B(rmxstal[0]), .Y(n3244) );
  INV_X0P5B_A12TR u3201 ( .A(rmxstal[1]), .Y(n3159) );
  AOI221_X0P5M_A12TR u3202 ( .A0(n3246), .A1(qfsm[0]), .B0(n3239), .B1(n3247), 
        .C0(n3248), .Y(n3140) );
  MXIT2_X0P5M_A12TR u3203 ( .A(n3249), .B(n3250), .S0(n3092), .Y(n2706) );
  INV_X0P5B_A12TR u3204 ( .A(rsfrdat[0]), .Y(n3250) );
  NOR3_X0P5A_A12TR u3205 ( .A(n3251), .B(n3252), .C(n3253), .Y(n3249) );
  OAI211_X0P5M_A12TR u3206 ( .A0(n3254), .A1(n3255), .B0(n3256), .C0(n3257), 
        .Y(n3253) );
  AOI222_X0P5M_A12TR u3207 ( .A0(rfsr2h[0]), .A1(n3124), .B0(rfsr2l[0]), .B1(
        n3122), .C0(rprodh[0]), .C1(n3120), .Y(n3257) );
  AOI22_X0P5M_A12TR u3208 ( .A0(rprng[0]), .A1(n3126), .B0(rfsr0l[0]), .B1(
        n3123), .Y(n3256) );
  OAI211_X0P5M_A12TR u3209 ( .A0(n3258), .A1(n3259), .B0(n3260), .C0(n3261), 
        .Y(n3252) );
  AOI222_X0P5M_A12TR u3210 ( .A0(rfsr1l[0]), .A1(n3121), .B0(wtblat[0]), .B1(
        n3119), .C0(rfsr1h[0]), .C1(n3117), .Y(n3261) );
  AOI32_X0P5M_A12TR u3211 ( .A0(n3262), .A1(n3263), .A2(rswdten), .B0(wrrc_7_), 
        .B1(n3177), .Y(n3260) );
  NAND4_X0P5A_A12TR u3212 ( .A(n3264), .B(n3265), .C(n3266), .D(n3267), .Y(
        n3251) );
  AOI222_X0P5M_A12TR u3213 ( .A0(rwreg[0]), .A1(n3112), .B0(rprodl[0]), .B1(
        n3128), .C0(wfilebsr[8]), .C1(n3111), .Y(n3267) );
  AOI222_X0P5M_A12TR u3214 ( .A0(n3110), .A1(wstkw[0]), .B0(wtblat[16]), .B1(
        n3268), .C0(iwb_dat_o[8]), .C1(n3109), .Y(n3266) );
  AOI222_X0P5M_A12TR u3215 ( .A0(rpclatu[0]), .A1(n3103), .B0(rpclath[0]), 
        .B1(n3108), .C0(wstkw[8]), .C1(n3102), .Y(n3265) );
  AOI222_X0P5M_A12TR u3216 ( .A0(n214), .A1(n3269), .B0(rpcl_0_), .B1(n3101), 
        .C0(wstkw[16]), .C1(n3270), .Y(n3264) );
  MXIT2_X0P5M_A12TR u3217 ( .A(n3271), .B(n3272), .S0(n3092), .Y(n2705) );
  INV_X0P5B_A12TR u3218 ( .A(rsfrdat[1]), .Y(n3272) );
  NOR3_X0P5A_A12TR u3219 ( .A(n3273), .B(n3274), .C(n3275), .Y(n3271) );
  OAI221_X0P5M_A12TR u3220 ( .A0(n3096), .A1(n3276), .B0(n3098), .B1(n3277), 
        .C0(n3278), .Y(n3275) );
  AOI222_X0P5M_A12TR u3221 ( .A0(wpclat[0]), .A1(n3101), .B0(wstkw[9]), .B1(
        n3102), .C0(rpclatu[1]), .C1(n3103), .Y(n3278) );
  INV_X0P5B_A12TR u3222 ( .A(n215), .Y(n3277) );
  OAI211_X0P5M_A12TR u3223 ( .A0(n3104), .A1(n3279), .B0(n3280), .C0(n3281), 
        .Y(n3274) );
  AOI222_X0P5M_A12TR u3224 ( .A0(rpclath[1]), .A1(n3108), .B0(iwb_dat_o[9]), 
        .B1(n3109), .C0(wstkw[1]), .C1(n3110), .Y(n3281) );
  AOI22_X0P5M_A12TR u3225 ( .A0(wfilebsr[9]), .A1(n3111), .B0(rwreg[1]), .B1(
        n3112), .Y(n3280) );
  NAND4_X0P5A_A12TR u3226 ( .A(n3282), .B(n3283), .C(n3284), .D(n3285), .Y(
        n3273) );
  AOI222_X0P5M_A12TR u3227 ( .A0(wtblat[1]), .A1(n3119), .B0(rdc), .B1(n3177), 
        .C0(wtblat[9]), .C1(n3118), .Y(n3285) );
  AOI222_X0P5M_A12TR u3228 ( .A0(rfsr2l[1]), .A1(n3122), .B0(rfsr1h[1]), .B1(
        n3117), .C0(rfsr1l[1]), .C1(n3121), .Y(n3284) );
  AOI222_X0P5M_A12TR u3229 ( .A0(rprng[1]), .A1(n3126), .B0(rprodh[1]), .B1(
        n3120), .C0(rfsr2h[1]), .C1(n3124), .Y(n3283) );
  AOI222_X0P5M_A12TR u3230 ( .A0(rprodl[1]), .A1(n3128), .B0(rfsr0l[1]), .B1(
        n3123), .C0(rfsr0h[1]), .C1(n3127), .Y(n3282) );
  MXIT2_X0P5M_A12TR u3231 ( .A(n3286), .B(n3287), .S0(n3092), .Y(n2704) );
  INV_X0P5B_A12TR u3232 ( .A(rsfrdat[2]), .Y(n3287) );
  NOR3_X0P5A_A12TR u3233 ( .A(n3288), .B(n3289), .C(n3290), .Y(n3286) );
  OAI221_X0P5M_A12TR u3234 ( .A0(n3096), .A1(n3291), .B0(n3098), .B1(n3292), 
        .C0(n3293), .Y(n3290) );
  AOI222_X0P5M_A12TR u3235 ( .A0(wpclat[1]), .A1(n3101), .B0(wstkw[10]), .B1(
        n3102), .C0(rpclatu[2]), .C1(n3103), .Y(n3293) );
  INV_X0P5B_A12TR u3236 ( .A(n216), .Y(n3292) );
  OAI211_X0P5M_A12TR u3237 ( .A0(n3104), .A1(n3294), .B0(n3295), .C0(n3296), 
        .Y(n3289) );
  AOI222_X0P5M_A12TR u3238 ( .A0(rpclath[2]), .A1(n3108), .B0(iwb_dat_o[10]), 
        .B1(n3109), .C0(wstkw[2]), .C1(n3110), .Y(n3296) );
  AOI22_X0P5M_A12TR u3239 ( .A0(wfilebsr[10]), .A1(n3111), .B0(rwreg[2]), .B1(
        n3112), .Y(n3295) );
  NAND4_X0P5A_A12TR u3240 ( .A(n3297), .B(n3298), .C(n3299), .D(n3300), .Y(
        n3288) );
  AOI222_X0P5M_A12TR u3241 ( .A0(wtblat[2]), .A1(n3119), .B0(rz), .B1(n3177), 
        .C0(wtblat[10]), .C1(n3118), .Y(n3300) );
  AOI222_X0P5M_A12TR u3242 ( .A0(rfsr2l[2]), .A1(n3122), .B0(rfsr1h[2]), .B1(
        n3117), .C0(rfsr1l[2]), .C1(n3121), .Y(n3299) );
  AOI222_X0P5M_A12TR u3243 ( .A0(rprng[2]), .A1(n3126), .B0(rprodh[2]), .B1(
        n3120), .C0(rfsr2h[2]), .C1(n3124), .Y(n3298) );
  AOI222_X0P5M_A12TR u3244 ( .A0(rprodl[2]), .A1(n3128), .B0(rfsr0l[2]), .B1(
        n3123), .C0(rfsr0h[2]), .C1(n3127), .Y(n3297) );
  MXIT2_X0P5M_A12TR u3245 ( .A(n3301), .B(n3302), .S0(n3092), .Y(n2703) );
  INV_X0P5B_A12TR u3246 ( .A(rsfrdat[3]), .Y(n3302) );
  NOR3_X0P5A_A12TR u3247 ( .A(n3303), .B(n3304), .C(n3305), .Y(n3301) );
  OAI221_X0P5M_A12TR u3248 ( .A0(n3096), .A1(n3306), .B0(n3098), .B1(n3307), 
        .C0(n3308), .Y(n3305) );
  AOI222_X0P5M_A12TR u3249 ( .A0(wpclat[2]), .A1(n3101), .B0(wstkw[11]), .B1(
        n3102), .C0(rpclatu[3]), .C1(n3103), .Y(n3308) );
  INV_X0P5B_A12TR u3250 ( .A(n217), .Y(n3307) );
  OAI211_X0P5M_A12TR u3251 ( .A0(n3104), .A1(n3309), .B0(n3310), .C0(n3311), 
        .Y(n3304) );
  AOI222_X0P5M_A12TR u3252 ( .A0(rpclath[3]), .A1(n3108), .B0(iwb_dat_o[11]), 
        .B1(n3109), .C0(wstkw[3]), .C1(n3110), .Y(n3311) );
  AOI22_X0P5M_A12TR u3253 ( .A0(wfilebsr[11]), .A1(n3111), .B0(rwreg[3]), .B1(
        n3112), .Y(n3310) );
  NAND4_X0P5A_A12TR u3254 ( .A(n3312), .B(n3313), .C(n3314), .D(n3315), .Y(
        n3303) );
  AOI222_X0P5M_A12TR u3255 ( .A0(wtblat[3]), .A1(n3119), .B0(rov), .B1(n3177), 
        .C0(wtblat[11]), .C1(n3118), .Y(n3315) );
  INV_X0P5B_A12TR u3256 ( .A(n3246), .Y(n3177) );
  NAND2_X0P5A_A12TR u3257 ( .A(n3316), .B(n3317), .Y(n3246) );
  AOI222_X0P5M_A12TR u3258 ( .A0(rfsr2l[3]), .A1(n3122), .B0(rfsr1h[3]), .B1(
        n3117), .C0(rfsr1l[3]), .C1(n3121), .Y(n3314) );
  AOI222_X0P5M_A12TR u3259 ( .A0(rprng[3]), .A1(n3126), .B0(rprodh[3]), .B1(
        n3120), .C0(rfsr2h[3]), .C1(n3124), .Y(n3313) );
  AOI222_X0P5M_A12TR u3260 ( .A0(rprodl[3]), .A1(n3128), .B0(rfsr0l[3]), .B1(
        n3123), .C0(rfsr0h[3]), .C1(n3127), .Y(n3312) );
  MXIT2_X0P5M_A12TR u3261 ( .A(n3318), .B(n3319), .S0(n3092), .Y(n2702) );
  INV_X0P5B_A12TR u3262 ( .A(rsfrdat[6]), .Y(n3319) );
  NOR3_X0P5A_A12TR u3263 ( .A(n3320), .B(n3321), .C(n3322), .Y(n3318) );
  OAI221_X0P5M_A12TR u3264 ( .A0(n3096), .A1(n3323), .B0(n3098), .B1(n3324), 
        .C0(n3325), .Y(n3322) );
  AOI222_X0P5M_A12TR u3265 ( .A0(wpclat[5]), .A1(n3101), .B0(wstkw[14]), .B1(
        n3102), .C0(rpclatu[6]), .C1(n3103), .Y(n3325) );
  OAI211_X0P5M_A12TR u3266 ( .A0(n3104), .A1(n3326), .B0(n3327), .C0(n3328), 
        .Y(n3321) );
  AOI222_X0P5M_A12TR u3267 ( .A0(rpclath[6]), .A1(n3108), .B0(iwb_dat_o[14]), 
        .B1(n3109), .C0(wstkw[6]), .C1(n3110), .Y(n3328) );
  AOI22_X0P5M_A12TR u3268 ( .A0(wfilebsr[14]), .A1(n3111), .B0(rwreg[6]), .B1(
        n3112), .Y(n3327) );
  NAND4_X0P5A_A12TR u3269 ( .A(n3329), .B(n3330), .C(n3331), .D(n3332), .Y(
        n3320) );
  AOI222_X0P5M_A12TR u3270 ( .A0(rfsr1h[6]), .A1(n3117), .B0(wtblat[14]), .B1(
        n3118), .C0(wtblat[6]), .C1(n3119), .Y(n3332) );
  AOI222_X0P5M_A12TR u3271 ( .A0(rprodh[6]), .A1(n3120), .B0(rfsr1l[6]), .B1(
        n3121), .C0(rfsr2l[6]), .C1(n3122), .Y(n3331) );
  AOI222_X0P5M_A12TR u3272 ( .A0(rfsr0l[6]), .A1(n3123), .B0(n3124), .B1(n3333), .C0(rprng[6]), .C1(n3126), .Y(n3330) );
  AOI22_X0P5M_A12TR u3273 ( .A0(rfsr0h[6]), .A1(n3127), .B0(rprodl[6]), .B1(
        n3128), .Y(n3329) );
  MXT2_X0P5M_A12TR u3274 ( .A(rstkram[636]), .B(wstkw[16]), .S0(n3334), .Y(
        n2701) );
  MXT2_X0P5M_A12TR u3275 ( .A(rstkram[616]), .B(wstkw[16]), .S0(n3335), .Y(
        n2700) );
  MXT2_X0P5M_A12TR u3276 ( .A(rstkram[596]), .B(wstkw[16]), .S0(n3336), .Y(
        n2699) );
  MXT2_X0P5M_A12TR u3277 ( .A(rstkram[576]), .B(wstkw[16]), .S0(n3337), .Y(
        n2698) );
  MXT2_X0P5M_A12TR u3278 ( .A(rstkram[556]), .B(wstkw[16]), .S0(n3338), .Y(
        n2697) );
  MXT2_X0P5M_A12TR u3279 ( .A(rstkram[536]), .B(wstkw[16]), .S0(n3339), .Y(
        n2696) );
  MXT2_X0P5M_A12TR u3280 ( .A(rstkram[516]), .B(wstkw[16]), .S0(n3340), .Y(
        n2695) );
  MXT2_X0P5M_A12TR u3281 ( .A(rstkram[496]), .B(wstkw[16]), .S0(n3341), .Y(
        n2694) );
  MXT2_X0P5M_A12TR u3282 ( .A(rstkram[476]), .B(wstkw[16]), .S0(n3342), .Y(
        n2693) );
  MXT2_X0P5M_A12TR u3283 ( .A(rstkram[456]), .B(wstkw[16]), .S0(n3343), .Y(
        n2692) );
  MXT2_X0P5M_A12TR u3284 ( .A(rstkram[436]), .B(wstkw[16]), .S0(n3344), .Y(
        n2691) );
  MXT2_X0P5M_A12TR u3285 ( .A(rstkram[416]), .B(wstkw[16]), .S0(n3345), .Y(
        n2690) );
  MXT2_X0P5M_A12TR u3286 ( .A(rstkram[396]), .B(wstkw[16]), .S0(n3346), .Y(
        n2689) );
  MXT2_X0P5M_A12TR u3287 ( .A(rstkram[376]), .B(wstkw[16]), .S0(n3347), .Y(
        n2688) );
  MXT2_X0P5M_A12TR u3288 ( .A(rstkram[356]), .B(wstkw[16]), .S0(n3348), .Y(
        n2687) );
  MXT2_X0P5M_A12TR u3289 ( .A(rstkram[336]), .B(wstkw[16]), .S0(n3349), .Y(
        n2686) );
  MXT2_X0P5M_A12TR u3290 ( .A(rstkram[316]), .B(wstkw[16]), .S0(n3350), .Y(
        n2685) );
  MXT2_X0P5M_A12TR u3291 ( .A(rstkram[296]), .B(wstkw[16]), .S0(n3351), .Y(
        n2684) );
  MXT2_X0P5M_A12TR u3292 ( .A(rstkram[276]), .B(wstkw[16]), .S0(n3352), .Y(
        n2683) );
  MXT2_X0P5M_A12TR u3293 ( .A(rstkram[256]), .B(wstkw[16]), .S0(n3353), .Y(
        n2682) );
  MXT2_X0P5M_A12TR u3294 ( .A(rstkram[236]), .B(wstkw[16]), .S0(n3354), .Y(
        n2681) );
  MXT2_X0P5M_A12TR u3295 ( .A(rstkram[216]), .B(wstkw[16]), .S0(n3355), .Y(
        n2680) );
  MXT2_X0P5M_A12TR u3296 ( .A(rstkram[196]), .B(wstkw[16]), .S0(n3356), .Y(
        n2679) );
  MXT2_X0P5M_A12TR u3297 ( .A(rstkram[176]), .B(wstkw[16]), .S0(n3357), .Y(
        n2678) );
  MXT2_X0P5M_A12TR u3298 ( .A(rstkram[156]), .B(wstkw[16]), .S0(n3358), .Y(
        n2677) );
  MXT2_X0P5M_A12TR u3299 ( .A(rstkram[136]), .B(wstkw[16]), .S0(n3359), .Y(
        n2676) );
  MXT2_X0P5M_A12TR u3300 ( .A(rstkram[116]), .B(wstkw[16]), .S0(n3360), .Y(
        n2675) );
  MXT2_X0P5M_A12TR u3301 ( .A(rstkram[96]), .B(wstkw[16]), .S0(n3361), .Y(
        n2674) );
  MXT2_X0P5M_A12TR u3302 ( .A(rstkram[76]), .B(wstkw[16]), .S0(n3362), .Y(
        n2673) );
  MXT2_X0P5M_A12TR u3303 ( .A(rstkram[56]), .B(wstkw[16]), .S0(n3363), .Y(
        n2672) );
  MXT2_X0P5M_A12TR u3304 ( .A(rstkram[36]), .B(wstkw[16]), .S0(n3364), .Y(
        n2671) );
  MXT2_X0P5M_A12TR u3305 ( .A(rstkram[16]), .B(wstkw[16]), .S0(n3365), .Y(
        n2670) );
  MXT2_X0P5M_A12TR u3306 ( .A(rstkram[637]), .B(wstkw[17]), .S0(n3334), .Y(
        n2669) );
  MXT2_X0P5M_A12TR u3307 ( .A(rstkram[617]), .B(wstkw[17]), .S0(n3335), .Y(
        n2668) );
  MXT2_X0P5M_A12TR u3308 ( .A(rstkram[597]), .B(wstkw[17]), .S0(n3336), .Y(
        n2667) );
  MXT2_X0P5M_A12TR u3309 ( .A(rstkram[577]), .B(wstkw[17]), .S0(n3337), .Y(
        n2666) );
  MXT2_X0P5M_A12TR u3310 ( .A(rstkram[557]), .B(wstkw[17]), .S0(n3338), .Y(
        n2665) );
  MXT2_X0P5M_A12TR u3311 ( .A(rstkram[537]), .B(wstkw[17]), .S0(n3339), .Y(
        n2664) );
  MXT2_X0P5M_A12TR u3312 ( .A(rstkram[517]), .B(wstkw[17]), .S0(n3340), .Y(
        n2663) );
  MXT2_X0P5M_A12TR u3313 ( .A(rstkram[497]), .B(wstkw[17]), .S0(n3341), .Y(
        n2662) );
  MXT2_X0P5M_A12TR u3314 ( .A(rstkram[477]), .B(wstkw[17]), .S0(n3342), .Y(
        n2661) );
  MXT2_X0P5M_A12TR u3315 ( .A(rstkram[457]), .B(wstkw[17]), .S0(n3343), .Y(
        n2660) );
  MXT2_X0P5M_A12TR u3316 ( .A(rstkram[437]), .B(wstkw[17]), .S0(n3344), .Y(
        n2659) );
  MXT2_X0P5M_A12TR u3317 ( .A(rstkram[417]), .B(wstkw[17]), .S0(n3345), .Y(
        n2658) );
  MXT2_X0P5M_A12TR u3318 ( .A(rstkram[397]), .B(wstkw[17]), .S0(n3346), .Y(
        n2657) );
  MXT2_X0P5M_A12TR u3319 ( .A(rstkram[377]), .B(wstkw[17]), .S0(n3347), .Y(
        n2656) );
  MXT2_X0P5M_A12TR u3320 ( .A(rstkram[357]), .B(wstkw[17]), .S0(n3348), .Y(
        n2655) );
  MXT2_X0P5M_A12TR u3321 ( .A(rstkram[337]), .B(wstkw[17]), .S0(n3349), .Y(
        n2654) );
  MXT2_X0P5M_A12TR u3322 ( .A(rstkram[317]), .B(wstkw[17]), .S0(n3350), .Y(
        n2653) );
  MXT2_X0P5M_A12TR u3323 ( .A(rstkram[297]), .B(wstkw[17]), .S0(n3351), .Y(
        n2652) );
  MXT2_X0P5M_A12TR u3324 ( .A(rstkram[277]), .B(wstkw[17]), .S0(n3352), .Y(
        n2651) );
  MXT2_X0P5M_A12TR u3325 ( .A(rstkram[257]), .B(wstkw[17]), .S0(n3353), .Y(
        n2650) );
  MXT2_X0P5M_A12TR u3326 ( .A(rstkram[237]), .B(wstkw[17]), .S0(n3354), .Y(
        n2649) );
  MXT2_X0P5M_A12TR u3327 ( .A(rstkram[217]), .B(wstkw[17]), .S0(n3355), .Y(
        n2648) );
  MXT2_X0P5M_A12TR u3328 ( .A(rstkram[197]), .B(wstkw[17]), .S0(n3356), .Y(
        n2647) );
  MXT2_X0P5M_A12TR u3329 ( .A(rstkram[177]), .B(wstkw[17]), .S0(n3357), .Y(
        n2646) );
  MXT2_X0P5M_A12TR u3330 ( .A(rstkram[157]), .B(wstkw[17]), .S0(n3358), .Y(
        n2645) );
  MXT2_X0P5M_A12TR u3331 ( .A(rstkram[137]), .B(wstkw[17]), .S0(n3359), .Y(
        n2644) );
  MXT2_X0P5M_A12TR u3332 ( .A(rstkram[117]), .B(wstkw[17]), .S0(n3360), .Y(
        n2643) );
  MXT2_X0P5M_A12TR u3333 ( .A(rstkram[97]), .B(wstkw[17]), .S0(n3361), .Y(
        n2642) );
  MXT2_X0P5M_A12TR u3334 ( .A(rstkram[77]), .B(wstkw[17]), .S0(n3362), .Y(
        n2641) );
  MXT2_X0P5M_A12TR u3335 ( .A(rstkram[57]), .B(wstkw[17]), .S0(n3363), .Y(
        n2640) );
  MXT2_X0P5M_A12TR u3336 ( .A(rstkram[37]), .B(wstkw[17]), .S0(n3364), .Y(
        n2639) );
  MXT2_X0P5M_A12TR u3337 ( .A(rstkram[17]), .B(wstkw[17]), .S0(n3365), .Y(
        n2638) );
  MXT2_X0P5M_A12TR u3338 ( .A(rstkram[638]), .B(wstkw[18]), .S0(n3334), .Y(
        n2637) );
  MXT2_X0P5M_A12TR u3339 ( .A(rstkram[618]), .B(wstkw[18]), .S0(n3335), .Y(
        n2636) );
  MXT2_X0P5M_A12TR u3340 ( .A(rstkram[598]), .B(wstkw[18]), .S0(n3336), .Y(
        n2635) );
  MXT2_X0P5M_A12TR u3341 ( .A(rstkram[578]), .B(wstkw[18]), .S0(n3337), .Y(
        n2634) );
  MXT2_X0P5M_A12TR u3342 ( .A(rstkram[558]), .B(wstkw[18]), .S0(n3338), .Y(
        n2633) );
  MXT2_X0P5M_A12TR u3343 ( .A(rstkram[538]), .B(wstkw[18]), .S0(n3339), .Y(
        n2632) );
  MXT2_X0P5M_A12TR u3344 ( .A(rstkram[518]), .B(wstkw[18]), .S0(n3340), .Y(
        n2631) );
  MXT2_X0P5M_A12TR u3345 ( .A(rstkram[498]), .B(wstkw[18]), .S0(n3341), .Y(
        n2630) );
  MXT2_X0P5M_A12TR u3346 ( .A(rstkram[478]), .B(wstkw[18]), .S0(n3342), .Y(
        n2629) );
  MXT2_X0P5M_A12TR u3347 ( .A(rstkram[458]), .B(wstkw[18]), .S0(n3343), .Y(
        n2628) );
  MXT2_X0P5M_A12TR u3348 ( .A(rstkram[438]), .B(wstkw[18]), .S0(n3344), .Y(
        n2627) );
  MXT2_X0P5M_A12TR u3349 ( .A(rstkram[418]), .B(wstkw[18]), .S0(n3345), .Y(
        n2626) );
  MXT2_X0P5M_A12TR u3350 ( .A(rstkram[398]), .B(wstkw[18]), .S0(n3346), .Y(
        n2625) );
  MXT2_X0P5M_A12TR u3351 ( .A(rstkram[378]), .B(wstkw[18]), .S0(n3347), .Y(
        n2624) );
  MXT2_X0P5M_A12TR u3352 ( .A(rstkram[358]), .B(wstkw[18]), .S0(n3348), .Y(
        n2623) );
  MXT2_X0P5M_A12TR u3353 ( .A(rstkram[338]), .B(wstkw[18]), .S0(n3349), .Y(
        n2622) );
  MXT2_X0P5M_A12TR u3354 ( .A(rstkram[318]), .B(wstkw[18]), .S0(n3350), .Y(
        n2621) );
  MXT2_X0P5M_A12TR u3355 ( .A(rstkram[298]), .B(wstkw[18]), .S0(n3351), .Y(
        n2620) );
  MXT2_X0P5M_A12TR u3356 ( .A(rstkram[278]), .B(wstkw[18]), .S0(n3352), .Y(
        n2619) );
  MXT2_X0P5M_A12TR u3357 ( .A(rstkram[258]), .B(wstkw[18]), .S0(n3353), .Y(
        n2618) );
  MXT2_X0P5M_A12TR u3358 ( .A(rstkram[238]), .B(wstkw[18]), .S0(n3354), .Y(
        n2617) );
  MXT2_X0P5M_A12TR u3359 ( .A(rstkram[218]), .B(wstkw[18]), .S0(n3355), .Y(
        n2616) );
  MXT2_X0P5M_A12TR u3360 ( .A(rstkram[198]), .B(wstkw[18]), .S0(n3356), .Y(
        n2615) );
  MXT2_X0P5M_A12TR u3361 ( .A(rstkram[178]), .B(wstkw[18]), .S0(n3357), .Y(
        n2614) );
  MXT2_X0P5M_A12TR u3362 ( .A(rstkram[158]), .B(wstkw[18]), .S0(n3358), .Y(
        n2613) );
  MXT2_X0P5M_A12TR u3363 ( .A(rstkram[138]), .B(wstkw[18]), .S0(n3359), .Y(
        n2612) );
  MXT2_X0P5M_A12TR u3364 ( .A(rstkram[118]), .B(wstkw[18]), .S0(n3360), .Y(
        n2611) );
  MXT2_X0P5M_A12TR u3365 ( .A(rstkram[98]), .B(wstkw[18]), .S0(n3361), .Y(
        n2610) );
  MXT2_X0P5M_A12TR u3366 ( .A(rstkram[78]), .B(wstkw[18]), .S0(n3362), .Y(
        n2609) );
  MXT2_X0P5M_A12TR u3367 ( .A(rstkram[58]), .B(wstkw[18]), .S0(n3363), .Y(
        n2608) );
  MXT2_X0P5M_A12TR u3368 ( .A(rstkram[38]), .B(wstkw[18]), .S0(n3364), .Y(
        n2607) );
  MXT2_X0P5M_A12TR u3369 ( .A(rstkram[18]), .B(wstkw[18]), .S0(n3365), .Y(
        n2606) );
  MXT2_X0P5M_A12TR u3370 ( .A(rstkram[639]), .B(wstkw[19]), .S0(n3334), .Y(
        n2605) );
  MXT2_X0P5M_A12TR u3371 ( .A(rstkram[619]), .B(wstkw[19]), .S0(n3335), .Y(
        n2604) );
  MXT2_X0P5M_A12TR u3372 ( .A(rstkram[599]), .B(wstkw[19]), .S0(n3336), .Y(
        n2603) );
  MXT2_X0P5M_A12TR u3373 ( .A(rstkram[579]), .B(wstkw[19]), .S0(n3337), .Y(
        n2602) );
  MXT2_X0P5M_A12TR u3374 ( .A(rstkram[559]), .B(wstkw[19]), .S0(n3338), .Y(
        n2601) );
  MXT2_X0P5M_A12TR u3375 ( .A(rstkram[539]), .B(wstkw[19]), .S0(n3339), .Y(
        n2600) );
  MXT2_X0P5M_A12TR u3376 ( .A(rstkram[519]), .B(wstkw[19]), .S0(n3340), .Y(
        n2599) );
  MXT2_X0P5M_A12TR u3377 ( .A(rstkram[499]), .B(wstkw[19]), .S0(n3341), .Y(
        n2598) );
  MXT2_X0P5M_A12TR u3378 ( .A(rstkram[479]), .B(wstkw[19]), .S0(n3342), .Y(
        n2597) );
  MXT2_X0P5M_A12TR u3379 ( .A(rstkram[459]), .B(wstkw[19]), .S0(n3343), .Y(
        n2596) );
  MXT2_X0P5M_A12TR u3380 ( .A(rstkram[439]), .B(wstkw[19]), .S0(n3344), .Y(
        n2595) );
  MXT2_X0P5M_A12TR u3381 ( .A(rstkram[419]), .B(wstkw[19]), .S0(n3345), .Y(
        n2594) );
  MXT2_X0P5M_A12TR u3382 ( .A(rstkram[399]), .B(wstkw[19]), .S0(n3346), .Y(
        n2593) );
  MXT2_X0P5M_A12TR u3383 ( .A(rstkram[379]), .B(wstkw[19]), .S0(n3347), .Y(
        n2592) );
  MXT2_X0P5M_A12TR u3384 ( .A(rstkram[359]), .B(wstkw[19]), .S0(n3348), .Y(
        n2591) );
  MXT2_X0P5M_A12TR u3385 ( .A(rstkram[339]), .B(wstkw[19]), .S0(n3349), .Y(
        n2590) );
  MXT2_X0P5M_A12TR u3386 ( .A(rstkram[319]), .B(wstkw[19]), .S0(n3350), .Y(
        n2589) );
  MXT2_X0P5M_A12TR u3387 ( .A(rstkram[299]), .B(wstkw[19]), .S0(n3351), .Y(
        n2588) );
  MXT2_X0P5M_A12TR u3388 ( .A(rstkram[279]), .B(wstkw[19]), .S0(n3352), .Y(
        n2587) );
  MXT2_X0P5M_A12TR u3389 ( .A(rstkram[259]), .B(wstkw[19]), .S0(n3353), .Y(
        n2586) );
  MXT2_X0P5M_A12TR u3390 ( .A(rstkram[239]), .B(wstkw[19]), .S0(n3354), .Y(
        n2585) );
  MXT2_X0P5M_A12TR u3391 ( .A(rstkram[219]), .B(wstkw[19]), .S0(n3355), .Y(
        n2584) );
  MXT2_X0P5M_A12TR u3392 ( .A(rstkram[199]), .B(wstkw[19]), .S0(n3356), .Y(
        n2583) );
  MXT2_X0P5M_A12TR u3393 ( .A(rstkram[179]), .B(wstkw[19]), .S0(n3357), .Y(
        n2582) );
  MXT2_X0P5M_A12TR u3394 ( .A(rstkram[159]), .B(wstkw[19]), .S0(n3358), .Y(
        n2581) );
  MXT2_X0P5M_A12TR u3395 ( .A(rstkram[139]), .B(wstkw[19]), .S0(n3359), .Y(
        n2580) );
  MXT2_X0P5M_A12TR u3396 ( .A(rstkram[119]), .B(wstkw[19]), .S0(n3360), .Y(
        n2579) );
  MXT2_X0P5M_A12TR u3397 ( .A(rstkram[99]), .B(wstkw[19]), .S0(n3361), .Y(
        n2578) );
  MXT2_X0P5M_A12TR u3398 ( .A(rstkram[79]), .B(wstkw[19]), .S0(n3362), .Y(
        n2577) );
  MXT2_X0P5M_A12TR u3399 ( .A(rstkram[59]), .B(wstkw[19]), .S0(n3363), .Y(
        n2576) );
  MXT2_X0P5M_A12TR u3400 ( .A(rstkram[39]), .B(wstkw[19]), .S0(n3364), .Y(
        n2575) );
  MXT2_X0P5M_A12TR u3401 ( .A(rstkram[19]), .B(wstkw[19]), .S0(n3365), .Y(
        n2574) );
  MXT2_X0P5M_A12TR u3402 ( .A(rstkram[628]), .B(wstkw[8]), .S0(n3334), .Y(
        n2573) );
  MXT2_X0P5M_A12TR u3403 ( .A(rstkram[608]), .B(wstkw[8]), .S0(n3335), .Y(
        n2572) );
  MXT2_X0P5M_A12TR u3404 ( .A(rstkram[588]), .B(wstkw[8]), .S0(n3336), .Y(
        n2571) );
  MXT2_X0P5M_A12TR u3405 ( .A(rstkram[568]), .B(wstkw[8]), .S0(n3337), .Y(
        n2570) );
  MXT2_X0P5M_A12TR u3406 ( .A(rstkram[548]), .B(wstkw[8]), .S0(n3338), .Y(
        n2569) );
  MXT2_X0P5M_A12TR u3407 ( .A(rstkram[528]), .B(wstkw[8]), .S0(n3339), .Y(
        n2568) );
  MXT2_X0P5M_A12TR u3408 ( .A(rstkram[508]), .B(wstkw[8]), .S0(n3340), .Y(
        n2567) );
  MXT2_X0P5M_A12TR u3409 ( .A(rstkram[488]), .B(wstkw[8]), .S0(n3341), .Y(
        n2566) );
  MXT2_X0P5M_A12TR u3410 ( .A(rstkram[468]), .B(wstkw[8]), .S0(n3342), .Y(
        n2565) );
  MXT2_X0P5M_A12TR u3411 ( .A(rstkram[448]), .B(wstkw[8]), .S0(n3343), .Y(
        n2564) );
  MXT2_X0P5M_A12TR u3412 ( .A(rstkram[428]), .B(wstkw[8]), .S0(n3344), .Y(
        n2563) );
  MXT2_X0P5M_A12TR u3413 ( .A(rstkram[408]), .B(wstkw[8]), .S0(n3345), .Y(
        n2562) );
  MXT2_X0P5M_A12TR u3414 ( .A(rstkram[388]), .B(wstkw[8]), .S0(n3346), .Y(
        n2561) );
  MXT2_X0P5M_A12TR u3415 ( .A(rstkram[368]), .B(wstkw[8]), .S0(n3347), .Y(
        n2560) );
  MXT2_X0P5M_A12TR u3416 ( .A(rstkram[348]), .B(wstkw[8]), .S0(n3348), .Y(
        n2559) );
  MXT2_X0P5M_A12TR u3417 ( .A(rstkram[328]), .B(wstkw[8]), .S0(n3349), .Y(
        n2558) );
  MXT2_X0P5M_A12TR u3418 ( .A(rstkram[308]), .B(wstkw[8]), .S0(n3350), .Y(
        n2557) );
  MXT2_X0P5M_A12TR u3419 ( .A(rstkram[288]), .B(wstkw[8]), .S0(n3351), .Y(
        n2556) );
  MXT2_X0P5M_A12TR u3420 ( .A(rstkram[268]), .B(wstkw[8]), .S0(n3352), .Y(
        n2555) );
  MXT2_X0P5M_A12TR u3421 ( .A(rstkram[248]), .B(wstkw[8]), .S0(n3353), .Y(
        n2554) );
  MXT2_X0P5M_A12TR u3422 ( .A(rstkram[228]), .B(wstkw[8]), .S0(n3354), .Y(
        n2553) );
  MXT2_X0P5M_A12TR u3423 ( .A(rstkram[208]), .B(wstkw[8]), .S0(n3355), .Y(
        n2552) );
  MXT2_X0P5M_A12TR u3424 ( .A(rstkram[188]), .B(wstkw[8]), .S0(n3356), .Y(
        n2551) );
  MXT2_X0P5M_A12TR u3425 ( .A(rstkram[168]), .B(wstkw[8]), .S0(n3357), .Y(
        n2550) );
  MXT2_X0P5M_A12TR u3426 ( .A(rstkram[148]), .B(wstkw[8]), .S0(n3358), .Y(
        n2549) );
  MXT2_X0P5M_A12TR u3427 ( .A(rstkram[128]), .B(wstkw[8]), .S0(n3359), .Y(
        n2548) );
  MXT2_X0P5M_A12TR u3428 ( .A(rstkram[108]), .B(wstkw[8]), .S0(n3360), .Y(
        n2547) );
  MXT2_X0P5M_A12TR u3429 ( .A(rstkram[88]), .B(wstkw[8]), .S0(n3361), .Y(n2546) );
  MXT2_X0P5M_A12TR u3430 ( .A(rstkram[68]), .B(wstkw[8]), .S0(n3362), .Y(n2545) );
  MXT2_X0P5M_A12TR u3431 ( .A(rstkram[48]), .B(wstkw[8]), .S0(n3363), .Y(n2544) );
  MXT2_X0P5M_A12TR u3432 ( .A(rstkram[28]), .B(wstkw[8]), .S0(n3364), .Y(n2543) );
  MXT2_X0P5M_A12TR u3433 ( .A(rstkram[8]), .B(wstkw[8]), .S0(n3365), .Y(n2542)
         );
  MXT2_X0P5M_A12TR u3434 ( .A(rstkram[629]), .B(wstkw[9]), .S0(n3334), .Y(
        n2541) );
  MXT2_X0P5M_A12TR u3435 ( .A(rstkram[609]), .B(wstkw[9]), .S0(n3335), .Y(
        n2540) );
  MXT2_X0P5M_A12TR u3436 ( .A(rstkram[589]), .B(wstkw[9]), .S0(n3336), .Y(
        n2539) );
  MXT2_X0P5M_A12TR u3437 ( .A(rstkram[569]), .B(wstkw[9]), .S0(n3337), .Y(
        n2538) );
  MXT2_X0P5M_A12TR u3438 ( .A(rstkram[549]), .B(wstkw[9]), .S0(n3338), .Y(
        n2537) );
  MXT2_X0P5M_A12TR u3439 ( .A(rstkram[529]), .B(wstkw[9]), .S0(n3339), .Y(
        n2536) );
  MXT2_X0P5M_A12TR u3440 ( .A(rstkram[509]), .B(wstkw[9]), .S0(n3340), .Y(
        n2535) );
  MXT2_X0P5M_A12TR u3441 ( .A(rstkram[489]), .B(wstkw[9]), .S0(n3341), .Y(
        n2534) );
  MXT2_X0P5M_A12TR u3442 ( .A(rstkram[469]), .B(wstkw[9]), .S0(n3342), .Y(
        n2533) );
  MXT2_X0P5M_A12TR u3443 ( .A(rstkram[449]), .B(wstkw[9]), .S0(n3343), .Y(
        n2532) );
  MXT2_X0P5M_A12TR u3444 ( .A(rstkram[429]), .B(wstkw[9]), .S0(n3344), .Y(
        n2531) );
  MXT2_X0P5M_A12TR u3445 ( .A(rstkram[409]), .B(wstkw[9]), .S0(n3345), .Y(
        n2530) );
  MXT2_X0P5M_A12TR u3446 ( .A(rstkram[389]), .B(wstkw[9]), .S0(n3346), .Y(
        n2529) );
  MXT2_X0P5M_A12TR u3447 ( .A(rstkram[369]), .B(wstkw[9]), .S0(n3347), .Y(
        n2528) );
  MXT2_X0P5M_A12TR u3448 ( .A(rstkram[349]), .B(wstkw[9]), .S0(n3348), .Y(
        n2527) );
  MXT2_X0P5M_A12TR u3449 ( .A(rstkram[329]), .B(wstkw[9]), .S0(n3349), .Y(
        n2526) );
  MXT2_X0P5M_A12TR u3450 ( .A(rstkram[309]), .B(wstkw[9]), .S0(n3350), .Y(
        n2525) );
  MXT2_X0P5M_A12TR u3451 ( .A(rstkram[289]), .B(wstkw[9]), .S0(n3351), .Y(
        n2524) );
  MXT2_X0P5M_A12TR u3452 ( .A(rstkram[269]), .B(wstkw[9]), .S0(n3352), .Y(
        n2523) );
  MXT2_X0P5M_A12TR u3453 ( .A(rstkram[249]), .B(wstkw[9]), .S0(n3353), .Y(
        n2522) );
  MXT2_X0P5M_A12TR u3454 ( .A(rstkram[229]), .B(wstkw[9]), .S0(n3354), .Y(
        n2521) );
  MXT2_X0P5M_A12TR u3455 ( .A(rstkram[209]), .B(wstkw[9]), .S0(n3355), .Y(
        n2520) );
  MXT2_X0P5M_A12TR u3456 ( .A(rstkram[189]), .B(wstkw[9]), .S0(n3356), .Y(
        n2519) );
  MXT2_X0P5M_A12TR u3457 ( .A(rstkram[169]), .B(wstkw[9]), .S0(n3357), .Y(
        n2518) );
  MXT2_X0P5M_A12TR u3458 ( .A(rstkram[149]), .B(wstkw[9]), .S0(n3358), .Y(
        n2517) );
  MXT2_X0P5M_A12TR u3459 ( .A(rstkram[129]), .B(wstkw[9]), .S0(n3359), .Y(
        n2516) );
  MXT2_X0P5M_A12TR u3460 ( .A(rstkram[109]), .B(wstkw[9]), .S0(n3360), .Y(
        n2515) );
  MXT2_X0P5M_A12TR u3461 ( .A(rstkram[89]), .B(wstkw[9]), .S0(n3361), .Y(n2514) );
  MXT2_X0P5M_A12TR u3462 ( .A(rstkram[69]), .B(wstkw[9]), .S0(n3362), .Y(n2513) );
  MXT2_X0P5M_A12TR u3463 ( .A(rstkram[49]), .B(wstkw[9]), .S0(n3363), .Y(n2512) );
  MXT2_X0P5M_A12TR u3464 ( .A(rstkram[29]), .B(wstkw[9]), .S0(n3364), .Y(n2511) );
  MXT2_X0P5M_A12TR u3465 ( .A(rstkram[9]), .B(wstkw[9]), .S0(n3365), .Y(n2510)
         );
  MXT2_X0P5M_A12TR u3466 ( .A(rstkram[630]), .B(wstkw[10]), .S0(n3334), .Y(
        n2509) );
  MXT2_X0P5M_A12TR u3467 ( .A(rstkram[610]), .B(wstkw[10]), .S0(n3335), .Y(
        n2508) );
  MXT2_X0P5M_A12TR u3468 ( .A(rstkram[590]), .B(wstkw[10]), .S0(n3336), .Y(
        n2507) );
  MXT2_X0P5M_A12TR u3469 ( .A(rstkram[570]), .B(wstkw[10]), .S0(n3337), .Y(
        n2506) );
  MXT2_X0P5M_A12TR u3470 ( .A(rstkram[550]), .B(wstkw[10]), .S0(n3338), .Y(
        n2505) );
  MXT2_X0P5M_A12TR u3471 ( .A(rstkram[530]), .B(wstkw[10]), .S0(n3339), .Y(
        n2504) );
  MXT2_X0P5M_A12TR u3472 ( .A(rstkram[510]), .B(wstkw[10]), .S0(n3340), .Y(
        n2503) );
  MXT2_X0P5M_A12TR u3473 ( .A(rstkram[490]), .B(wstkw[10]), .S0(n3341), .Y(
        n2502) );
  MXT2_X0P5M_A12TR u3474 ( .A(rstkram[470]), .B(wstkw[10]), .S0(n3342), .Y(
        n2501) );
  MXT2_X0P5M_A12TR u3475 ( .A(rstkram[450]), .B(wstkw[10]), .S0(n3343), .Y(
        n2500) );
  MXT2_X0P5M_A12TR u3476 ( .A(rstkram[430]), .B(wstkw[10]), .S0(n3344), .Y(
        n2499) );
  MXT2_X0P5M_A12TR u3477 ( .A(rstkram[410]), .B(wstkw[10]), .S0(n3345), .Y(
        n2498) );
  MXT2_X0P5M_A12TR u3478 ( .A(rstkram[390]), .B(wstkw[10]), .S0(n3346), .Y(
        n2497) );
  MXT2_X0P5M_A12TR u3479 ( .A(rstkram[370]), .B(wstkw[10]), .S0(n3347), .Y(
        n2496) );
  MXT2_X0P5M_A12TR u3480 ( .A(rstkram[350]), .B(wstkw[10]), .S0(n3348), .Y(
        n2495) );
  MXT2_X0P5M_A12TR u3481 ( .A(rstkram[330]), .B(wstkw[10]), .S0(n3349), .Y(
        n2494) );
  MXT2_X0P5M_A12TR u3482 ( .A(rstkram[310]), .B(wstkw[10]), .S0(n3350), .Y(
        n2493) );
  MXT2_X0P5M_A12TR u3483 ( .A(rstkram[290]), .B(wstkw[10]), .S0(n3351), .Y(
        n2492) );
  MXT2_X0P5M_A12TR u3484 ( .A(rstkram[270]), .B(wstkw[10]), .S0(n3352), .Y(
        n2491) );
  MXT2_X0P5M_A12TR u3485 ( .A(rstkram[250]), .B(wstkw[10]), .S0(n3353), .Y(
        n2490) );
  MXT2_X0P5M_A12TR u3486 ( .A(rstkram[230]), .B(wstkw[10]), .S0(n3354), .Y(
        n2489) );
  MXT2_X0P5M_A12TR u3487 ( .A(rstkram[210]), .B(wstkw[10]), .S0(n3355), .Y(
        n2488) );
  MXT2_X0P5M_A12TR u3488 ( .A(rstkram[190]), .B(wstkw[10]), .S0(n3356), .Y(
        n2487) );
  MXT2_X0P5M_A12TR u3489 ( .A(rstkram[170]), .B(wstkw[10]), .S0(n3357), .Y(
        n2486) );
  MXT2_X0P5M_A12TR u3490 ( .A(rstkram[150]), .B(wstkw[10]), .S0(n3358), .Y(
        n2485) );
  MXT2_X0P5M_A12TR u3491 ( .A(rstkram[130]), .B(wstkw[10]), .S0(n3359), .Y(
        n2484) );
  MXT2_X0P5M_A12TR u3492 ( .A(rstkram[110]), .B(wstkw[10]), .S0(n3360), .Y(
        n2483) );
  MXT2_X0P5M_A12TR u3493 ( .A(rstkram[90]), .B(wstkw[10]), .S0(n3361), .Y(
        n2482) );
  MXT2_X0P5M_A12TR u3494 ( .A(rstkram[70]), .B(wstkw[10]), .S0(n3362), .Y(
        n2481) );
  MXT2_X0P5M_A12TR u3495 ( .A(rstkram[50]), .B(wstkw[10]), .S0(n3363), .Y(
        n2480) );
  MXT2_X0P5M_A12TR u3496 ( .A(rstkram[30]), .B(wstkw[10]), .S0(n3364), .Y(
        n2479) );
  MXT2_X0P5M_A12TR u3497 ( .A(rstkram[10]), .B(wstkw[10]), .S0(n3365), .Y(
        n2478) );
  MXT2_X0P5M_A12TR u3498 ( .A(rstkram[631]), .B(wstkw[11]), .S0(n3334), .Y(
        n2477) );
  MXT2_X0P5M_A12TR u3499 ( .A(rstkram[611]), .B(wstkw[11]), .S0(n3335), .Y(
        n2476) );
  MXT2_X0P5M_A12TR u3500 ( .A(rstkram[591]), .B(wstkw[11]), .S0(n3336), .Y(
        n2475) );
  MXT2_X0P5M_A12TR u3501 ( .A(rstkram[571]), .B(wstkw[11]), .S0(n3337), .Y(
        n2474) );
  MXT2_X0P5M_A12TR u3502 ( .A(rstkram[551]), .B(wstkw[11]), .S0(n3338), .Y(
        n2473) );
  MXT2_X0P5M_A12TR u3503 ( .A(rstkram[531]), .B(wstkw[11]), .S0(n3339), .Y(
        n2472) );
  MXT2_X0P5M_A12TR u3504 ( .A(rstkram[511]), .B(wstkw[11]), .S0(n3340), .Y(
        n2471) );
  MXT2_X0P5M_A12TR u3505 ( .A(rstkram[491]), .B(wstkw[11]), .S0(n3341), .Y(
        n2470) );
  MXT2_X0P5M_A12TR u3506 ( .A(rstkram[471]), .B(wstkw[11]), .S0(n3342), .Y(
        n2469) );
  MXT2_X0P5M_A12TR u3507 ( .A(rstkram[451]), .B(wstkw[11]), .S0(n3343), .Y(
        n2468) );
  MXT2_X0P5M_A12TR u3508 ( .A(rstkram[431]), .B(wstkw[11]), .S0(n3344), .Y(
        n2467) );
  MXT2_X0P5M_A12TR u3509 ( .A(rstkram[411]), .B(wstkw[11]), .S0(n3345), .Y(
        n2466) );
  MXT2_X0P5M_A12TR u3510 ( .A(rstkram[391]), .B(wstkw[11]), .S0(n3346), .Y(
        n2465) );
  MXT2_X0P5M_A12TR u3511 ( .A(rstkram[371]), .B(wstkw[11]), .S0(n3347), .Y(
        n2464) );
  MXT2_X0P5M_A12TR u3512 ( .A(rstkram[351]), .B(wstkw[11]), .S0(n3348), .Y(
        n2463) );
  MXT2_X0P5M_A12TR u3513 ( .A(rstkram[331]), .B(wstkw[11]), .S0(n3349), .Y(
        n2462) );
  MXT2_X0P5M_A12TR u3514 ( .A(rstkram[311]), .B(wstkw[11]), .S0(n3350), .Y(
        n2461) );
  MXT2_X0P5M_A12TR u3515 ( .A(rstkram[291]), .B(wstkw[11]), .S0(n3351), .Y(
        n2460) );
  MXT2_X0P5M_A12TR u3516 ( .A(rstkram[271]), .B(wstkw[11]), .S0(n3352), .Y(
        n2459) );
  MXT2_X0P5M_A12TR u3517 ( .A(rstkram[251]), .B(wstkw[11]), .S0(n3353), .Y(
        n2458) );
  MXT2_X0P5M_A12TR u3518 ( .A(rstkram[231]), .B(wstkw[11]), .S0(n3354), .Y(
        n2457) );
  MXT2_X0P5M_A12TR u3519 ( .A(rstkram[211]), .B(wstkw[11]), .S0(n3355), .Y(
        n2456) );
  MXT2_X0P5M_A12TR u3520 ( .A(rstkram[191]), .B(wstkw[11]), .S0(n3356), .Y(
        n2455) );
  MXT2_X0P5M_A12TR u3521 ( .A(rstkram[171]), .B(wstkw[11]), .S0(n3357), .Y(
        n2454) );
  MXT2_X0P5M_A12TR u3522 ( .A(rstkram[151]), .B(wstkw[11]), .S0(n3358), .Y(
        n2453) );
  MXT2_X0P5M_A12TR u3523 ( .A(rstkram[131]), .B(wstkw[11]), .S0(n3359), .Y(
        n2452) );
  MXT2_X0P5M_A12TR u3524 ( .A(rstkram[111]), .B(wstkw[11]), .S0(n3360), .Y(
        n2451) );
  MXT2_X0P5M_A12TR u3525 ( .A(rstkram[91]), .B(wstkw[11]), .S0(n3361), .Y(
        n2450) );
  MXT2_X0P5M_A12TR u3526 ( .A(rstkram[71]), .B(wstkw[11]), .S0(n3362), .Y(
        n2449) );
  MXT2_X0P5M_A12TR u3527 ( .A(rstkram[51]), .B(wstkw[11]), .S0(n3363), .Y(
        n2448) );
  MXT2_X0P5M_A12TR u3528 ( .A(rstkram[31]), .B(wstkw[11]), .S0(n3364), .Y(
        n2447) );
  MXT2_X0P5M_A12TR u3529 ( .A(rstkram[11]), .B(wstkw[11]), .S0(n3365), .Y(
        n2446) );
  MXT2_X0P5M_A12TR u3530 ( .A(rstkram[632]), .B(wstkw[12]), .S0(n3334), .Y(
        n2445) );
  MXT2_X0P5M_A12TR u3531 ( .A(rstkram[612]), .B(wstkw[12]), .S0(n3335), .Y(
        n2444) );
  MXT2_X0P5M_A12TR u3532 ( .A(rstkram[592]), .B(wstkw[12]), .S0(n3336), .Y(
        n2443) );
  MXT2_X0P5M_A12TR u3533 ( .A(rstkram[572]), .B(wstkw[12]), .S0(n3337), .Y(
        n2442) );
  MXT2_X0P5M_A12TR u3534 ( .A(rstkram[552]), .B(wstkw[12]), .S0(n3338), .Y(
        n2441) );
  MXT2_X0P5M_A12TR u3535 ( .A(rstkram[532]), .B(wstkw[12]), .S0(n3339), .Y(
        n2440) );
  MXT2_X0P5M_A12TR u3536 ( .A(rstkram[512]), .B(wstkw[12]), .S0(n3340), .Y(
        n2439) );
  MXT2_X0P5M_A12TR u3537 ( .A(rstkram[492]), .B(wstkw[12]), .S0(n3341), .Y(
        n2438) );
  MXT2_X0P5M_A12TR u3538 ( .A(rstkram[472]), .B(wstkw[12]), .S0(n3342), .Y(
        n2437) );
  MXT2_X0P5M_A12TR u3539 ( .A(rstkram[452]), .B(wstkw[12]), .S0(n3343), .Y(
        n2436) );
  MXT2_X0P5M_A12TR u3540 ( .A(rstkram[432]), .B(wstkw[12]), .S0(n3344), .Y(
        n2435) );
  MXT2_X0P5M_A12TR u3541 ( .A(rstkram[412]), .B(wstkw[12]), .S0(n3345), .Y(
        n2434) );
  MXT2_X0P5M_A12TR u3542 ( .A(rstkram[392]), .B(wstkw[12]), .S0(n3346), .Y(
        n2433) );
  MXT2_X0P5M_A12TR u3543 ( .A(rstkram[372]), .B(wstkw[12]), .S0(n3347), .Y(
        n2432) );
  MXT2_X0P5M_A12TR u3544 ( .A(rstkram[352]), .B(wstkw[12]), .S0(n3348), .Y(
        n2431) );
  MXT2_X0P5M_A12TR u3545 ( .A(rstkram[332]), .B(wstkw[12]), .S0(n3349), .Y(
        n2430) );
  MXT2_X0P5M_A12TR u3546 ( .A(rstkram[312]), .B(wstkw[12]), .S0(n3350), .Y(
        n2429) );
  MXT2_X0P5M_A12TR u3547 ( .A(rstkram[292]), .B(wstkw[12]), .S0(n3351), .Y(
        n2428) );
  MXT2_X0P5M_A12TR u3548 ( .A(rstkram[272]), .B(wstkw[12]), .S0(n3352), .Y(
        n2427) );
  MXT2_X0P5M_A12TR u3549 ( .A(rstkram[252]), .B(wstkw[12]), .S0(n3353), .Y(
        n2426) );
  MXT2_X0P5M_A12TR u3550 ( .A(rstkram[232]), .B(wstkw[12]), .S0(n3354), .Y(
        n2425) );
  MXT2_X0P5M_A12TR u3551 ( .A(rstkram[212]), .B(wstkw[12]), .S0(n3355), .Y(
        n2424) );
  MXT2_X0P5M_A12TR u3552 ( .A(rstkram[192]), .B(wstkw[12]), .S0(n3356), .Y(
        n2423) );
  MXT2_X0P5M_A12TR u3553 ( .A(rstkram[172]), .B(wstkw[12]), .S0(n3357), .Y(
        n2422) );
  MXT2_X0P5M_A12TR u3554 ( .A(rstkram[152]), .B(wstkw[12]), .S0(n3358), .Y(
        n2421) );
  MXT2_X0P5M_A12TR u3555 ( .A(rstkram[132]), .B(wstkw[12]), .S0(n3359), .Y(
        n2420) );
  MXT2_X0P5M_A12TR u3556 ( .A(rstkram[112]), .B(wstkw[12]), .S0(n3360), .Y(
        n2419) );
  MXT2_X0P5M_A12TR u3557 ( .A(rstkram[92]), .B(wstkw[12]), .S0(n3361), .Y(
        n2418) );
  MXT2_X0P5M_A12TR u3558 ( .A(rstkram[72]), .B(wstkw[12]), .S0(n3362), .Y(
        n2417) );
  MXT2_X0P5M_A12TR u3559 ( .A(rstkram[52]), .B(wstkw[12]), .S0(n3363), .Y(
        n2416) );
  MXT2_X0P5M_A12TR u3560 ( .A(rstkram[32]), .B(wstkw[12]), .S0(n3364), .Y(
        n2415) );
  MXT2_X0P5M_A12TR u3561 ( .A(rstkram[12]), .B(wstkw[12]), .S0(n3365), .Y(
        n2414) );
  MXT2_X0P5M_A12TR u3562 ( .A(rstkram[633]), .B(wstkw[13]), .S0(n3334), .Y(
        n2413) );
  MXT2_X0P5M_A12TR u3563 ( .A(rstkram[613]), .B(wstkw[13]), .S0(n3335), .Y(
        n2412) );
  MXT2_X0P5M_A12TR u3564 ( .A(rstkram[593]), .B(wstkw[13]), .S0(n3336), .Y(
        n2411) );
  MXT2_X0P5M_A12TR u3565 ( .A(rstkram[573]), .B(wstkw[13]), .S0(n3337), .Y(
        n2410) );
  MXT2_X0P5M_A12TR u3566 ( .A(rstkram[553]), .B(wstkw[13]), .S0(n3338), .Y(
        n2409) );
  MXT2_X0P5M_A12TR u3567 ( .A(rstkram[533]), .B(wstkw[13]), .S0(n3339), .Y(
        n2408) );
  MXT2_X0P5M_A12TR u3568 ( .A(rstkram[513]), .B(wstkw[13]), .S0(n3340), .Y(
        n2407) );
  MXT2_X0P5M_A12TR u3569 ( .A(rstkram[493]), .B(wstkw[13]), .S0(n3341), .Y(
        n2406) );
  MXT2_X0P5M_A12TR u3570 ( .A(rstkram[473]), .B(wstkw[13]), .S0(n3342), .Y(
        n2405) );
  MXT2_X0P5M_A12TR u3571 ( .A(rstkram[453]), .B(wstkw[13]), .S0(n3343), .Y(
        n2404) );
  MXT2_X0P5M_A12TR u3572 ( .A(rstkram[433]), .B(wstkw[13]), .S0(n3344), .Y(
        n2403) );
  MXT2_X0P5M_A12TR u3573 ( .A(rstkram[413]), .B(wstkw[13]), .S0(n3345), .Y(
        n2402) );
  MXT2_X0P5M_A12TR u3574 ( .A(rstkram[393]), .B(wstkw[13]), .S0(n3346), .Y(
        n2401) );
  MXT2_X0P5M_A12TR u3575 ( .A(rstkram[373]), .B(wstkw[13]), .S0(n3347), .Y(
        n2400) );
  MXT2_X0P5M_A12TR u3576 ( .A(rstkram[353]), .B(wstkw[13]), .S0(n3348), .Y(
        n2399) );
  MXT2_X0P5M_A12TR u3577 ( .A(rstkram[333]), .B(wstkw[13]), .S0(n3349), .Y(
        n2398) );
  MXT2_X0P5M_A12TR u3578 ( .A(rstkram[313]), .B(wstkw[13]), .S0(n3350), .Y(
        n2397) );
  MXT2_X0P5M_A12TR u3579 ( .A(rstkram[293]), .B(wstkw[13]), .S0(n3351), .Y(
        n2396) );
  MXT2_X0P5M_A12TR u3580 ( .A(rstkram[273]), .B(wstkw[13]), .S0(n3352), .Y(
        n2395) );
  MXT2_X0P5M_A12TR u3581 ( .A(rstkram[253]), .B(wstkw[13]), .S0(n3353), .Y(
        n2394) );
  MXT2_X0P5M_A12TR u3582 ( .A(rstkram[233]), .B(wstkw[13]), .S0(n3354), .Y(
        n2393) );
  MXT2_X0P5M_A12TR u3583 ( .A(rstkram[213]), .B(wstkw[13]), .S0(n3355), .Y(
        n2392) );
  MXT2_X0P5M_A12TR u3584 ( .A(rstkram[193]), .B(wstkw[13]), .S0(n3356), .Y(
        n2391) );
  MXT2_X0P5M_A12TR u3585 ( .A(rstkram[173]), .B(wstkw[13]), .S0(n3357), .Y(
        n2390) );
  MXT2_X0P5M_A12TR u3586 ( .A(rstkram[153]), .B(wstkw[13]), .S0(n3358), .Y(
        n2389) );
  MXT2_X0P5M_A12TR u3587 ( .A(rstkram[133]), .B(wstkw[13]), .S0(n3359), .Y(
        n2388) );
  MXT2_X0P5M_A12TR u3588 ( .A(rstkram[113]), .B(wstkw[13]), .S0(n3360), .Y(
        n2387) );
  MXT2_X0P5M_A12TR u3589 ( .A(rstkram[93]), .B(wstkw[13]), .S0(n3361), .Y(
        n2386) );
  MXT2_X0P5M_A12TR u3590 ( .A(rstkram[73]), .B(wstkw[13]), .S0(n3362), .Y(
        n2385) );
  MXT2_X0P5M_A12TR u3591 ( .A(rstkram[53]), .B(wstkw[13]), .S0(n3363), .Y(
        n2384) );
  MXT2_X0P5M_A12TR u3592 ( .A(rstkram[33]), .B(wstkw[13]), .S0(n3364), .Y(
        n2383) );
  MXT2_X0P5M_A12TR u3593 ( .A(rstkram[13]), .B(wstkw[13]), .S0(n3365), .Y(
        n2382) );
  MXT2_X0P5M_A12TR u3594 ( .A(rstkram[634]), .B(wstkw[14]), .S0(n3334), .Y(
        n2381) );
  MXT2_X0P5M_A12TR u3595 ( .A(rstkram[614]), .B(wstkw[14]), .S0(n3335), .Y(
        n2380) );
  MXT2_X0P5M_A12TR u3596 ( .A(rstkram[594]), .B(wstkw[14]), .S0(n3336), .Y(
        n2379) );
  MXT2_X0P5M_A12TR u3597 ( .A(rstkram[574]), .B(wstkw[14]), .S0(n3337), .Y(
        n2378) );
  MXT2_X0P5M_A12TR u3598 ( .A(rstkram[554]), .B(wstkw[14]), .S0(n3338), .Y(
        n2377) );
  MXT2_X0P5M_A12TR u3599 ( .A(rstkram[534]), .B(wstkw[14]), .S0(n3339), .Y(
        n2376) );
  MXT2_X0P5M_A12TR u3600 ( .A(rstkram[514]), .B(wstkw[14]), .S0(n3340), .Y(
        n2375) );
  MXT2_X0P5M_A12TR u3601 ( .A(rstkram[494]), .B(wstkw[14]), .S0(n3341), .Y(
        n2374) );
  MXT2_X0P5M_A12TR u3602 ( .A(rstkram[474]), .B(wstkw[14]), .S0(n3342), .Y(
        n2373) );
  MXT2_X0P5M_A12TR u3603 ( .A(rstkram[454]), .B(wstkw[14]), .S0(n3343), .Y(
        n2372) );
  MXT2_X0P5M_A12TR u3604 ( .A(rstkram[434]), .B(wstkw[14]), .S0(n3344), .Y(
        n2371) );
  MXT2_X0P5M_A12TR u3605 ( .A(rstkram[414]), .B(wstkw[14]), .S0(n3345), .Y(
        n2370) );
  MXT2_X0P5M_A12TR u3606 ( .A(rstkram[394]), .B(wstkw[14]), .S0(n3346), .Y(
        n2369) );
  MXT2_X0P5M_A12TR u3607 ( .A(rstkram[374]), .B(wstkw[14]), .S0(n3347), .Y(
        n2368) );
  MXT2_X0P5M_A12TR u3608 ( .A(rstkram[354]), .B(wstkw[14]), .S0(n3348), .Y(
        n2367) );
  MXT2_X0P5M_A12TR u3609 ( .A(rstkram[334]), .B(wstkw[14]), .S0(n3349), .Y(
        n2366) );
  MXT2_X0P5M_A12TR u3610 ( .A(rstkram[314]), .B(wstkw[14]), .S0(n3350), .Y(
        n2365) );
  MXT2_X0P5M_A12TR u3611 ( .A(rstkram[294]), .B(wstkw[14]), .S0(n3351), .Y(
        n2364) );
  MXT2_X0P5M_A12TR u3612 ( .A(rstkram[274]), .B(wstkw[14]), .S0(n3352), .Y(
        n2363) );
  MXT2_X0P5M_A12TR u3613 ( .A(rstkram[254]), .B(wstkw[14]), .S0(n3353), .Y(
        n2362) );
  MXT2_X0P5M_A12TR u3614 ( .A(rstkram[234]), .B(wstkw[14]), .S0(n3354), .Y(
        n2361) );
  MXT2_X0P5M_A12TR u3615 ( .A(rstkram[214]), .B(wstkw[14]), .S0(n3355), .Y(
        n2360) );
  MXT2_X0P5M_A12TR u3616 ( .A(rstkram[194]), .B(wstkw[14]), .S0(n3356), .Y(
        n2359) );
  MXT2_X0P5M_A12TR u3617 ( .A(rstkram[174]), .B(wstkw[14]), .S0(n3357), .Y(
        n2358) );
  MXT2_X0P5M_A12TR u3618 ( .A(rstkram[154]), .B(wstkw[14]), .S0(n3358), .Y(
        n2357) );
  MXT2_X0P5M_A12TR u3619 ( .A(rstkram[134]), .B(wstkw[14]), .S0(n3359), .Y(
        n2356) );
  MXT2_X0P5M_A12TR u3620 ( .A(rstkram[114]), .B(wstkw[14]), .S0(n3360), .Y(
        n2355) );
  MXT2_X0P5M_A12TR u3621 ( .A(rstkram[94]), .B(wstkw[14]), .S0(n3361), .Y(
        n2354) );
  MXT2_X0P5M_A12TR u3622 ( .A(rstkram[74]), .B(wstkw[14]), .S0(n3362), .Y(
        n2353) );
  MXT2_X0P5M_A12TR u3623 ( .A(rstkram[54]), .B(wstkw[14]), .S0(n3363), .Y(
        n2352) );
  MXT2_X0P5M_A12TR u3624 ( .A(rstkram[34]), .B(wstkw[14]), .S0(n3364), .Y(
        n2351) );
  MXT2_X0P5M_A12TR u3625 ( .A(rstkram[14]), .B(wstkw[14]), .S0(n3365), .Y(
        n2350) );
  MXT2_X0P5M_A12TR u3626 ( .A(rstkram[635]), .B(wstkw[15]), .S0(n3334), .Y(
        n2349) );
  MXT2_X0P5M_A12TR u3627 ( .A(rstkram[615]), .B(wstkw[15]), .S0(n3335), .Y(
        n2348) );
  MXT2_X0P5M_A12TR u3628 ( .A(rstkram[595]), .B(wstkw[15]), .S0(n3336), .Y(
        n2347) );
  MXT2_X0P5M_A12TR u3629 ( .A(rstkram[575]), .B(wstkw[15]), .S0(n3337), .Y(
        n2346) );
  MXT2_X0P5M_A12TR u3630 ( .A(rstkram[555]), .B(wstkw[15]), .S0(n3338), .Y(
        n2345) );
  MXT2_X0P5M_A12TR u3631 ( .A(rstkram[535]), .B(wstkw[15]), .S0(n3339), .Y(
        n2344) );
  MXT2_X0P5M_A12TR u3632 ( .A(rstkram[515]), .B(wstkw[15]), .S0(n3340), .Y(
        n2343) );
  MXT2_X0P5M_A12TR u3633 ( .A(rstkram[495]), .B(wstkw[15]), .S0(n3341), .Y(
        n2342) );
  MXT2_X0P5M_A12TR u3634 ( .A(rstkram[475]), .B(wstkw[15]), .S0(n3342), .Y(
        n2341) );
  MXT2_X0P5M_A12TR u3635 ( .A(rstkram[455]), .B(wstkw[15]), .S0(n3343), .Y(
        n2340) );
  MXT2_X0P5M_A12TR u3636 ( .A(rstkram[435]), .B(wstkw[15]), .S0(n3344), .Y(
        n2339) );
  MXT2_X0P5M_A12TR u3637 ( .A(rstkram[415]), .B(wstkw[15]), .S0(n3345), .Y(
        n2338) );
  MXT2_X0P5M_A12TR u3638 ( .A(rstkram[395]), .B(wstkw[15]), .S0(n3346), .Y(
        n2337) );
  MXT2_X0P5M_A12TR u3639 ( .A(rstkram[375]), .B(wstkw[15]), .S0(n3347), .Y(
        n2336) );
  MXT2_X0P5M_A12TR u3640 ( .A(rstkram[355]), .B(wstkw[15]), .S0(n3348), .Y(
        n2335) );
  MXT2_X0P5M_A12TR u3641 ( .A(rstkram[335]), .B(wstkw[15]), .S0(n3349), .Y(
        n2334) );
  MXT2_X0P5M_A12TR u3642 ( .A(rstkram[315]), .B(wstkw[15]), .S0(n3350), .Y(
        n2333) );
  MXT2_X0P5M_A12TR u3643 ( .A(rstkram[295]), .B(wstkw[15]), .S0(n3351), .Y(
        n2332) );
  MXT2_X0P5M_A12TR u3644 ( .A(rstkram[275]), .B(wstkw[15]), .S0(n3352), .Y(
        n2331) );
  MXT2_X0P5M_A12TR u3645 ( .A(rstkram[255]), .B(wstkw[15]), .S0(n3353), .Y(
        n2330) );
  MXT2_X0P5M_A12TR u3646 ( .A(rstkram[235]), .B(wstkw[15]), .S0(n3354), .Y(
        n2329) );
  MXT2_X0P5M_A12TR u3647 ( .A(rstkram[215]), .B(wstkw[15]), .S0(n3355), .Y(
        n2328) );
  MXT2_X0P5M_A12TR u3648 ( .A(rstkram[195]), .B(wstkw[15]), .S0(n3356), .Y(
        n2327) );
  MXT2_X0P5M_A12TR u3649 ( .A(rstkram[175]), .B(wstkw[15]), .S0(n3357), .Y(
        n2326) );
  MXT2_X0P5M_A12TR u3650 ( .A(rstkram[155]), .B(wstkw[15]), .S0(n3358), .Y(
        n2325) );
  MXT2_X0P5M_A12TR u3651 ( .A(rstkram[135]), .B(wstkw[15]), .S0(n3359), .Y(
        n2324) );
  MXT2_X0P5M_A12TR u3652 ( .A(rstkram[115]), .B(wstkw[15]), .S0(n3360), .Y(
        n2323) );
  MXT2_X0P5M_A12TR u3653 ( .A(rstkram[95]), .B(wstkw[15]), .S0(n3361), .Y(
        n2322) );
  MXT2_X0P5M_A12TR u3654 ( .A(rstkram[75]), .B(wstkw[15]), .S0(n3362), .Y(
        n2321) );
  MXT2_X0P5M_A12TR u3655 ( .A(rstkram[55]), .B(wstkw[15]), .S0(n3363), .Y(
        n2320) );
  MXT2_X0P5M_A12TR u3656 ( .A(rstkram[35]), .B(wstkw[15]), .S0(n3364), .Y(
        n2319) );
  MXT2_X0P5M_A12TR u3657 ( .A(rstkram[15]), .B(wstkw[15]), .S0(n3365), .Y(
        n2318) );
  MXT2_X0P5M_A12TR u3658 ( .A(rstkram[620]), .B(wstkw[0]), .S0(n3334), .Y(
        n2317) );
  MXT2_X0P5M_A12TR u3659 ( .A(rstkram[600]), .B(wstkw[0]), .S0(n3335), .Y(
        n2316) );
  MXT2_X0P5M_A12TR u3660 ( .A(rstkram[580]), .B(wstkw[0]), .S0(n3336), .Y(
        n2315) );
  MXT2_X0P5M_A12TR u3661 ( .A(rstkram[560]), .B(wstkw[0]), .S0(n3337), .Y(
        n2314) );
  MXT2_X0P5M_A12TR u3662 ( .A(rstkram[540]), .B(wstkw[0]), .S0(n3338), .Y(
        n2313) );
  MXT2_X0P5M_A12TR u3663 ( .A(rstkram[520]), .B(wstkw[0]), .S0(n3339), .Y(
        n2312) );
  MXT2_X0P5M_A12TR u3664 ( .A(rstkram[500]), .B(wstkw[0]), .S0(n3340), .Y(
        n2311) );
  MXT2_X0P5M_A12TR u3665 ( .A(rstkram[480]), .B(wstkw[0]), .S0(n3341), .Y(
        n2310) );
  MXT2_X0P5M_A12TR u3666 ( .A(rstkram[460]), .B(wstkw[0]), .S0(n3342), .Y(
        n2309) );
  MXT2_X0P5M_A12TR u3667 ( .A(rstkram[440]), .B(wstkw[0]), .S0(n3343), .Y(
        n2308) );
  MXT2_X0P5M_A12TR u3668 ( .A(rstkram[420]), .B(wstkw[0]), .S0(n3344), .Y(
        n2307) );
  MXT2_X0P5M_A12TR u3669 ( .A(rstkram[400]), .B(wstkw[0]), .S0(n3345), .Y(
        n2306) );
  MXT2_X0P5M_A12TR u3670 ( .A(rstkram[380]), .B(wstkw[0]), .S0(n3346), .Y(
        n2305) );
  MXT2_X0P5M_A12TR u3671 ( .A(rstkram[360]), .B(wstkw[0]), .S0(n3347), .Y(
        n2304) );
  MXT2_X0P5M_A12TR u3672 ( .A(rstkram[340]), .B(wstkw[0]), .S0(n3348), .Y(
        n2303) );
  MXT2_X0P5M_A12TR u3673 ( .A(rstkram[320]), .B(wstkw[0]), .S0(n3349), .Y(
        n2302) );
  MXT2_X0P5M_A12TR u3674 ( .A(rstkram[300]), .B(wstkw[0]), .S0(n3350), .Y(
        n2301) );
  MXT2_X0P5M_A12TR u3675 ( .A(rstkram[280]), .B(wstkw[0]), .S0(n3351), .Y(
        n2300) );
  MXT2_X0P5M_A12TR u3676 ( .A(rstkram[260]), .B(wstkw[0]), .S0(n3352), .Y(
        n2299) );
  MXT2_X0P5M_A12TR u3677 ( .A(rstkram[240]), .B(wstkw[0]), .S0(n3353), .Y(
        n2298) );
  MXT2_X0P5M_A12TR u3678 ( .A(rstkram[220]), .B(wstkw[0]), .S0(n3354), .Y(
        n2297) );
  MXT2_X0P5M_A12TR u3679 ( .A(rstkram[200]), .B(wstkw[0]), .S0(n3355), .Y(
        n2296) );
  MXT2_X0P5M_A12TR u3680 ( .A(rstkram[180]), .B(wstkw[0]), .S0(n3356), .Y(
        n2295) );
  MXT2_X0P5M_A12TR u3681 ( .A(rstkram[160]), .B(wstkw[0]), .S0(n3357), .Y(
        n2294) );
  MXT2_X0P5M_A12TR u3682 ( .A(rstkram[140]), .B(wstkw[0]), .S0(n3358), .Y(
        n2293) );
  MXT2_X0P5M_A12TR u3683 ( .A(rstkram[120]), .B(wstkw[0]), .S0(n3359), .Y(
        n2292) );
  MXT2_X0P5M_A12TR u3684 ( .A(rstkram[100]), .B(wstkw[0]), .S0(n3360), .Y(
        n2291) );
  MXT2_X0P5M_A12TR u3685 ( .A(rstkram[80]), .B(wstkw[0]), .S0(n3361), .Y(n2290) );
  MXT2_X0P5M_A12TR u3686 ( .A(rstkram[60]), .B(wstkw[0]), .S0(n3362), .Y(n2289) );
  MXT2_X0P5M_A12TR u3687 ( .A(rstkram[40]), .B(wstkw[0]), .S0(n3363), .Y(n2288) );
  MXT2_X0P5M_A12TR u3688 ( .A(rstkram[20]), .B(wstkw[0]), .S0(n3364), .Y(n2287) );
  MXT2_X0P5M_A12TR u3689 ( .A(rstkram[0]), .B(wstkw[0]), .S0(n3365), .Y(n2286)
         );
  MXT2_X0P5M_A12TR u3690 ( .A(rstkram[621]), .B(wstkw[1]), .S0(n3334), .Y(
        n2285) );
  MXT2_X0P5M_A12TR u3691 ( .A(rstkram[601]), .B(wstkw[1]), .S0(n3335), .Y(
        n2284) );
  MXT2_X0P5M_A12TR u3692 ( .A(rstkram[581]), .B(wstkw[1]), .S0(n3336), .Y(
        n2283) );
  MXT2_X0P5M_A12TR u3693 ( .A(rstkram[561]), .B(wstkw[1]), .S0(n3337), .Y(
        n2282) );
  MXT2_X0P5M_A12TR u3694 ( .A(rstkram[541]), .B(wstkw[1]), .S0(n3338), .Y(
        n2281) );
  MXT2_X0P5M_A12TR u3695 ( .A(rstkram[521]), .B(wstkw[1]), .S0(n3339), .Y(
        n2280) );
  MXT2_X0P5M_A12TR u3696 ( .A(rstkram[501]), .B(wstkw[1]), .S0(n3340), .Y(
        n2279) );
  MXT2_X0P5M_A12TR u3697 ( .A(rstkram[481]), .B(wstkw[1]), .S0(n3341), .Y(
        n2278) );
  MXT2_X0P5M_A12TR u3698 ( .A(rstkram[461]), .B(wstkw[1]), .S0(n3342), .Y(
        n2277) );
  MXT2_X0P5M_A12TR u3699 ( .A(rstkram[441]), .B(wstkw[1]), .S0(n3343), .Y(
        n2276) );
  MXT2_X0P5M_A12TR u3700 ( .A(rstkram[421]), .B(wstkw[1]), .S0(n3344), .Y(
        n2275) );
  MXT2_X0P5M_A12TR u3701 ( .A(rstkram[401]), .B(wstkw[1]), .S0(n3345), .Y(
        n2274) );
  MXT2_X0P5M_A12TR u3702 ( .A(rstkram[381]), .B(wstkw[1]), .S0(n3346), .Y(
        n2273) );
  MXT2_X0P5M_A12TR u3703 ( .A(rstkram[361]), .B(wstkw[1]), .S0(n3347), .Y(
        n2272) );
  MXT2_X0P5M_A12TR u3704 ( .A(rstkram[341]), .B(wstkw[1]), .S0(n3348), .Y(
        n2271) );
  MXT2_X0P5M_A12TR u3705 ( .A(rstkram[321]), .B(wstkw[1]), .S0(n3349), .Y(
        n2270) );
  MXT2_X0P5M_A12TR u3706 ( .A(rstkram[301]), .B(wstkw[1]), .S0(n3350), .Y(
        n2269) );
  MXT2_X0P5M_A12TR u3707 ( .A(rstkram[281]), .B(wstkw[1]), .S0(n3351), .Y(
        n2268) );
  MXT2_X0P5M_A12TR u3708 ( .A(rstkram[261]), .B(wstkw[1]), .S0(n3352), .Y(
        n2267) );
  MXT2_X0P5M_A12TR u3709 ( .A(rstkram[241]), .B(wstkw[1]), .S0(n3353), .Y(
        n2266) );
  MXT2_X0P5M_A12TR u3710 ( .A(rstkram[221]), .B(wstkw[1]), .S0(n3354), .Y(
        n2265) );
  MXT2_X0P5M_A12TR u3711 ( .A(rstkram[201]), .B(wstkw[1]), .S0(n3355), .Y(
        n2264) );
  MXT2_X0P5M_A12TR u3712 ( .A(rstkram[181]), .B(wstkw[1]), .S0(n3356), .Y(
        n2263) );
  MXT2_X0P5M_A12TR u3713 ( .A(rstkram[161]), .B(wstkw[1]), .S0(n3357), .Y(
        n2262) );
  MXT2_X0P5M_A12TR u3714 ( .A(rstkram[141]), .B(wstkw[1]), .S0(n3358), .Y(
        n2261) );
  MXT2_X0P5M_A12TR u3715 ( .A(rstkram[121]), .B(wstkw[1]), .S0(n3359), .Y(
        n2260) );
  MXT2_X0P5M_A12TR u3716 ( .A(rstkram[101]), .B(wstkw[1]), .S0(n3360), .Y(
        n2259) );
  MXT2_X0P5M_A12TR u3717 ( .A(rstkram[81]), .B(wstkw[1]), .S0(n3361), .Y(n2258) );
  MXT2_X0P5M_A12TR u3718 ( .A(rstkram[61]), .B(wstkw[1]), .S0(n3362), .Y(n2257) );
  MXT2_X0P5M_A12TR u3719 ( .A(rstkram[41]), .B(wstkw[1]), .S0(n3363), .Y(n2256) );
  MXT2_X0P5M_A12TR u3720 ( .A(rstkram[21]), .B(wstkw[1]), .S0(n3364), .Y(n2255) );
  MXT2_X0P5M_A12TR u3721 ( .A(rstkram[1]), .B(wstkw[1]), .S0(n3365), .Y(n2254)
         );
  MXT2_X0P5M_A12TR u3722 ( .A(rstkram[622]), .B(wstkw[2]), .S0(n3334), .Y(
        n2253) );
  MXT2_X0P5M_A12TR u3723 ( .A(rstkram[602]), .B(wstkw[2]), .S0(n3335), .Y(
        n2252) );
  MXT2_X0P5M_A12TR u3724 ( .A(rstkram[582]), .B(wstkw[2]), .S0(n3336), .Y(
        n2251) );
  MXT2_X0P5M_A12TR u3725 ( .A(rstkram[562]), .B(wstkw[2]), .S0(n3337), .Y(
        n2250) );
  MXT2_X0P5M_A12TR u3726 ( .A(rstkram[542]), .B(wstkw[2]), .S0(n3338), .Y(
        n2249) );
  MXT2_X0P5M_A12TR u3727 ( .A(rstkram[522]), .B(wstkw[2]), .S0(n3339), .Y(
        n2248) );
  MXT2_X0P5M_A12TR u3728 ( .A(rstkram[502]), .B(wstkw[2]), .S0(n3340), .Y(
        n2247) );
  MXT2_X0P5M_A12TR u3729 ( .A(rstkram[482]), .B(wstkw[2]), .S0(n3341), .Y(
        n2246) );
  MXT2_X0P5M_A12TR u3730 ( .A(rstkram[462]), .B(wstkw[2]), .S0(n3342), .Y(
        n2245) );
  MXT2_X0P5M_A12TR u3731 ( .A(rstkram[442]), .B(wstkw[2]), .S0(n3343), .Y(
        n2244) );
  MXT2_X0P5M_A12TR u3732 ( .A(rstkram[422]), .B(wstkw[2]), .S0(n3344), .Y(
        n2243) );
  MXT2_X0P5M_A12TR u3733 ( .A(rstkram[402]), .B(wstkw[2]), .S0(n3345), .Y(
        n2242) );
  MXT2_X0P5M_A12TR u3734 ( .A(rstkram[382]), .B(wstkw[2]), .S0(n3346), .Y(
        n2241) );
  MXT2_X0P5M_A12TR u3735 ( .A(rstkram[362]), .B(wstkw[2]), .S0(n3347), .Y(
        n2240) );
  MXT2_X0P5M_A12TR u3736 ( .A(rstkram[342]), .B(wstkw[2]), .S0(n3348), .Y(
        n2239) );
  MXT2_X0P5M_A12TR u3737 ( .A(rstkram[322]), .B(wstkw[2]), .S0(n3349), .Y(
        n2238) );
  MXT2_X0P5M_A12TR u3738 ( .A(rstkram[302]), .B(wstkw[2]), .S0(n3350), .Y(
        n2237) );
  MXT2_X0P5M_A12TR u3739 ( .A(rstkram[282]), .B(wstkw[2]), .S0(n3351), .Y(
        n2236) );
  MXT2_X0P5M_A12TR u3740 ( .A(rstkram[262]), .B(wstkw[2]), .S0(n3352), .Y(
        n2235) );
  MXT2_X0P5M_A12TR u3741 ( .A(rstkram[242]), .B(wstkw[2]), .S0(n3353), .Y(
        n2234) );
  MXT2_X0P5M_A12TR u3742 ( .A(rstkram[222]), .B(wstkw[2]), .S0(n3354), .Y(
        n2233) );
  MXT2_X0P5M_A12TR u3743 ( .A(rstkram[202]), .B(wstkw[2]), .S0(n3355), .Y(
        n2232) );
  MXT2_X0P5M_A12TR u3744 ( .A(rstkram[182]), .B(wstkw[2]), .S0(n3356), .Y(
        n2231) );
  MXT2_X0P5M_A12TR u3745 ( .A(rstkram[162]), .B(wstkw[2]), .S0(n3357), .Y(
        n2230) );
  MXT2_X0P5M_A12TR u3746 ( .A(rstkram[142]), .B(wstkw[2]), .S0(n3358), .Y(
        n2229) );
  MXT2_X0P5M_A12TR u3747 ( .A(rstkram[122]), .B(wstkw[2]), .S0(n3359), .Y(
        n2228) );
  MXT2_X0P5M_A12TR u3748 ( .A(rstkram[102]), .B(wstkw[2]), .S0(n3360), .Y(
        n2227) );
  MXT2_X0P5M_A12TR u3749 ( .A(rstkram[82]), .B(wstkw[2]), .S0(n3361), .Y(n2226) );
  MXT2_X0P5M_A12TR u3750 ( .A(rstkram[62]), .B(wstkw[2]), .S0(n3362), .Y(n2225) );
  MXT2_X0P5M_A12TR u3751 ( .A(rstkram[42]), .B(wstkw[2]), .S0(n3363), .Y(n2224) );
  MXT2_X0P5M_A12TR u3752 ( .A(rstkram[22]), .B(wstkw[2]), .S0(n3364), .Y(n2223) );
  MXT2_X0P5M_A12TR u3753 ( .A(rstkram[2]), .B(wstkw[2]), .S0(n3365), .Y(n2222)
         );
  MXT2_X0P5M_A12TR u3754 ( .A(rstkram[623]), .B(wstkw[3]), .S0(n3334), .Y(
        n2221) );
  MXT2_X0P5M_A12TR u3755 ( .A(rstkram[603]), .B(wstkw[3]), .S0(n3335), .Y(
        n2220) );
  MXT2_X0P5M_A12TR u3756 ( .A(rstkram[583]), .B(wstkw[3]), .S0(n3336), .Y(
        n2219) );
  MXT2_X0P5M_A12TR u3757 ( .A(rstkram[563]), .B(wstkw[3]), .S0(n3337), .Y(
        n2218) );
  MXT2_X0P5M_A12TR u3758 ( .A(rstkram[543]), .B(wstkw[3]), .S0(n3338), .Y(
        n2217) );
  MXT2_X0P5M_A12TR u3759 ( .A(rstkram[523]), .B(wstkw[3]), .S0(n3339), .Y(
        n2216) );
  MXT2_X0P5M_A12TR u3760 ( .A(rstkram[503]), .B(wstkw[3]), .S0(n3340), .Y(
        n2215) );
  MXT2_X0P5M_A12TR u3761 ( .A(rstkram[483]), .B(wstkw[3]), .S0(n3341), .Y(
        n2214) );
  MXT2_X0P5M_A12TR u3762 ( .A(rstkram[463]), .B(wstkw[3]), .S0(n3342), .Y(
        n2213) );
  MXT2_X0P5M_A12TR u3763 ( .A(rstkram[443]), .B(wstkw[3]), .S0(n3343), .Y(
        n2212) );
  MXT2_X0P5M_A12TR u3764 ( .A(rstkram[423]), .B(wstkw[3]), .S0(n3344), .Y(
        n2211) );
  MXT2_X0P5M_A12TR u3765 ( .A(rstkram[403]), .B(wstkw[3]), .S0(n3345), .Y(
        n2210) );
  MXT2_X0P5M_A12TR u3766 ( .A(rstkram[383]), .B(wstkw[3]), .S0(n3346), .Y(
        n2209) );
  MXT2_X0P5M_A12TR u3767 ( .A(rstkram[363]), .B(wstkw[3]), .S0(n3347), .Y(
        n2208) );
  MXT2_X0P5M_A12TR u3768 ( .A(rstkram[343]), .B(wstkw[3]), .S0(n3348), .Y(
        n2207) );
  MXT2_X0P5M_A12TR u3769 ( .A(rstkram[323]), .B(wstkw[3]), .S0(n3349), .Y(
        n2206) );
  MXT2_X0P5M_A12TR u3770 ( .A(rstkram[303]), .B(wstkw[3]), .S0(n3350), .Y(
        n2205) );
  MXT2_X0P5M_A12TR u3771 ( .A(rstkram[283]), .B(wstkw[3]), .S0(n3351), .Y(
        n2204) );
  MXT2_X0P5M_A12TR u3772 ( .A(rstkram[263]), .B(wstkw[3]), .S0(n3352), .Y(
        n2203) );
  MXT2_X0P5M_A12TR u3773 ( .A(rstkram[243]), .B(wstkw[3]), .S0(n3353), .Y(
        n2202) );
  MXT2_X0P5M_A12TR u3774 ( .A(rstkram[223]), .B(wstkw[3]), .S0(n3354), .Y(
        n2201) );
  MXT2_X0P5M_A12TR u3775 ( .A(rstkram[203]), .B(wstkw[3]), .S0(n3355), .Y(
        n2200) );
  MXT2_X0P5M_A12TR u3776 ( .A(rstkram[183]), .B(wstkw[3]), .S0(n3356), .Y(
        n2199) );
  MXT2_X0P5M_A12TR u3777 ( .A(rstkram[163]), .B(wstkw[3]), .S0(n3357), .Y(
        n2198) );
  MXT2_X0P5M_A12TR u3778 ( .A(rstkram[143]), .B(wstkw[3]), .S0(n3358), .Y(
        n2197) );
  MXT2_X0P5M_A12TR u3779 ( .A(rstkram[123]), .B(wstkw[3]), .S0(n3359), .Y(
        n2196) );
  MXT2_X0P5M_A12TR u3780 ( .A(rstkram[103]), .B(wstkw[3]), .S0(n3360), .Y(
        n2195) );
  MXT2_X0P5M_A12TR u3781 ( .A(rstkram[83]), .B(wstkw[3]), .S0(n3361), .Y(n2194) );
  MXT2_X0P5M_A12TR u3782 ( .A(rstkram[63]), .B(wstkw[3]), .S0(n3362), .Y(n2193) );
  MXT2_X0P5M_A12TR u3783 ( .A(rstkram[43]), .B(wstkw[3]), .S0(n3363), .Y(n2192) );
  MXT2_X0P5M_A12TR u3784 ( .A(rstkram[23]), .B(wstkw[3]), .S0(n3364), .Y(n2191) );
  MXT2_X0P5M_A12TR u3785 ( .A(rstkram[3]), .B(wstkw[3]), .S0(n3365), .Y(n2190)
         );
  MXT2_X0P5M_A12TR u3786 ( .A(rstkram[624]), .B(wstkw[4]), .S0(n3334), .Y(
        n2189) );
  MXT2_X0P5M_A12TR u3787 ( .A(rstkram[604]), .B(wstkw[4]), .S0(n3335), .Y(
        n2188) );
  MXT2_X0P5M_A12TR u3788 ( .A(rstkram[584]), .B(wstkw[4]), .S0(n3336), .Y(
        n2187) );
  MXT2_X0P5M_A12TR u3789 ( .A(rstkram[564]), .B(wstkw[4]), .S0(n3337), .Y(
        n2186) );
  MXT2_X0P5M_A12TR u3790 ( .A(rstkram[544]), .B(wstkw[4]), .S0(n3338), .Y(
        n2185) );
  MXT2_X0P5M_A12TR u3791 ( .A(rstkram[524]), .B(wstkw[4]), .S0(n3339), .Y(
        n2184) );
  MXT2_X0P5M_A12TR u3792 ( .A(rstkram[504]), .B(wstkw[4]), .S0(n3340), .Y(
        n2183) );
  MXT2_X0P5M_A12TR u3793 ( .A(rstkram[484]), .B(wstkw[4]), .S0(n3341), .Y(
        n2182) );
  MXT2_X0P5M_A12TR u3794 ( .A(rstkram[464]), .B(wstkw[4]), .S0(n3342), .Y(
        n2181) );
  MXT2_X0P5M_A12TR u3795 ( .A(rstkram[444]), .B(wstkw[4]), .S0(n3343), .Y(
        n2180) );
  MXT2_X0P5M_A12TR u3796 ( .A(rstkram[424]), .B(wstkw[4]), .S0(n3344), .Y(
        n2179) );
  MXT2_X0P5M_A12TR u3797 ( .A(rstkram[404]), .B(wstkw[4]), .S0(n3345), .Y(
        n2178) );
  MXT2_X0P5M_A12TR u3798 ( .A(rstkram[384]), .B(wstkw[4]), .S0(n3346), .Y(
        n2177) );
  MXT2_X0P5M_A12TR u3799 ( .A(rstkram[364]), .B(wstkw[4]), .S0(n3347), .Y(
        n2176) );
  MXT2_X0P5M_A12TR u3800 ( .A(rstkram[344]), .B(wstkw[4]), .S0(n3348), .Y(
        n2175) );
  MXT2_X0P5M_A12TR u3801 ( .A(rstkram[324]), .B(wstkw[4]), .S0(n3349), .Y(
        n2174) );
  MXT2_X0P5M_A12TR u3802 ( .A(rstkram[304]), .B(wstkw[4]), .S0(n3350), .Y(
        n2173) );
  MXT2_X0P5M_A12TR u3803 ( .A(rstkram[284]), .B(wstkw[4]), .S0(n3351), .Y(
        n2172) );
  MXT2_X0P5M_A12TR u3804 ( .A(rstkram[264]), .B(wstkw[4]), .S0(n3352), .Y(
        n2171) );
  MXT2_X0P5M_A12TR u3805 ( .A(rstkram[244]), .B(wstkw[4]), .S0(n3353), .Y(
        n2170) );
  MXT2_X0P5M_A12TR u3806 ( .A(rstkram[224]), .B(wstkw[4]), .S0(n3354), .Y(
        n2169) );
  MXT2_X0P5M_A12TR u3807 ( .A(rstkram[204]), .B(wstkw[4]), .S0(n3355), .Y(
        n2168) );
  MXT2_X0P5M_A12TR u3808 ( .A(rstkram[184]), .B(wstkw[4]), .S0(n3356), .Y(
        n2167) );
  MXT2_X0P5M_A12TR u3809 ( .A(rstkram[164]), .B(wstkw[4]), .S0(n3357), .Y(
        n2166) );
  MXT2_X0P5M_A12TR u3810 ( .A(rstkram[144]), .B(wstkw[4]), .S0(n3358), .Y(
        n2165) );
  MXT2_X0P5M_A12TR u3811 ( .A(rstkram[124]), .B(wstkw[4]), .S0(n3359), .Y(
        n2164) );
  MXT2_X0P5M_A12TR u3812 ( .A(rstkram[104]), .B(wstkw[4]), .S0(n3360), .Y(
        n2163) );
  MXT2_X0P5M_A12TR u3813 ( .A(rstkram[84]), .B(wstkw[4]), .S0(n3361), .Y(n2162) );
  MXT2_X0P5M_A12TR u3814 ( .A(rstkram[64]), .B(wstkw[4]), .S0(n3362), .Y(n2161) );
  MXT2_X0P5M_A12TR u3815 ( .A(rstkram[44]), .B(wstkw[4]), .S0(n3363), .Y(n2160) );
  MXT2_X0P5M_A12TR u3816 ( .A(rstkram[24]), .B(wstkw[4]), .S0(n3364), .Y(n2159) );
  MXT2_X0P5M_A12TR u3817 ( .A(rstkram[4]), .B(wstkw[4]), .S0(n3365), .Y(n2158)
         );
  MXT2_X0P5M_A12TR u3818 ( .A(rstkram[625]), .B(wstkw[5]), .S0(n3334), .Y(
        n2157) );
  MXT2_X0P5M_A12TR u3819 ( .A(rstkram[605]), .B(wstkw[5]), .S0(n3335), .Y(
        n2156) );
  MXT2_X0P5M_A12TR u3820 ( .A(rstkram[585]), .B(wstkw[5]), .S0(n3336), .Y(
        n2155) );
  MXT2_X0P5M_A12TR u3821 ( .A(rstkram[565]), .B(wstkw[5]), .S0(n3337), .Y(
        n2154) );
  MXT2_X0P5M_A12TR u3822 ( .A(rstkram[545]), .B(wstkw[5]), .S0(n3338), .Y(
        n2153) );
  MXT2_X0P5M_A12TR u3823 ( .A(rstkram[525]), .B(wstkw[5]), .S0(n3339), .Y(
        n2152) );
  MXT2_X0P5M_A12TR u3824 ( .A(rstkram[505]), .B(wstkw[5]), .S0(n3340), .Y(
        n2151) );
  MXT2_X0P5M_A12TR u3825 ( .A(rstkram[485]), .B(wstkw[5]), .S0(n3341), .Y(
        n2150) );
  MXT2_X0P5M_A12TR u3826 ( .A(rstkram[465]), .B(wstkw[5]), .S0(n3342), .Y(
        n2149) );
  MXT2_X0P5M_A12TR u3827 ( .A(rstkram[445]), .B(wstkw[5]), .S0(n3343), .Y(
        n2148) );
  MXT2_X0P5M_A12TR u3828 ( .A(rstkram[425]), .B(wstkw[5]), .S0(n3344), .Y(
        n2147) );
  MXT2_X0P5M_A12TR u3829 ( .A(rstkram[405]), .B(wstkw[5]), .S0(n3345), .Y(
        n2146) );
  MXT2_X0P5M_A12TR u3830 ( .A(rstkram[385]), .B(wstkw[5]), .S0(n3346), .Y(
        n2145) );
  MXT2_X0P5M_A12TR u3831 ( .A(rstkram[365]), .B(wstkw[5]), .S0(n3347), .Y(
        n2144) );
  MXT2_X0P5M_A12TR u3832 ( .A(rstkram[345]), .B(wstkw[5]), .S0(n3348), .Y(
        n2143) );
  MXT2_X0P5M_A12TR u3833 ( .A(rstkram[325]), .B(wstkw[5]), .S0(n3349), .Y(
        n2142) );
  MXT2_X0P5M_A12TR u3834 ( .A(rstkram[305]), .B(wstkw[5]), .S0(n3350), .Y(
        n2141) );
  MXT2_X0P5M_A12TR u3835 ( .A(rstkram[285]), .B(wstkw[5]), .S0(n3351), .Y(
        n2140) );
  MXT2_X0P5M_A12TR u3836 ( .A(rstkram[265]), .B(wstkw[5]), .S0(n3352), .Y(
        n2139) );
  MXT2_X0P5M_A12TR u3837 ( .A(rstkram[245]), .B(wstkw[5]), .S0(n3353), .Y(
        n2138) );
  MXT2_X0P5M_A12TR u3838 ( .A(rstkram[225]), .B(wstkw[5]), .S0(n3354), .Y(
        n2137) );
  MXT2_X0P5M_A12TR u3839 ( .A(rstkram[205]), .B(wstkw[5]), .S0(n3355), .Y(
        n2136) );
  MXT2_X0P5M_A12TR u3840 ( .A(rstkram[185]), .B(wstkw[5]), .S0(n3356), .Y(
        n2135) );
  MXT2_X0P5M_A12TR u3841 ( .A(rstkram[165]), .B(wstkw[5]), .S0(n3357), .Y(
        n2134) );
  MXT2_X0P5M_A12TR u3842 ( .A(rstkram[145]), .B(wstkw[5]), .S0(n3358), .Y(
        n2133) );
  MXT2_X0P5M_A12TR u3843 ( .A(rstkram[125]), .B(wstkw[5]), .S0(n3359), .Y(
        n2132) );
  MXT2_X0P5M_A12TR u3844 ( .A(rstkram[105]), .B(wstkw[5]), .S0(n3360), .Y(
        n2131) );
  MXT2_X0P5M_A12TR u3845 ( .A(rstkram[85]), .B(wstkw[5]), .S0(n3361), .Y(n2130) );
  MXT2_X0P5M_A12TR u3846 ( .A(rstkram[65]), .B(wstkw[5]), .S0(n3362), .Y(n2129) );
  MXT2_X0P5M_A12TR u3847 ( .A(rstkram[45]), .B(wstkw[5]), .S0(n3363), .Y(n2128) );
  MXT2_X0P5M_A12TR u3848 ( .A(rstkram[25]), .B(wstkw[5]), .S0(n3364), .Y(n2127) );
  MXT2_X0P5M_A12TR u3849 ( .A(rstkram[5]), .B(wstkw[5]), .S0(n3365), .Y(n2126)
         );
  MXT2_X0P5M_A12TR u3850 ( .A(rstkram[626]), .B(wstkw[6]), .S0(n3334), .Y(
        n2125) );
  MXT2_X0P5M_A12TR u3851 ( .A(rstkram[606]), .B(wstkw[6]), .S0(n3335), .Y(
        n2124) );
  MXT2_X0P5M_A12TR u3852 ( .A(rstkram[586]), .B(wstkw[6]), .S0(n3336), .Y(
        n2123) );
  MXT2_X0P5M_A12TR u3853 ( .A(rstkram[566]), .B(wstkw[6]), .S0(n3337), .Y(
        n2122) );
  MXT2_X0P5M_A12TR u3854 ( .A(rstkram[546]), .B(wstkw[6]), .S0(n3338), .Y(
        n2121) );
  MXT2_X0P5M_A12TR u3855 ( .A(rstkram[526]), .B(wstkw[6]), .S0(n3339), .Y(
        n2120) );
  MXT2_X0P5M_A12TR u3856 ( .A(rstkram[506]), .B(wstkw[6]), .S0(n3340), .Y(
        n2119) );
  MXT2_X0P5M_A12TR u3857 ( .A(rstkram[486]), .B(wstkw[6]), .S0(n3341), .Y(
        n2118) );
  MXT2_X0P5M_A12TR u3858 ( .A(rstkram[466]), .B(wstkw[6]), .S0(n3342), .Y(
        n2117) );
  MXT2_X0P5M_A12TR u3859 ( .A(rstkram[446]), .B(wstkw[6]), .S0(n3343), .Y(
        n2116) );
  MXT2_X0P5M_A12TR u3860 ( .A(rstkram[426]), .B(wstkw[6]), .S0(n3344), .Y(
        n2115) );
  MXT2_X0P5M_A12TR u3861 ( .A(rstkram[406]), .B(wstkw[6]), .S0(n3345), .Y(
        n2114) );
  MXT2_X0P5M_A12TR u3862 ( .A(rstkram[386]), .B(wstkw[6]), .S0(n3346), .Y(
        n2113) );
  MXT2_X0P5M_A12TR u3863 ( .A(rstkram[366]), .B(wstkw[6]), .S0(n3347), .Y(
        n2112) );
  MXT2_X0P5M_A12TR u3864 ( .A(rstkram[346]), .B(wstkw[6]), .S0(n3348), .Y(
        n2111) );
  MXT2_X0P5M_A12TR u3865 ( .A(rstkram[326]), .B(wstkw[6]), .S0(n3349), .Y(
        n2110) );
  MXT2_X0P5M_A12TR u3866 ( .A(rstkram[306]), .B(wstkw[6]), .S0(n3350), .Y(
        n2109) );
  MXT2_X0P5M_A12TR u3867 ( .A(rstkram[286]), .B(wstkw[6]), .S0(n3351), .Y(
        n2108) );
  MXT2_X0P5M_A12TR u3868 ( .A(rstkram[266]), .B(wstkw[6]), .S0(n3352), .Y(
        n2107) );
  MXT2_X0P5M_A12TR u3869 ( .A(rstkram[246]), .B(wstkw[6]), .S0(n3353), .Y(
        n2106) );
  MXT2_X0P5M_A12TR u3870 ( .A(rstkram[226]), .B(wstkw[6]), .S0(n3354), .Y(
        n2105) );
  MXT2_X0P5M_A12TR u3871 ( .A(rstkram[206]), .B(wstkw[6]), .S0(n3355), .Y(
        n2104) );
  MXT2_X0P5M_A12TR u3872 ( .A(rstkram[186]), .B(wstkw[6]), .S0(n3356), .Y(
        n2103) );
  MXT2_X0P5M_A12TR u3873 ( .A(rstkram[166]), .B(wstkw[6]), .S0(n3357), .Y(
        n2102) );
  MXT2_X0P5M_A12TR u3874 ( .A(rstkram[146]), .B(wstkw[6]), .S0(n3358), .Y(
        n2101) );
  MXT2_X0P5M_A12TR u3875 ( .A(rstkram[126]), .B(wstkw[6]), .S0(n3359), .Y(
        n2100) );
  MXT2_X0P5M_A12TR u3876 ( .A(rstkram[106]), .B(wstkw[6]), .S0(n3360), .Y(
        n2099) );
  MXT2_X0P5M_A12TR u3877 ( .A(rstkram[86]), .B(wstkw[6]), .S0(n3361), .Y(n2098) );
  MXT2_X0P5M_A12TR u3878 ( .A(rstkram[66]), .B(wstkw[6]), .S0(n3362), .Y(n2097) );
  MXT2_X0P5M_A12TR u3879 ( .A(rstkram[46]), .B(wstkw[6]), .S0(n3363), .Y(n2096) );
  MXT2_X0P5M_A12TR u3880 ( .A(rstkram[26]), .B(wstkw[6]), .S0(n3364), .Y(n2095) );
  MXT2_X0P5M_A12TR u3881 ( .A(rstkram[6]), .B(wstkw[6]), .S0(n3365), .Y(n2094)
         );
  MXT2_X0P5M_A12TR u3882 ( .A(rstkram[627]), .B(wstkw[7]), .S0(n3334), .Y(
        n2093) );
  AND2_X0P5M_A12TR u3883 ( .A(n3366), .B(n3367), .Y(n3334) );
  MXT2_X0P5M_A12TR u3884 ( .A(rstkram[607]), .B(wstkw[7]), .S0(n3335), .Y(
        n2092) );
  AND2_X0P5M_A12TR u3885 ( .A(n3368), .B(n3367), .Y(n3335) );
  MXT2_X0P5M_A12TR u3886 ( .A(rstkram[587]), .B(wstkw[7]), .S0(n3336), .Y(
        n2091) );
  AND2_X0P5M_A12TR u3887 ( .A(n3369), .B(n3367), .Y(n3336) );
  MXT2_X0P5M_A12TR u3888 ( .A(rstkram[567]), .B(wstkw[7]), .S0(n3337), .Y(
        n2090) );
  AND2_X0P5M_A12TR u3889 ( .A(n3370), .B(n3367), .Y(n3337) );
  MXT2_X0P5M_A12TR u3890 ( .A(rstkram[547]), .B(wstkw[7]), .S0(n3338), .Y(
        n2089) );
  AND2_X0P5M_A12TR u3891 ( .A(n3371), .B(n3367), .Y(n3338) );
  MXT2_X0P5M_A12TR u3892 ( .A(rstkram[527]), .B(wstkw[7]), .S0(n3339), .Y(
        n2088) );
  AND2_X0P5M_A12TR u3893 ( .A(n3372), .B(n3367), .Y(n3339) );
  MXT2_X0P5M_A12TR u3894 ( .A(rstkram[507]), .B(wstkw[7]), .S0(n3340), .Y(
        n2087) );
  AND2_X0P5M_A12TR u3895 ( .A(n3373), .B(n3367), .Y(n3340) );
  MXT2_X0P5M_A12TR u3896 ( .A(rstkram[487]), .B(wstkw[7]), .S0(n3341), .Y(
        n2086) );
  AND2_X0P5M_A12TR u3897 ( .A(n3374), .B(n3367), .Y(n3341) );
  NOR3_X0P5A_A12TR u3898 ( .A(rstkptr_[3]), .B(rstkptr_[4]), .C(n3375), .Y(
        n3367) );
  MXT2_X0P5M_A12TR u3899 ( .A(rstkram[467]), .B(wstkw[7]), .S0(n3342), .Y(
        n2085) );
  AND2_X0P5M_A12TR u3900 ( .A(n3376), .B(n3366), .Y(n3342) );
  MXT2_X0P5M_A12TR u3901 ( .A(rstkram[447]), .B(wstkw[7]), .S0(n3343), .Y(
        n2084) );
  AND2_X0P5M_A12TR u3902 ( .A(n3376), .B(n3368), .Y(n3343) );
  MXT2_X0P5M_A12TR u3903 ( .A(rstkram[427]), .B(wstkw[7]), .S0(n3344), .Y(
        n2083) );
  AND2_X0P5M_A12TR u3904 ( .A(n3376), .B(n3369), .Y(n3344) );
  MXT2_X0P5M_A12TR u3905 ( .A(rstkram[407]), .B(wstkw[7]), .S0(n3345), .Y(
        n2082) );
  AND2_X0P5M_A12TR u3906 ( .A(n3376), .B(n3370), .Y(n3345) );
  MXT2_X0P5M_A12TR u3907 ( .A(rstkram[387]), .B(wstkw[7]), .S0(n3346), .Y(
        n2081) );
  AND2_X0P5M_A12TR u3908 ( .A(n3376), .B(n3371), .Y(n3346) );
  MXT2_X0P5M_A12TR u3909 ( .A(rstkram[367]), .B(wstkw[7]), .S0(n3347), .Y(
        n2080) );
  AND2_X0P5M_A12TR u3910 ( .A(n3376), .B(n3372), .Y(n3347) );
  MXT2_X0P5M_A12TR u3911 ( .A(rstkram[347]), .B(wstkw[7]), .S0(n3348), .Y(
        n2079) );
  AND2_X0P5M_A12TR u3912 ( .A(n3376), .B(n3373), .Y(n3348) );
  MXT2_X0P5M_A12TR u3913 ( .A(rstkram[327]), .B(wstkw[7]), .S0(n3349), .Y(
        n2078) );
  AND2_X0P5M_A12TR u3914 ( .A(n3376), .B(n3374), .Y(n3349) );
  NOR3_X0P5A_A12TR u3915 ( .A(n3375), .B(rstkptr_[4]), .C(n3377), .Y(n3376) );
  MXT2_X0P5M_A12TR u3916 ( .A(rstkram[307]), .B(wstkw[7]), .S0(n3350), .Y(
        n2077) );
  AND2_X0P5M_A12TR u3917 ( .A(n3378), .B(n3366), .Y(n3350) );
  MXT2_X0P5M_A12TR u3918 ( .A(rstkram[287]), .B(wstkw[7]), .S0(n3351), .Y(
        n2076) );
  AND2_X0P5M_A12TR u3919 ( .A(n3378), .B(n3368), .Y(n3351) );
  MXT2_X0P5M_A12TR u3920 ( .A(rstkram[267]), .B(wstkw[7]), .S0(n3352), .Y(
        n2075) );
  AND2_X0P5M_A12TR u3921 ( .A(n3378), .B(n3369), .Y(n3352) );
  MXT2_X0P5M_A12TR u3922 ( .A(rstkram[247]), .B(wstkw[7]), .S0(n3353), .Y(
        n2074) );
  AND2_X0P5M_A12TR u3923 ( .A(n3378), .B(n3370), .Y(n3353) );
  MXT2_X0P5M_A12TR u3924 ( .A(rstkram[227]), .B(wstkw[7]), .S0(n3354), .Y(
        n2073) );
  AND2_X0P5M_A12TR u3925 ( .A(n3378), .B(n3371), .Y(n3354) );
  MXT2_X0P5M_A12TR u3926 ( .A(rstkram[207]), .B(wstkw[7]), .S0(n3355), .Y(
        n2072) );
  AND2_X0P5M_A12TR u3927 ( .A(n3378), .B(n3372), .Y(n3355) );
  MXT2_X0P5M_A12TR u3928 ( .A(rstkram[187]), .B(wstkw[7]), .S0(n3356), .Y(
        n2071) );
  AND2_X0P5M_A12TR u3929 ( .A(n3378), .B(n3373), .Y(n3356) );
  MXT2_X0P5M_A12TR u3930 ( .A(rstkram[167]), .B(wstkw[7]), .S0(n3357), .Y(
        n2070) );
  AND2_X0P5M_A12TR u3931 ( .A(n3378), .B(n3374), .Y(n3357) );
  NOR3_X0P5A_A12TR u3932 ( .A(n3375), .B(rstkptr_[3]), .C(n3379), .Y(n3378) );
  MXT2_X0P5M_A12TR u3933 ( .A(rstkram[147]), .B(wstkw[7]), .S0(n3358), .Y(
        n2069) );
  AND2_X0P5M_A12TR u3934 ( .A(n3380), .B(n3366), .Y(n3358) );
  NOR3_X0P5A_A12TR u3935 ( .A(rstkptr_[1]), .B(rstkptr_[2]), .C(rstkptr_[0]), 
        .Y(n3366) );
  MXT2_X0P5M_A12TR u3936 ( .A(rstkram[127]), .B(wstkw[7]), .S0(n3359), .Y(
        n2068) );
  AND2_X0P5M_A12TR u3937 ( .A(n3380), .B(n3368), .Y(n3359) );
  NOR3_X0P5A_A12TR u3938 ( .A(rstkptr_[1]), .B(rstkptr_[2]), .C(n3381), .Y(
        n3368) );
  MXT2_X0P5M_A12TR u3939 ( .A(rstkram[107]), .B(wstkw[7]), .S0(n3360), .Y(
        n2067) );
  AND2_X0P5M_A12TR u3940 ( .A(n3380), .B(n3369), .Y(n3360) );
  NOR3_X0P5A_A12TR u3941 ( .A(rstkptr_[0]), .B(rstkptr_[2]), .C(n3382), .Y(
        n3369) );
  MXT2_X0P5M_A12TR u3942 ( .A(rstkram[87]), .B(wstkw[7]), .S0(n3361), .Y(n2066) );
  AND2_X0P5M_A12TR u3943 ( .A(n3380), .B(n3370), .Y(n3361) );
  NOR3_X0P5A_A12TR u3944 ( .A(n3381), .B(rstkptr_[2]), .C(n3382), .Y(n3370) );
  MXT2_X0P5M_A12TR u3945 ( .A(rstkram[67]), .B(wstkw[7]), .S0(n3362), .Y(n2065) );
  AND2_X0P5M_A12TR u3946 ( .A(n3380), .B(n3371), .Y(n3362) );
  NOR3_X0P5A_A12TR u3947 ( .A(rstkptr_[0]), .B(rstkptr_[1]), .C(n3383), .Y(
        n3371) );
  MXT2_X0P5M_A12TR u3948 ( .A(rstkram[47]), .B(wstkw[7]), .S0(n3363), .Y(n2064) );
  AND2_X0P5M_A12TR u3949 ( .A(n3380), .B(n3372), .Y(n3363) );
  NOR3_X0P5A_A12TR u3950 ( .A(n3381), .B(rstkptr_[1]), .C(n3383), .Y(n3372) );
  MXT2_X0P5M_A12TR u3951 ( .A(rstkram[27]), .B(wstkw[7]), .S0(n3364), .Y(n2063) );
  AND2_X0P5M_A12TR u3952 ( .A(n3380), .B(n3373), .Y(n3364) );
  NOR3_X0P5A_A12TR u3953 ( .A(n3382), .B(rstkptr_[0]), .C(n3383), .Y(n3373) );
  MXT2_X0P5M_A12TR u3954 ( .A(rstkram[7]), .B(wstkw[7]), .S0(n3365), .Y(n2062)
         );
  AND2_X0P5M_A12TR u3955 ( .A(n3380), .B(n3374), .Y(n3365) );
  NOR3_X0P5A_A12TR u3956 ( .A(n3382), .B(n3381), .C(n3383), .Y(n3374) );
  NOR3_X0P5A_A12TR u3957 ( .A(n3377), .B(n3375), .C(n3379), .Y(n3380) );
  OAI211_X0P5M_A12TR u3958 ( .A0(n3384), .A1(n3385), .B0(n3386), .C0(n3387), 
        .Y(n2061) );
  AOI22_X0P5M_A12TR u3959 ( .A0(n3388), .A1(rromlat[8]), .B0(reaptr[8]), .B1(
        n3389), .Y(n3387) );
  OAI211_X0P5M_A12TR u3960 ( .A0(n3390), .A1(n3385), .B0(n3386), .C0(n3391), 
        .Y(n2060) );
  AOI22_X0P5M_A12TR u3961 ( .A0(n3388), .A1(rromlat[9]), .B0(reaptr[9]), .B1(
        n3389), .Y(n3391) );
  OAI211_X0P5M_A12TR u3962 ( .A0(n3392), .A1(n3385), .B0(n3386), .C0(n3393), 
        .Y(n2059) );
  AOI22_X0P5M_A12TR u3963 ( .A0(n3388), .A1(rromlat[10]), .B0(reaptr[10]), 
        .B1(n3389), .Y(n3393) );
  OAI211_X0P5M_A12TR u3964 ( .A0(n3394), .A1(n3385), .B0(n3386), .C0(n3395), 
        .Y(n2058) );
  AOI22_X0P5M_A12TR u3965 ( .A0(n3388), .A1(rromlat[11]), .B0(reaptr[11]), 
        .B1(n3389), .Y(n3395) );
  NOR2_X0P5A_A12TR u3966 ( .A(n3396), .B(rmxbsr[1]), .Y(n3388) );
  NAND2B_X0P5M_A12TR u3967 ( .AN(n3396), .B(rmxbsr[1]), .Y(n3385) );
  OAI221_X0P5M_A12TR u3968 ( .A0(n3397), .A1(n3396), .B0(n3398), .B1(n3399), 
        .C0(n3386), .Y(n2057) );
  OAI221_X0P5M_A12TR u3969 ( .A0(n3396), .A1(n3400), .B0(n3398), .B1(n3401), 
        .C0(n3386), .Y(n2056) );
  OAI221_X0P5M_A12TR u3970 ( .A0(n3402), .A1(n3396), .B0(n3398), .B1(n3403), 
        .C0(n3386), .Y(n2055) );
  OAI221_X0P5M_A12TR u3971 ( .A0(n3404), .A1(n3396), .B0(n3398), .B1(n3405), 
        .C0(n3386), .Y(n2054) );
  NAND3_X0P5A_A12TR u3972 ( .A(rromlat[7]), .B(n3406), .C(n3398), .Y(n3386) );
  NAND2_X0P5A_A12TR u3973 ( .A(rmxbsr[0]), .B(n3398), .Y(n3396) );
  OAI221_X0P5M_A12TR u3974 ( .A0(n3192), .A1(n3183), .B0(n3184), .B1(n3407), 
        .C0(n3408), .Y(n2053) );
  AOI222_X0P5M_A12TR u3975 ( .A0(wfsrdec2[0]), .A1(n3187), .B0(rfsr2l[0]), 
        .B1(n3188), .C0(n3189), .C1(dwb_dat_o[0]), .Y(n3408) );
  INV_X0P5B_A12TR u3976 ( .A(wfsrinc2[0]), .Y(n3407) );
  OAI221_X0P5M_A12TR u3977 ( .A0(n3083), .A1(n3183), .B0(n3184), .B1(n3409), 
        .C0(n3410), .Y(n2052) );
  AOI222_X0P5M_A12TR u3978 ( .A0(wfsrdec2[1]), .A1(n3187), .B0(rfsr2l[1]), 
        .B1(n3188), .C0(dwb_dat_o[1]), .C1(n3189), .Y(n3410) );
  INV_X0P5B_A12TR u3979 ( .A(wfsrinc2[1]), .Y(n3409) );
  OAI221_X0P5M_A12TR u3980 ( .A0(n3084), .A1(n3183), .B0(n3184), .B1(n3411), 
        .C0(n3412), .Y(n2051) );
  AOI222_X0P5M_A12TR u3981 ( .A0(wfsrdec2[2]), .A1(n3187), .B0(rfsr2l[2]), 
        .B1(n3188), .C0(n3189), .C1(dwb_dat_o[2]), .Y(n3412) );
  INV_X0P5B_A12TR u3982 ( .A(wfsrinc2[2]), .Y(n3411) );
  OAI221_X0P5M_A12TR u3983 ( .A0(n3197), .A1(n3183), .B0(n3184), .B1(n3413), 
        .C0(n3414), .Y(n2050) );
  AOI222_X0P5M_A12TR u3984 ( .A0(wfsrdec2[3]), .A1(n3187), .B0(rfsr2l[3]), 
        .B1(n3188), .C0(n3189), .C1(dwb_dat_o[3]), .Y(n3414) );
  INV_X0P5B_A12TR u3985 ( .A(wfsrinc2[3]), .Y(n3413) );
  OAI221_X0P5M_A12TR u3986 ( .A0(n3199), .A1(n3183), .B0(n3184), .B1(n3415), 
        .C0(n3416), .Y(n2049) );
  AOI222_X0P5M_A12TR u3987 ( .A0(wfsrdec2[4]), .A1(n3187), .B0(rfsr2l[4]), 
        .B1(n3188), .C0(n3189), .C1(dwb_dat_o[4]), .Y(n3416) );
  INV_X0P5B_A12TR u3988 ( .A(wfsrinc2[4]), .Y(n3415) );
  OAI221_X0P5M_A12TR u3989 ( .A0(n3201), .A1(n3183), .B0(n3184), .B1(n3417), 
        .C0(n3418), .Y(n2048) );
  AOI222_X0P5M_A12TR u3990 ( .A0(wfsrdec2[5]), .A1(n3187), .B0(rfsr2l[5]), 
        .B1(n3188), .C0(dwb_dat_o[5]), .C1(n3189), .Y(n3418) );
  INV_X0P5B_A12TR u3991 ( .A(wfsrinc2[5]), .Y(n3417) );
  OAI221_X0P5M_A12TR u3992 ( .A0(n3088), .A1(n3183), .B0(n3184), .B1(n3419), 
        .C0(n3420), .Y(n2047) );
  AOI222_X0P5M_A12TR u3993 ( .A0(wfsrdec2[6]), .A1(n3187), .B0(rfsr2l[6]), 
        .B1(n3188), .C0(dwb_dat_o[6]), .C1(n3189), .Y(n3420) );
  AND3_X0P5M_A12TR u3994 ( .A(n3421), .B(n3122), .C(n3422), .Y(n3189) );
  OAI211_X0P5M_A12TR u3995 ( .A0(n3122), .A1(n3423), .B0(n3424), .C0(n3421), 
        .Y(n3188) );
  INV_X0P5B_A12TR u3996 ( .A(wfsrinc2[6]), .Y(n3419) );
  OAI221_X0P5M_A12TR u3997 ( .A0(n3192), .A1(n3425), .B0(n3426), .B1(n3427), 
        .C0(n3428), .Y(n2046) );
  AOI222_X0P5M_A12TR u3998 ( .A0(wfsrdec0[0]), .A1(n3429), .B0(rfsr0l[0]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[0]), .Y(n3428) );
  INV_X0P5B_A12TR u3999 ( .A(wfsrinc0[0]), .Y(n3427) );
  OAI221_X0P5M_A12TR u4000 ( .A0(n3083), .A1(n3425), .B0(n3426), .B1(n3432), 
        .C0(n3433), .Y(n2045) );
  AOI222_X0P5M_A12TR u4001 ( .A0(wfsrdec0[1]), .A1(n3429), .B0(rfsr0l[1]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[1]), .Y(n3433) );
  INV_X0P5B_A12TR u4002 ( .A(wfsrinc0[1]), .Y(n3432) );
  OAI221_X0P5M_A12TR u4003 ( .A0(n3084), .A1(n3425), .B0(n3426), .B1(n3434), 
        .C0(n3435), .Y(n2044) );
  AOI222_X0P5M_A12TR u4004 ( .A0(wfsrdec0[2]), .A1(n3429), .B0(rfsr0l[2]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[2]), .Y(n3435) );
  INV_X0P5B_A12TR u4005 ( .A(wfsrinc0[2]), .Y(n3434) );
  OAI221_X0P5M_A12TR u4006 ( .A0(n3197), .A1(n3425), .B0(n3426), .B1(n3436), 
        .C0(n3437), .Y(n2043) );
  AOI222_X0P5M_A12TR u4007 ( .A0(wfsrdec0[3]), .A1(n3429), .B0(rfsr0l[3]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[3]), .Y(n3437) );
  INV_X0P5B_A12TR u4008 ( .A(wfsrinc0[3]), .Y(n3436) );
  OAI221_X0P5M_A12TR u4009 ( .A0(n3199), .A1(n3425), .B0(n3426), .B1(n3438), 
        .C0(n3439), .Y(n2042) );
  AOI222_X0P5M_A12TR u4010 ( .A0(wfsrdec0[4]), .A1(n3429), .B0(rfsr0l[4]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[4]), .Y(n3439) );
  INV_X0P5B_A12TR u4011 ( .A(wfsrinc0[4]), .Y(n3438) );
  OAI221_X0P5M_A12TR u4012 ( .A0(n3201), .A1(n3425), .B0(n3426), .B1(n3440), 
        .C0(n3441), .Y(n2041) );
  AOI222_X0P5M_A12TR u4013 ( .A0(wfsrdec0[5]), .A1(n3429), .B0(rfsr0l[5]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[5]), .Y(n3441) );
  INV_X0P5B_A12TR u4014 ( .A(wfsrinc0[5]), .Y(n3440) );
  OAI221_X0P5M_A12TR u4015 ( .A0(n3088), .A1(n3425), .B0(n3426), .B1(n3442), 
        .C0(n3443), .Y(n2040) );
  AOI222_X0P5M_A12TR u4016 ( .A0(wfsrdec0[6]), .A1(n3429), .B0(rfsr0l[6]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[6]), .Y(n3443) );
  INV_X0P5B_A12TR u4017 ( .A(wfsrinc0[6]), .Y(n3442) );
  OAI221_X0P5M_A12TR u4018 ( .A0(n3089), .A1(n3425), .B0(n3426), .B1(n3444), 
        .C0(n3445), .Y(n2039) );
  AOI222_X0P5M_A12TR u4019 ( .A0(wfsrdec0[7]), .A1(n3429), .B0(rfsr0l[7]), 
        .B1(n3430), .C0(n3431), .C1(dwb_dat_o[7]), .Y(n3445) );
  AND3_X0P5M_A12TR u4020 ( .A(n3422), .B(n3123), .C(n3446), .Y(n3431) );
  OAI211_X0P5M_A12TR u4021 ( .A0(n3123), .A1(n3423), .B0(n3424), .C0(n3446), 
        .Y(n3430) );
  INV_X0P5B_A12TR u4022 ( .A(wfsrinc0[7]), .Y(n3444) );
  OAI221_X0P5M_A12TR u4023 ( .A0(n3447), .A1(n3255), .B0(n3067), .B1(n3448), 
        .C0(n3449), .Y(n2038) );
  AOI222_X0P5M_A12TR u4024 ( .A0(wfsrinc0[8]), .A1(n3450), .B0(wfsrdec0[8]), 
        .B1(n3429), .C0(n3451), .C1(rireg[0]), .Y(n3449) );
  INV_X0P5B_A12TR u4025 ( .A(rfsr0h[0]), .Y(n3255) );
  OAI221_X0P5M_A12TR u4026 ( .A0(n3447), .A1(n3452), .B0(n3453), .B1(n3448), 
        .C0(n3454), .Y(n2037) );
  AOI222_X0P5M_A12TR u4027 ( .A0(wfsrinc0[9]), .A1(n3450), .B0(wfsrdec0[9]), 
        .B1(n3429), .C0(n3451), .C1(rireg[1]), .Y(n3454) );
  INV_X0P5B_A12TR u4028 ( .A(rfsr0h[1]), .Y(n3452) );
  OAI221_X0P5M_A12TR u4029 ( .A0(n3447), .A1(n3455), .B0(n3158), .B1(n3448), 
        .C0(n3456), .Y(n2036) );
  AOI222_X0P5M_A12TR u4030 ( .A0(wfsrinc0[10]), .A1(n3450), .B0(wfsrdec0[10]), 
        .B1(n3429), .C0(n3451), .C1(rireg[2]), .Y(n3456) );
  INV_X0P5B_A12TR u4031 ( .A(rfsr0h[2]), .Y(n3455) );
  OAI221_X0P5M_A12TR u4032 ( .A0(n3447), .A1(n3457), .B0(n3458), .B1(n3448), 
        .C0(n3459), .Y(n2035) );
  AOI222_X0P5M_A12TR u4033 ( .A0(wfsrinc0[11]), .A1(n3450), .B0(wfsrdec0[11]), 
        .B1(n3429), .C0(n3451), .C1(rireg[3]), .Y(n3459) );
  INV_X0P5B_A12TR u4034 ( .A(n3425), .Y(n3451) );
  NAND2_X0P5A_A12TR u4035 ( .A(n3446), .B(n3460), .Y(n3425) );
  AND2_X0P5M_A12TR u4036 ( .A(n3461), .B(n3462), .Y(n3429) );
  INV_X0P5B_A12TR u4037 ( .A(n3426), .Y(n3450) );
  AOI22_X0P5M_A12TR u4038 ( .A0(n3143), .A1(n3446), .B0(n3463), .B1(n3461), 
        .Y(n3426) );
  NOR2_X0P5A_A12TR u4039 ( .A(n3464), .B(n3238), .Y(n3461) );
  INV_X0P5B_A12TR u4040 ( .A(rfsr0h[3]), .Y(n3457) );
  OAI22_X0P5M_A12TR u4041 ( .A0(n3148), .A1(n3448), .B0(n3447), .B1(n3465), 
        .Y(n2034) );
  INV_X0P5B_A12TR u4042 ( .A(rfsr0h[4]), .Y(n3465) );
  OAI22_X0P5M_A12TR u4043 ( .A0(n3466), .A1(n3448), .B0(n3447), .B1(n3467), 
        .Y(n2033) );
  INV_X0P5B_A12TR u4044 ( .A(rfsr0h[5]), .Y(n3467) );
  OAI22_X0P5M_A12TR u4045 ( .A0(n3468), .A1(n3448), .B0(n3447), .B1(n3469), 
        .Y(n2032) );
  INV_X0P5B_A12TR u4046 ( .A(rfsr0h[6]), .Y(n3469) );
  OAI22_X0P5M_A12TR u4047 ( .A0(n3470), .A1(n3448), .B0(n3447), .B1(n3471), 
        .Y(n2031) );
  INV_X0P5B_A12TR u4048 ( .A(rfsr0h[7]), .Y(n3471) );
  AOI211_X0P5M_A12TR u4049 ( .A0(n3254), .A1(n3472), .B0(n3473), .C0(n3464), 
        .Y(n3447) );
  INV_X0P5B_A12TR u4050 ( .A(n3446), .Y(n3464) );
  NAND3_X0P5A_A12TR u4051 ( .A(n3422), .B(n3127), .C(n3446), .Y(n3448) );
  AOI21_X0P5M_A12TR u4052 ( .A0(n3474), .A1(n3475), .B0(n3476), .Y(n3446) );
  AOI31_X0P5M_A12TR u4053 ( .A0(n3477), .A1(n3233), .A2(n3232), .B0(n3478), 
        .Y(n3475) );
  AND3_X0P5M_A12TR u4054 ( .A(n3247), .B(n3479), .C(n3480), .Y(n3478) );
  MXIT2_X0P5M_A12TR u4055 ( .A(n3481), .B(n3482), .S0(n3483), .Y(n3480) );
  AOI31_X0P5M_A12TR u4056 ( .A0(n3484), .A1(n3483), .A2(n3143), .B0(n3472), 
        .Y(n3474) );
  OAI221_X0P5M_A12TR u4057 ( .A0(n3192), .A1(n3485), .B0(n3486), .B1(n3487), 
        .C0(n3488), .Y(n2030) );
  AOI222_X0P5M_A12TR u4058 ( .A0(wfsrdec1[0]), .A1(n3489), .B0(rfsr1l[0]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[0]), .Y(n3488) );
  INV_X0P5B_A12TR u4059 ( .A(wfsrinc1[0]), .Y(n3487) );
  OAI221_X0P5M_A12TR u4060 ( .A0(n3083), .A1(n3485), .B0(n3486), .B1(n3492), 
        .C0(n3493), .Y(n2029) );
  AOI222_X0P5M_A12TR u4061 ( .A0(wfsrdec1[1]), .A1(n3489), .B0(rfsr1l[1]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[1]), .Y(n3493) );
  INV_X0P5B_A12TR u4062 ( .A(wfsrinc1[1]), .Y(n3492) );
  OAI221_X0P5M_A12TR u4063 ( .A0(n3084), .A1(n3485), .B0(n3486), .B1(n3494), 
        .C0(n3495), .Y(n2028) );
  AOI222_X0P5M_A12TR u4064 ( .A0(wfsrdec1[2]), .A1(n3489), .B0(rfsr1l[2]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[2]), .Y(n3495) );
  INV_X0P5B_A12TR u4065 ( .A(wfsrinc1[2]), .Y(n3494) );
  OAI221_X0P5M_A12TR u4066 ( .A0(n3197), .A1(n3485), .B0(n3486), .B1(n3496), 
        .C0(n3497), .Y(n2027) );
  AOI222_X0P5M_A12TR u4067 ( .A0(wfsrdec1[3]), .A1(n3489), .B0(rfsr1l[3]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[3]), .Y(n3497) );
  INV_X0P5B_A12TR u4068 ( .A(wfsrinc1[3]), .Y(n3496) );
  OAI221_X0P5M_A12TR u4069 ( .A0(n3199), .A1(n3485), .B0(n3486), .B1(n3498), 
        .C0(n3499), .Y(n2026) );
  AOI222_X0P5M_A12TR u4070 ( .A0(wfsrdec1[4]), .A1(n3489), .B0(rfsr1l[4]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[4]), .Y(n3499) );
  INV_X0P5B_A12TR u4071 ( .A(wfsrinc1[4]), .Y(n3498) );
  OAI221_X0P5M_A12TR u4072 ( .A0(n3201), .A1(n3485), .B0(n3486), .B1(n3500), 
        .C0(n3501), .Y(n2025) );
  AOI222_X0P5M_A12TR u4073 ( .A0(wfsrdec1[5]), .A1(n3489), .B0(rfsr1l[5]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[5]), .Y(n3501) );
  INV_X0P5B_A12TR u4074 ( .A(wfsrinc1[5]), .Y(n3500) );
  OAI221_X0P5M_A12TR u4075 ( .A0(n3088), .A1(n3485), .B0(n3486), .B1(n3502), 
        .C0(n3503), .Y(n2024) );
  AOI222_X0P5M_A12TR u4076 ( .A0(wfsrdec1[6]), .A1(n3489), .B0(rfsr1l[6]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[6]), .Y(n3503) );
  INV_X0P5B_A12TR u4077 ( .A(wfsrinc1[6]), .Y(n3502) );
  OAI221_X0P5M_A12TR u4078 ( .A0(n3089), .A1(n3485), .B0(n3486), .B1(n3504), 
        .C0(n3505), .Y(n2023) );
  AOI222_X0P5M_A12TR u4079 ( .A0(wfsrdec1[7]), .A1(n3489), .B0(rfsr1l[7]), 
        .B1(n3490), .C0(n3491), .C1(dwb_dat_o[7]), .Y(n3505) );
  AND3_X0P5M_A12TR u4080 ( .A(n3121), .B(n3506), .C(n3422), .Y(n3491) );
  OAI211_X0P5M_A12TR u4081 ( .A0(n3121), .A1(n3423), .B0(n3506), .C0(n3424), 
        .Y(n3490) );
  INV_X0P5B_A12TR u4082 ( .A(wfsrinc1[7]), .Y(n3504) );
  OAI221_X0P5M_A12TR u4083 ( .A0(n3507), .A1(n3508), .B0(n3067), .B1(n3509), 
        .C0(n3510), .Y(n2022) );
  AOI222_X0P5M_A12TR u4084 ( .A0(wfsrinc1[8]), .A1(n3511), .B0(wfsrdec1[8]), 
        .B1(n3489), .C0(n3512), .C1(rireg[0]), .Y(n3510) );
  INV_X0P5B_A12TR u4085 ( .A(rfsr1h[0]), .Y(n3508) );
  OAI221_X0P5M_A12TR u4086 ( .A0(n3507), .A1(n3513), .B0(n3453), .B1(n3509), 
        .C0(n3514), .Y(n2021) );
  AOI222_X0P5M_A12TR u4087 ( .A0(wfsrinc1[9]), .A1(n3511), .B0(wfsrdec1[9]), 
        .B1(n3489), .C0(n3512), .C1(rireg[1]), .Y(n3514) );
  INV_X0P5B_A12TR u4088 ( .A(rfsr1h[1]), .Y(n3513) );
  OAI221_X0P5M_A12TR u4089 ( .A0(n3507), .A1(n3515), .B0(n3158), .B1(n3509), 
        .C0(n3516), .Y(n2020) );
  AOI222_X0P5M_A12TR u4090 ( .A0(wfsrinc1[10]), .A1(n3511), .B0(wfsrdec1[10]), 
        .B1(n3489), .C0(n3512), .C1(rireg[2]), .Y(n3516) );
  INV_X0P5B_A12TR u4091 ( .A(rfsr1h[2]), .Y(n3515) );
  OAI221_X0P5M_A12TR u4092 ( .A0(n3507), .A1(n3517), .B0(n3458), .B1(n3509), 
        .C0(n3518), .Y(n2019) );
  AOI222_X0P5M_A12TR u4093 ( .A0(wfsrinc1[11]), .A1(n3511), .B0(wfsrdec1[11]), 
        .B1(n3489), .C0(n3512), .C1(rireg[3]), .Y(n3518) );
  INV_X0P5B_A12TR u4094 ( .A(n3485), .Y(n3512) );
  NAND2_X0P5A_A12TR u4095 ( .A(n3460), .B(n3506), .Y(n3485) );
  AND3_X0P5M_A12TR u4096 ( .A(n3463), .B(n3506), .C(n3519), .Y(n3489) );
  INV_X0P5B_A12TR u4097 ( .A(n3486), .Y(n3511) );
  OAI21_X0P5M_A12TR u4098 ( .A0(n3143), .A1(n3520), .B0(n3506), .Y(n3486) );
  INV_X0P5B_A12TR u4099 ( .A(rfsr1h[3]), .Y(n3517) );
  OAI22_X0P5M_A12TR u4100 ( .A0(n3148), .A1(n3509), .B0(n3507), .B1(n3521), 
        .Y(n2018) );
  INV_X0P5B_A12TR u4101 ( .A(rfsr1h[4]), .Y(n3521) );
  OAI22_X0P5M_A12TR u4102 ( .A0(n3466), .A1(n3509), .B0(n3507), .B1(n3522), 
        .Y(n2017) );
  INV_X0P5B_A12TR u4103 ( .A(rfsr1h[5]), .Y(n3522) );
  OAI22_X0P5M_A12TR u4104 ( .A0(n3468), .A1(n3509), .B0(n3507), .B1(n3523), 
        .Y(n2016) );
  INV_X0P5B_A12TR u4105 ( .A(rfsr1h[6]), .Y(n3523) );
  OAI22_X0P5M_A12TR u4106 ( .A0(n3470), .A1(n3509), .B0(n3507), .B1(n3524), 
        .Y(n2015) );
  INV_X0P5B_A12TR u4107 ( .A(rfsr1h[7]), .Y(n3524) );
  OA211_X0P5M_A12TR u4108 ( .A0(n3117), .A1(n3423), .B0(n3506), .C0(n3424), 
        .Y(n3507) );
  NAND3_X0P5A_A12TR u4109 ( .A(n3117), .B(n3506), .C(n3422), .Y(n3509) );
  AO21A1AI2_X0P5M_A12TR u4110 ( .A0(n3525), .A1(n3526), .B0(n3476), .C0(n3527), 
        .Y(n3506) );
  NOR2_X0P5A_A12TR u4111 ( .A(n3472), .B(n3520), .Y(n3526) );
  AND3_X0P5M_A12TR u4112 ( .A(rmxfsr[0]), .B(n3528), .C(n3519), .Y(n3520) );
  AOI32_X0P5M_A12TR u4113 ( .A0(n3477), .A1(n3233), .A2(rireg[4]), .B0(n3519), 
        .B1(n3463), .Y(n3525) );
  NOR3_X0P5A_A12TR u4114 ( .A(n3238), .B(rmxfsr[2]), .C(n3479), .Y(n3519) );
  INV_X0P5B_A12TR u4115 ( .A(n3529), .Y(n3477) );
  OAI221_X0P5M_A12TR u4116 ( .A0(n3530), .A1(n3531), .B0(n3067), .B1(n3532), 
        .C0(n3533), .Y(n2014) );
  AOI222_X0P5M_A12TR u4117 ( .A0(wfsrinc2[8]), .A1(n3534), .B0(wfsrdec2[8]), 
        .B1(n3187), .C0(rireg[0]), .C1(n3535), .Y(n3533) );
  INV_X0P5B_A12TR u4118 ( .A(rfsr2h[0]), .Y(n3531) );
  OAI221_X0P5M_A12TR u4119 ( .A0(n3530), .A1(n3536), .B0(n3453), .B1(n3532), 
        .C0(n3537), .Y(n2013) );
  AOI222_X0P5M_A12TR u4120 ( .A0(wfsrinc2[9]), .A1(n3534), .B0(wfsrdec2[9]), 
        .B1(n3187), .C0(rireg[1]), .C1(n3535), .Y(n3537) );
  INV_X0P5B_A12TR u4121 ( .A(rfsr2h[1]), .Y(n3536) );
  OAI221_X0P5M_A12TR u4122 ( .A0(n3530), .A1(n3538), .B0(n3158), .B1(n3532), 
        .C0(n3539), .Y(n2012) );
  AOI222_X0P5M_A12TR u4123 ( .A0(wfsrinc2[10]), .A1(n3534), .B0(wfsrdec2[10]), 
        .B1(n3187), .C0(rireg[2]), .C1(n3535), .Y(n3539) );
  INV_X0P5B_A12TR u4124 ( .A(rfsr2h[2]), .Y(n3538) );
  OAI221_X0P5M_A12TR u4125 ( .A0(n3530), .A1(n3540), .B0(n3458), .B1(n3532), 
        .C0(n3541), .Y(n2011) );
  AOI222_X0P5M_A12TR u4126 ( .A0(wfsrinc2[11]), .A1(n3534), .B0(wfsrdec2[11]), 
        .B1(n3187), .C0(rireg[3]), .C1(n3535), .Y(n3541) );
  INV_X0P5B_A12TR u4127 ( .A(n3183), .Y(n3535) );
  NAND2_X0P5A_A12TR u4128 ( .A(n3421), .B(n3460), .Y(n3183) );
  AND2_X0P5M_A12TR u4129 ( .A(n3542), .B(rmxfsr[0]), .Y(n3187) );
  INV_X0P5B_A12TR u4130 ( .A(n3184), .Y(n3534) );
  AOI22_X0P5M_A12TR u4131 ( .A0(n3143), .A1(n3421), .B0(n3543), .B1(n3542), 
        .Y(n3184) );
  NOR2_X0P5A_A12TR u4132 ( .A(n3544), .B(n3238), .Y(n3542) );
  INV_X0P5B_A12TR u4133 ( .A(rfsr2h[3]), .Y(n3540) );
  OAI22_X0P5M_A12TR u4134 ( .A0(n3148), .A1(n3532), .B0(n3530), .B1(n3545), 
        .Y(n2010) );
  INV_X0P5B_A12TR u4135 ( .A(rfsr2h[4]), .Y(n3545) );
  OAI22_X0P5M_A12TR u4136 ( .A0(n3466), .A1(n3532), .B0(n1942), .B1(n3530), 
        .Y(n2009) );
  OAI22_X0P5M_A12TR u4137 ( .A0(n3468), .A1(n3532), .B0(n1941), .B1(n3530), 
        .Y(n2008) );
  OAI22_X0P5M_A12TR u4138 ( .A0(n3470), .A1(n3532), .B0(n1940), .B1(n3530), 
        .Y(n2007) );
  AOI211_X0P5M_A12TR u4139 ( .A0(n3546), .A1(n3472), .B0(n3473), .C0(n3544), 
        .Y(n3530) );
  NAND3_X0P5A_A12TR u4140 ( .A(n3421), .B(n3124), .C(n3422), .Y(n3532) );
  INV_X0P5B_A12TR u4141 ( .A(n3544), .Y(n3421) );
  OAI21_X0P5M_A12TR u4142 ( .A0(n3547), .A1(n3548), .B0(n3242), .Y(n3544) );
  OAI31_X0P5M_A12TR u4143 ( .A0(n3233), .A1(rireg[4]), .A2(n3529), .B0(n3423), 
        .Y(n3548) );
  NAND4_X0P5A_A12TR u4144 ( .A(n3460), .B(n3549), .C(n3550), .D(n3551), .Y(
        n3529) );
  MXIT2_X0P5M_A12TR u4145 ( .A(n3552), .B(n3553), .S0(n3481), .Y(n3547) );
  NAND3_X0P5A_A12TR u4146 ( .A(n3247), .B(n3482), .C(n3554), .Y(n3553) );
  NAND2_X0P5A_A12TR u4147 ( .A(n3554), .B(n3143), .Y(n3552) );
  AO22_X0P5M_A12TR u4148 ( .A0(n239), .A1(n3190), .B0(rwdt[15]), .B1(n3191), 
        .Y(n2006) );
  AO22_X0P5M_A12TR u4149 ( .A0(n238), .A1(n3190), .B0(rwdt[14]), .B1(n3191), 
        .Y(n2005) );
  AO22_X0P5M_A12TR u4150 ( .A0(n237), .A1(n3190), .B0(rwdt[13]), .B1(n3191), 
        .Y(n2004) );
  AO22_X0P5M_A12TR u4151 ( .A0(n236), .A1(n3190), .B0(rwdt[12]), .B1(n3191), 
        .Y(n2003) );
  AO22_X0P5M_A12TR u4152 ( .A0(n235), .A1(n3190), .B0(rwdt[11]), .B1(n3191), 
        .Y(n2002) );
  AO22_X0P5M_A12TR u4153 ( .A0(n234), .A1(n3190), .B0(rwdt[10]), .B1(n3191), 
        .Y(n2001) );
  AO22_X0P5M_A12TR u4154 ( .A0(n233), .A1(n3190), .B0(rwdt[9]), .B1(n3191), 
        .Y(n2000) );
  AO22_X0P5M_A12TR u4155 ( .A0(n232), .A1(n3190), .B0(rwdt[8]), .B1(n3191), 
        .Y(n1999) );
  AO22_X0P5M_A12TR u4156 ( .A0(n231), .A1(n3190), .B0(rwdt[7]), .B1(n3191), 
        .Y(n1998) );
  AO22_X0P5M_A12TR u4157 ( .A0(n230), .A1(n3190), .B0(rwdt[6]), .B1(n3191), 
        .Y(n1997) );
  AO22_X0P5M_A12TR u4158 ( .A0(n229), .A1(n3190), .B0(rwdt[5]), .B1(n3191), 
        .Y(n1996) );
  AO22_X0P5M_A12TR u4159 ( .A0(n228), .A1(n3190), .B0(rwdt[4]), .B1(n3191), 
        .Y(n1995) );
  AO22_X0P5M_A12TR u4160 ( .A0(n227), .A1(n3190), .B0(rwdt[3]), .B1(n3191), 
        .Y(n1994) );
  AO22_X0P5M_A12TR u4161 ( .A0(n226), .A1(n3190), .B0(rwdt[2]), .B1(n3191), 
        .Y(n1993) );
  AO22_X0P5M_A12TR u4162 ( .A0(n225), .A1(n3190), .B0(rwdt[1]), .B1(n3191), 
        .Y(n1992) );
  AO22_X0P5M_A12TR u4163 ( .A0(n224), .A1(n3190), .B0(rwdt[0]), .B1(n3191), 
        .Y(n1991) );
  NOR3_X0P5A_A12TR u4164 ( .A(rclrwdt), .B(rsleep), .C(n3190), .Y(n3191) );
  NOR3_X0P5A_A12TR u4165 ( .A(rclrwdt), .B(rsleep), .C(n3555), .Y(n3190) );
  OAI221_X0P5M_A12TR u4166 ( .A0(n3067), .A1(n3556), .B0(n3557), .B1(n3558), 
        .C0(n3559), .Y(n1990) );
  AOI22_X0P5M_A12TR u4167 ( .A0(wtbldec[0]), .A1(n3560), .B0(wtblinc[0]), .B1(
        n3561), .Y(n3559) );
  OAI222_X0P5M_A12TR u4168 ( .A0(n3193), .A1(n3562), .B0(n3206), .B1(n3563), 
        .C0(n3564), .C1(n3565), .Y(n1989) );
  INV_X0P5B_A12TR u4169 ( .A(iwb_dat_i[8]), .Y(n3206) );
  INV_X0P5B_A12TR u4170 ( .A(iwb_dat_i[0]), .Y(n3193) );
  OAI222_X0P5M_A12TR u4171 ( .A0(n3195), .A1(n3562), .B0(n3208), .B1(n3563), 
        .C0(n3564), .C1(n3566), .Y(n1988) );
  INV_X0P5B_A12TR u4172 ( .A(iwb_dat_i[9]), .Y(n3208) );
  INV_X0P5B_A12TR u4173 ( .A(iwb_dat_i[1]), .Y(n3195) );
  OAI222_X0P5M_A12TR u4174 ( .A0(n3196), .A1(n3562), .B0(n3210), .B1(n3563), 
        .C0(n3564), .C1(n3567), .Y(n1987) );
  INV_X0P5B_A12TR u4175 ( .A(iwb_dat_i[10]), .Y(n3210) );
  INV_X0P5B_A12TR u4176 ( .A(iwb_dat_i[2]), .Y(n3196) );
  OAI222_X0P5M_A12TR u4177 ( .A0(n3198), .A1(n3562), .B0(n3212), .B1(n3563), 
        .C0(n3564), .C1(n3568), .Y(n1986) );
  INV_X0P5B_A12TR u4178 ( .A(iwb_dat_i[11]), .Y(n3212) );
  INV_X0P5B_A12TR u4179 ( .A(iwb_dat_i[3]), .Y(n3198) );
  OAI222_X0P5M_A12TR u4180 ( .A0(n3200), .A1(n3562), .B0(n3214), .B1(n3563), 
        .C0(n3564), .C1(n3569), .Y(n1985) );
  INV_X0P5B_A12TR u4181 ( .A(iwb_dat_i[12]), .Y(n3214) );
  INV_X0P5B_A12TR u4182 ( .A(iwb_dat_i[4]), .Y(n3200) );
  OAI222_X0P5M_A12TR u4183 ( .A0(n3202), .A1(n3562), .B0(n3216), .B1(n3563), 
        .C0(n3564), .C1(n3570), .Y(n1984) );
  INV_X0P5B_A12TR u4184 ( .A(iwb_dat_i[13]), .Y(n3216) );
  INV_X0P5B_A12TR u4185 ( .A(iwb_dat_i[5]), .Y(n3202) );
  OAI222_X0P5M_A12TR u4186 ( .A0(n3203), .A1(n3562), .B0(n3218), .B1(n3563), 
        .C0(n3564), .C1(n3571), .Y(n1983) );
  INV_X0P5B_A12TR u4187 ( .A(iwb_dat_i[14]), .Y(n3218) );
  INV_X0P5B_A12TR u4188 ( .A(iwb_dat_i[6]), .Y(n3203) );
  OAI222_X0P5M_A12TR u4189 ( .A0(n3204), .A1(n3562), .B0(n3220), .B1(n3563), 
        .C0(n3564), .C1(n3572), .Y(n1982) );
  NAND2_X0P5A_A12TR u4190 ( .A(n3564), .B(n3558), .Y(n3563) );
  INV_X0P5B_A12TR u4191 ( .A(iwb_dat_i[15]), .Y(n3220) );
  NAND2_X0P5A_A12TR u4192 ( .A(n3564), .B(wtblat[0]), .Y(n3562) );
  NOR2_X0P5A_A12TR u4193 ( .A(n3238), .B(n3221), .Y(n3564) );
  INV_X0P5B_A12TR u4194 ( .A(iwb_dat_i[7]), .Y(n3204) );
  OAI221_X0P5M_A12TR u4195 ( .A0(n3453), .A1(n3556), .B0(n3557), .B1(n3573), 
        .C0(n3574), .Y(n1981) );
  AOI22_X0P5M_A12TR u4196 ( .A0(wtbldec[1]), .A1(n3560), .B0(wtblinc[1]), .B1(
        n3561), .Y(n3574) );
  OAI221_X0P5M_A12TR u4197 ( .A0(n3158), .A1(n3556), .B0(n3557), .B1(n3575), 
        .C0(n3576), .Y(n1980) );
  AOI22_X0P5M_A12TR u4198 ( .A0(wtbldec[2]), .A1(n3560), .B0(wtblinc[2]), .B1(
        n3561), .Y(n3576) );
  OAI221_X0P5M_A12TR u4199 ( .A0(n3458), .A1(n3556), .B0(n3557), .B1(n3577), 
        .C0(n3578), .Y(n1979) );
  AOI22_X0P5M_A12TR u4200 ( .A0(wtbldec[3]), .A1(n3560), .B0(wtblinc[3]), .B1(
        n3561), .Y(n3578) );
  OAI221_X0P5M_A12TR u4201 ( .A0(n3148), .A1(n3556), .B0(n3557), .B1(n3579), 
        .C0(n3580), .Y(n1978) );
  AOI22_X0P5M_A12TR u4202 ( .A0(wtbldec[4]), .A1(n3560), .B0(wtblinc[4]), .B1(
        n3561), .Y(n3580) );
  INV_X0P5B_A12TR u4203 ( .A(wtblat[4]), .Y(n3579) );
  OAI221_X0P5M_A12TR u4204 ( .A0(n3466), .A1(n3556), .B0(n3557), .B1(n3581), 
        .C0(n3582), .Y(n1977) );
  AOI22_X0P5M_A12TR u4205 ( .A0(wtbldec[5]), .A1(n3560), .B0(wtblinc[5]), .B1(
        n3561), .Y(n3582) );
  OAI221_X0P5M_A12TR u4206 ( .A0(n3468), .A1(n3556), .B0(n3557), .B1(n3583), 
        .C0(n3584), .Y(n1976) );
  AOI22_X0P5M_A12TR u4207 ( .A0(wtbldec[6]), .A1(n3560), .B0(wtblinc[6]), .B1(
        n3561), .Y(n3584) );
  OAI221_X0P5M_A12TR u4208 ( .A0(n3470), .A1(n3556), .B0(n3557), .B1(n3585), 
        .C0(n3586), .Y(n1975) );
  AOI22_X0P5M_A12TR u4209 ( .A0(wtbldec[7]), .A1(n3560), .B0(wtblinc[7]), .B1(
        n3561), .Y(n3586) );
  AOI211_X0P5M_A12TR u4210 ( .A0(n3587), .A1(qfsm[0]), .B0(n3248), .C0(n3588), 
        .Y(n3557) );
  NAND3_X0P5A_A12TR u4211 ( .A(n3119), .B(n3240), .C(n3589), .Y(n3556) );
  OAI221_X0P5M_A12TR u4212 ( .A0(n3067), .A1(n3590), .B0(n3591), .B1(n3592), 
        .C0(n3593), .Y(n1974) );
  AOI22_X0P5M_A12TR u4213 ( .A0(wtbldec[16]), .A1(n3560), .B0(wtblinc[16]), 
        .B1(n3561), .Y(n3593) );
  OAI221_X0P5M_A12TR u4214 ( .A0(n3453), .A1(n3590), .B0(n3591), .B1(n3279), 
        .C0(n3594), .Y(n1973) );
  AOI22_X0P5M_A12TR u4215 ( .A0(wtbldec[17]), .A1(n3560), .B0(wtblinc[17]), 
        .B1(n3561), .Y(n3594) );
  OAI221_X0P5M_A12TR u4216 ( .A0(n3158), .A1(n3590), .B0(n3591), .B1(n3294), 
        .C0(n3595), .Y(n1972) );
  AOI22_X0P5M_A12TR u4217 ( .A0(wtbldec[18]), .A1(n3560), .B0(wtblinc[18]), 
        .B1(n3561), .Y(n3595) );
  OAI221_X0P5M_A12TR u4218 ( .A0(n3458), .A1(n3590), .B0(n3591), .B1(n3309), 
        .C0(n3596), .Y(n1971) );
  AOI22_X0P5M_A12TR u4219 ( .A0(wtbldec[19]), .A1(n3560), .B0(wtblinc[19]), 
        .B1(n3561), .Y(n3596) );
  OA21A1OI2_X0P5M_A12TR u4220 ( .A0(n3104), .A1(n3597), .B0(qfsm[0]), .C0(
        n3588), .Y(n3591) );
  NAND3_X0P5A_A12TR u4221 ( .A(n3268), .B(n3240), .C(n3589), .Y(n3590) );
  OAI221_X0P5M_A12TR u4222 ( .A0(n3598), .A1(n3259), .B0(n3067), .B1(n3599), 
        .C0(n3600), .Y(n1970) );
  AOI22_X0P5M_A12TR u4223 ( .A0(wtbldec[8]), .A1(n3560), .B0(wtblinc[8]), .B1(
        n3561), .Y(n3600) );
  OAI221_X0P5M_A12TR u4224 ( .A0(n3598), .A1(n3601), .B0(n3453), .B1(n3599), 
        .C0(n3602), .Y(n1969) );
  AOI22_X0P5M_A12TR u4225 ( .A0(wtbldec[9]), .A1(n3560), .B0(wtblinc[9]), .B1(
        n3561), .Y(n3602) );
  OAI221_X0P5M_A12TR u4226 ( .A0(n3598), .A1(n3603), .B0(n3158), .B1(n3599), 
        .C0(n3604), .Y(n1968) );
  AOI22_X0P5M_A12TR u4227 ( .A0(wtbldec[10]), .A1(n3560), .B0(wtblinc[10]), 
        .B1(n3561), .Y(n3604) );
  OAI221_X0P5M_A12TR u4228 ( .A0(n3598), .A1(n3605), .B0(n3458), .B1(n3599), 
        .C0(n3606), .Y(n1967) );
  AOI22_X0P5M_A12TR u4229 ( .A0(wtbldec[11]), .A1(n3560), .B0(wtblinc[11]), 
        .B1(n3561), .Y(n3606) );
  OAI221_X0P5M_A12TR u4230 ( .A0(n3598), .A1(n3607), .B0(n3148), .B1(n3599), 
        .C0(n3608), .Y(n1966) );
  AOI22_X0P5M_A12TR u4231 ( .A0(wtbldec[12]), .A1(n3560), .B0(wtblinc[12]), 
        .B1(n3561), .Y(n3608) );
  OAI221_X0P5M_A12TR u4232 ( .A0(n3598), .A1(n3609), .B0(n3466), .B1(n3599), 
        .C0(n3610), .Y(n1965) );
  AOI22_X0P5M_A12TR u4233 ( .A0(wtbldec[13]), .A1(n3560), .B0(wtblinc[13]), 
        .B1(n3561), .Y(n3610) );
  OAI221_X0P5M_A12TR u4234 ( .A0(n3598), .A1(n3611), .B0(n3468), .B1(n3599), 
        .C0(n3612), .Y(n1964) );
  AOI22_X0P5M_A12TR u4235 ( .A0(wtbldec[14]), .A1(n3560), .B0(wtblinc[14]), 
        .B1(n3561), .Y(n3612) );
  OAI221_X0P5M_A12TR u4236 ( .A0(n3598), .A1(n3613), .B0(n3470), .B1(n3599), 
        .C0(n3614), .Y(n1963) );
  AOI22_X0P5M_A12TR u4237 ( .A0(wtbldec[15]), .A1(n3560), .B0(wtblinc[15]), 
        .B1(n3561), .Y(n3614) );
  AND3_X0P5M_A12TR u4238 ( .A(rmxtbl[0]), .B(n3615), .C(n3589), .Y(n3561) );
  OAI31_X0P5M_A12TR u4239 ( .A0(n3616), .A1(n3138), .A2(n3617), .B0(n3238), 
        .Y(n3615) );
  AND3_X0P5M_A12TR u4240 ( .A(n3247), .B(n3618), .C(n3589), .Y(n3560) );
  NAND3_X0P5A_A12TR u4241 ( .A(n3118), .B(n3240), .C(n3589), .Y(n3599) );
  AOI211_X0P5M_A12TR u4242 ( .A0(n3258), .A1(qfsm[0]), .B0(n3248), .C0(n3588), 
        .Y(n3598) );
  NAND2_X0P5A_A12TR u4243 ( .A(n3589), .B(n3619), .Y(n3588) );
  OAI31_X0P5M_A12TR u4244 ( .A0(n3616), .A1(n3617), .A2(n3618), .B0(n3143), 
        .Y(n3619) );
  OA21A1OI2_X0P5M_A12TR u4245 ( .A0(n3616), .A1(n3620), .B0(n3247), .C0(n3476), 
        .Y(n3589) );
  XNOR2_X0P5M_A12TR u4246 ( .A(rmxtbl[1]), .B(rmxtbl[0]), .Y(n3620) );
  OAI211_X0P5M_A12TR u4247 ( .A0(n3577), .A1(n3621), .B0(n3622), .C0(n3623), 
        .Y(n1962) );
  OAI21_X0P5M_A12TR u4248 ( .A0(rpcnxt[2]), .A1(n3624), .B0(n3625), .Y(n3623)
         );
  NAND2_X0P5A_A12TR u4249 ( .A(iwb_adr_o[3]), .B(n3626), .Y(n3622) );
  INV_X0P5B_A12TR u4250 ( .A(wtblat[3]), .Y(n3577) );
  OAI211_X0P5M_A12TR u4251 ( .A0(n3627), .A1(n3628), .B0(n3629), .C0(n3630), 
        .Y(n1961) );
  AOI22_X0P5M_A12TR u4252 ( .A0(iwb_adr_o[4]), .A1(n3626), .B0(n3631), .B1(
        wtblat[4]), .Y(n3630) );
  INV_X0P5B_A12TR u4253 ( .A(n3621), .Y(n3631) );
  NAND3B_X0P5M_A12TR u4254 ( .AN(rintf[1]), .B(rintf[0]), .C(n3625), .Y(n3629)
         );
  INV_X0P5B_A12TR u4255 ( .A(n3632), .Y(n3627) );
  AO1B2_X0P5M_A12TR u4256 ( .B0(rprodh[0]), .B1(n3633), .A0N(n3634), .Y(n1960)
         );
  AOI22_X0P5M_A12TR u4257 ( .A0(n17900), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[0]), .Y(n3634) );
  AO1B2_X0P5M_A12TR u4258 ( .B0(rprodh[1]), .B1(n3633), .A0N(n3637), .Y(n1959)
         );
  AOI22_X0P5M_A12TR u4259 ( .A0(n1791), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[1]), .Y(n3637) );
  AO1B2_X0P5M_A12TR u4260 ( .B0(rprodh[2]), .B1(n3633), .A0N(n3638), .Y(n1958)
         );
  AOI22_X0P5M_A12TR u4261 ( .A0(n1792), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[2]), .Y(n3638) );
  AO1B2_X0P5M_A12TR u4262 ( .B0(rprodh[3]), .B1(n3633), .A0N(n3639), .Y(n1957)
         );
  AOI22_X0P5M_A12TR u4263 ( .A0(n1793), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[3]), .Y(n3639) );
  AO1B2_X0P5M_A12TR u4264 ( .B0(rprodh[4]), .B1(n3633), .A0N(n3640), .Y(n1956)
         );
  AOI22_X0P5M_A12TR u4265 ( .A0(n1794), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[4]), .Y(n3640) );
  AO1B2_X0P5M_A12TR u4266 ( .B0(n3633), .B1(rprodh[5]), .A0N(n3641), .Y(n1955)
         );
  AOI22_X0P5M_A12TR u4267 ( .A0(n1795), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[5]), .Y(n3641) );
  AO1B2_X0P5M_A12TR u4268 ( .B0(rprodh[6]), .B1(n3633), .A0N(n3642), .Y(n1954)
         );
  AOI22_X0P5M_A12TR u4269 ( .A0(n1796), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[6]), .Y(n3642) );
  AO1B2_X0P5M_A12TR u4270 ( .B0(rprodh[7]), .B1(n3633), .A0N(n3643), .Y(n1953)
         );
  AOI22_X0P5M_A12TR u4271 ( .A0(n17970), .A1(n3635), .B0(n3636), .B1(
        dwb_dat_o[7]), .Y(n3643) );
  NOR3_X0P5A_A12TR u4272 ( .A(n3597), .B(n3633), .C(n3644), .Y(n3636) );
  AOI21_X0P5M_A12TR u4273 ( .A0(n3645), .A1(n3120), .B0(n3633), .Y(n3635) );
  AOI21_X0P5M_A12TR u4274 ( .A0(n3120), .A1(n3646), .B0(n3647), .Y(n3633) );
  AO1B2_X0P5M_A12TR u4275 ( .B0(rprodl[0]), .B1(n3648), .A0N(n3649), .Y(n1952)
         );
  AOI22_X0P5M_A12TR u4276 ( .A0(n17820), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[0]), .Y(n3649) );
  AO1B2_X0P5M_A12TR u4277 ( .B0(rprodl[1]), .B1(n3648), .A0N(n3652), .Y(n1951)
         );
  AOI22_X0P5M_A12TR u4278 ( .A0(n1783), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[1]), .Y(n3652) );
  AO1B2_X0P5M_A12TR u4279 ( .B0(rprodl[2]), .B1(n3648), .A0N(n3653), .Y(n1950)
         );
  AOI22_X0P5M_A12TR u4280 ( .A0(n17840), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[2]), .Y(n3653) );
  AO1B2_X0P5M_A12TR u4281 ( .B0(rprodl[3]), .B1(n3648), .A0N(n3654), .Y(n1949)
         );
  AOI22_X0P5M_A12TR u4282 ( .A0(n1785), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[3]), .Y(n3654) );
  AO1B2_X0P5M_A12TR u4283 ( .B0(rprodl[4]), .B1(n3648), .A0N(n3655), .Y(n1948)
         );
  AOI22_X0P5M_A12TR u4284 ( .A0(n1786), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[4]), .Y(n3655) );
  AO1B2_X0P5M_A12TR u4285 ( .B0(n3648), .B1(rprodl[5]), .A0N(n3656), .Y(n1947)
         );
  AOI22_X0P5M_A12TR u4286 ( .A0(n17870), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[5]), .Y(n3656) );
  MXIT2_X0P5M_A12TR u4287 ( .A(n3657), .B(n3658), .S0(n3092), .Y(n1946) );
  INV_X0P5B_A12TR u4288 ( .A(rsfrdat[5]), .Y(n3658) );
  NOR3_X0P5A_A12TR u4289 ( .A(n3659), .B(n3660), .C(n3661), .Y(n3657) );
  OAI221_X0P5M_A12TR u4290 ( .A0(n3662), .A1(n3663), .B0(n3096), .B1(n3664), 
        .C0(n3665), .Y(n3661) );
  AOI222_X0P5M_A12TR u4291 ( .A0(rpclatu[5]), .A1(n3103), .B0(rpclath[5]), 
        .B1(n3108), .C0(wstkw[13]), .C1(n3102), .Y(n3665) );
  OAI221_X0P5M_A12TR u4292 ( .A0(n3666), .A1(n3667), .B0(n3668), .B1(n3669), 
        .C0(n3670), .Y(n3660) );
  AOI222_X0P5M_A12TR u4293 ( .A0(rtblptru[5]), .A1(n3268), .B0(wfilebsr[13]), 
        .B1(n3111), .C0(rwreg[5]), .C1(n3112), .Y(n3670) );
  INV_X0P5B_A12TR u4294 ( .A(n3671), .Y(n3112) );
  NAND4_X0P5A_A12TR u4295 ( .A(n3672), .B(n3673), .C(n3674), .D(n3675), .Y(
        n3659) );
  AOI222_X0P5M_A12TR u4296 ( .A0(rfsr1h[5]), .A1(n3117), .B0(wtblat[13]), .B1(
        n3118), .C0(wtblat[5]), .C1(n3119), .Y(n3675) );
  INV_X0P5B_A12TR u4297 ( .A(n3587), .Y(n3119) );
  NAND2_X0P5A_A12TR u4298 ( .A(n3676), .B(n3677), .Y(n3587) );
  INV_X0P5B_A12TR u4299 ( .A(n3258), .Y(n3118) );
  NAND2_X0P5A_A12TR u4300 ( .A(n3678), .B(n3677), .Y(n3258) );
  AND3_X0P5M_A12TR u4301 ( .A(n3676), .B(n3679), .C(n3680), .Y(n3117) );
  AOI222_X0P5M_A12TR u4302 ( .A0(rprodh[5]), .A1(n3120), .B0(rfsr1l[5]), .B1(
        n3121), .C0(rfsr2l[5]), .C1(n3122), .Y(n3674) );
  AND2_X0P5M_A12TR u4303 ( .A(n3316), .B(n3263), .Y(n3122) );
  AND3_X0P5M_A12TR u4304 ( .A(n3263), .B(n3679), .C(n3680), .Y(n3121) );
  INV_X0P5B_A12TR u4305 ( .A(n3644), .Y(n3120) );
  NAND2_X0P5A_A12TR u4306 ( .A(n3677), .B(n3317), .Y(n3644) );
  AOI222_X0P5M_A12TR u4307 ( .A0(rfsr0l[5]), .A1(n3123), .B0(n3124), .B1(n3681), .C0(rprng[5]), .C1(n3126), .Y(n3673) );
  NOR2_X0P5A_A12TR u4308 ( .A(n3682), .B(dwb_adr_o[5]), .Y(n3126) );
  INV_X0P5B_A12TR u4309 ( .A(n3546), .Y(n3124) );
  NAND2_X0P5A_A12TR u4310 ( .A(n3316), .B(n3676), .Y(n3546) );
  AND4_X0P5M_A12TR u4311 ( .A(dwb_adr_o[3]), .B(dwb_adr_o[4]), .C(n3683), .D(
        n3684), .Y(n3316) );
  AND3_X0P5M_A12TR u4312 ( .A(n3263), .B(dwb_adr_o[3]), .C(n3680), .Y(n3123)
         );
  AOI22_X0P5M_A12TR u4313 ( .A0(rfsr0h[5]), .A1(n3127), .B0(rprodl[5]), .B1(
        n3128), .Y(n3672) );
  INV_X0P5B_A12TR u4314 ( .A(n3254), .Y(n3127) );
  NAND3_X0P5A_A12TR u4315 ( .A(n3676), .B(dwb_adr_o[3]), .C(n3680), .Y(n3254)
         );
  AO1B2_X0P5M_A12TR u4316 ( .B0(rprodl[6]), .B1(n3648), .A0N(n3685), .Y(n1945)
         );
  AOI22_X0P5M_A12TR u4317 ( .A0(n1788), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[6]), .Y(n3685) );
  AO1B2_X0P5M_A12TR u4318 ( .B0(rprodl[7]), .B1(n3648), .A0N(n3686), .Y(n1944)
         );
  AOI22_X0P5M_A12TR u4319 ( .A0(n1789), .A1(n3650), .B0(n3651), .B1(
        dwb_dat_o[7]), .Y(n3686) );
  NOR3_X0P5A_A12TR u4320 ( .A(n3597), .B(n3648), .C(n3687), .Y(n3651) );
  AOI21_X0P5M_A12TR u4321 ( .A0(n3645), .A1(n3128), .B0(n3648), .Y(n3650) );
  AOI21_X0P5M_A12TR u4322 ( .A0(n3128), .A1(n3646), .B0(n3647), .Y(n3648) );
  AND4_X0P5M_A12TR u4323 ( .A(rmxalu[0]), .B(n3688), .C(n3549), .D(n3551), .Y(
        n3647) );
  AND4_X0P5M_A12TR u4324 ( .A(rmxdst[0]), .B(rmxalu[3]), .C(rmxalu[1]), .D(
        rmxalu[2]), .Y(n3549) );
  INV_X0P5B_A12TR u4325 ( .A(n3687), .Y(n3128) );
  NAND3_X0P5A_A12TR u4326 ( .A(n3262), .B(dwb_adr_o[5]), .C(n3678), .Y(n3687)
         );
  OAI21_X0P5M_A12TR u4327 ( .A0(n3309), .A1(n3621), .B0(n3689), .Y(n1937) );
  AOI22_X0P5M_A12TR u4328 ( .A0(rpcnxt[18]), .A1(n3632), .B0(iwb_adr_o[19]), 
        .B1(n3626), .Y(n3689) );
  INV_X0P5B_A12TR u4329 ( .A(wtblat[19]), .Y(n3309) );
  OAI21_X0P5M_A12TR u4330 ( .A0(n3294), .A1(n3621), .B0(n3690), .Y(n1936) );
  AOI22_X0P5M_A12TR u4331 ( .A0(rpcnxt[17]), .A1(n3632), .B0(iwb_adr_o[18]), 
        .B1(n3626), .Y(n3690) );
  INV_X0P5B_A12TR u4332 ( .A(wtblat[18]), .Y(n3294) );
  OAI21_X0P5M_A12TR u4333 ( .A0(n3279), .A1(n3621), .B0(n3691), .Y(n1935) );
  AOI22_X0P5M_A12TR u4334 ( .A0(rpcnxt[16]), .A1(n3632), .B0(iwb_adr_o[17]), 
        .B1(n3626), .Y(n3691) );
  INV_X0P5B_A12TR u4335 ( .A(wtblat[17]), .Y(n3279) );
  OAI21_X0P5M_A12TR u4336 ( .A0(n3592), .A1(n3621), .B0(n3692), .Y(n1934) );
  AOI22_X0P5M_A12TR u4337 ( .A0(rpcnxt[15]), .A1(n3632), .B0(iwb_adr_o[16]), 
        .B1(n3626), .Y(n3692) );
  INV_X0P5B_A12TR u4338 ( .A(wtblat[16]), .Y(n3592) );
  OAI21_X0P5M_A12TR u4339 ( .A0(n3613), .A1(n3621), .B0(n3693), .Y(n1933) );
  AOI22_X0P5M_A12TR u4340 ( .A0(rpcnxt[14]), .A1(n3632), .B0(iwb_adr_o[15]), 
        .B1(n3626), .Y(n3693) );
  INV_X0P5B_A12TR u4341 ( .A(wtblat[15]), .Y(n3613) );
  OAI21_X0P5M_A12TR u4342 ( .A0(n3611), .A1(n3621), .B0(n3694), .Y(n1932) );
  AOI22_X0P5M_A12TR u4343 ( .A0(rpcnxt[13]), .A1(n3632), .B0(iwb_adr_o[14]), 
        .B1(n3626), .Y(n3694) );
  INV_X0P5B_A12TR u4344 ( .A(wtblat[14]), .Y(n3611) );
  OAI21_X0P5M_A12TR u4345 ( .A0(n3609), .A1(n3621), .B0(n3695), .Y(n1931) );
  AOI22_X0P5M_A12TR u4346 ( .A0(rpcnxt[12]), .A1(n3632), .B0(iwb_adr_o[13]), 
        .B1(n3626), .Y(n3695) );
  INV_X0P5B_A12TR u4347 ( .A(wtblat[13]), .Y(n3609) );
  OAI21_X0P5M_A12TR u4348 ( .A0(n3607), .A1(n3621), .B0(n3696), .Y(n1930) );
  AOI22_X0P5M_A12TR u4349 ( .A0(rpcnxt[11]), .A1(n3632), .B0(iwb_adr_o[12]), 
        .B1(n3626), .Y(n3696) );
  INV_X0P5B_A12TR u4350 ( .A(wtblat[12]), .Y(n3607) );
  OAI21_X0P5M_A12TR u4351 ( .A0(n3605), .A1(n3621), .B0(n3697), .Y(n1929) );
  AOI22_X0P5M_A12TR u4352 ( .A0(rpcnxt[10]), .A1(n3632), .B0(iwb_adr_o[11]), 
        .B1(n3626), .Y(n3697) );
  INV_X0P5B_A12TR u4353 ( .A(wtblat[11]), .Y(n3605) );
  OAI21_X0P5M_A12TR u4354 ( .A0(n3603), .A1(n3621), .B0(n3698), .Y(n1928) );
  AOI22_X0P5M_A12TR u4355 ( .A0(rpcnxt[9]), .A1(n3632), .B0(iwb_adr_o[10]), 
        .B1(n3626), .Y(n3698) );
  INV_X0P5B_A12TR u4356 ( .A(wtblat[10]), .Y(n3603) );
  OAI21_X0P5M_A12TR u4357 ( .A0(n3601), .A1(n3621), .B0(n3699), .Y(n1927) );
  AOI22_X0P5M_A12TR u4358 ( .A0(rpcnxt[8]), .A1(n3632), .B0(iwb_adr_o[9]), 
        .B1(n3626), .Y(n3699) );
  INV_X0P5B_A12TR u4359 ( .A(wtblat[9]), .Y(n3601) );
  OAI21_X0P5M_A12TR u4360 ( .A0(n3259), .A1(n3621), .B0(n3700), .Y(n1926) );
  AOI22_X0P5M_A12TR u4361 ( .A0(rpcnxt[7]), .A1(n3632), .B0(iwb_adr_o[8]), 
        .B1(n3626), .Y(n3700) );
  INV_X0P5B_A12TR u4362 ( .A(wtblat[8]), .Y(n3259) );
  OAI21_X0P5M_A12TR u4363 ( .A0(n3585), .A1(n3621), .B0(n3701), .Y(n1925) );
  AOI22_X0P5M_A12TR u4364 ( .A0(rpcnxt[6]), .A1(n3632), .B0(iwb_adr_o[7]), 
        .B1(n3626), .Y(n3701) );
  INV_X0P5B_A12TR u4365 ( .A(wtblat[7]), .Y(n3585) );
  OAI21_X0P5M_A12TR u4366 ( .A0(n3583), .A1(n3621), .B0(n3702), .Y(n1924) );
  AOI22_X0P5M_A12TR u4367 ( .A0(rpcnxt[5]), .A1(n3632), .B0(iwb_adr_o[6]), 
        .B1(n3626), .Y(n3702) );
  INV_X0P5B_A12TR u4368 ( .A(wtblat[6]), .Y(n3583) );
  OAI21_X0P5M_A12TR u4369 ( .A0(n3581), .A1(n3621), .B0(n3703), .Y(n1923) );
  AOI22_X0P5M_A12TR u4370 ( .A0(rpcnxt[4]), .A1(n3632), .B0(iwb_adr_o[5]), 
        .B1(n3626), .Y(n3703) );
  INV_X0P5B_A12TR u4371 ( .A(wtblat[5]), .Y(n3581) );
  OAI21_X0P5M_A12TR u4372 ( .A0(n3575), .A1(n3621), .B0(n3704), .Y(n1922) );
  AOI22_X0P5M_A12TR u4373 ( .A0(rpcnxt[1]), .A1(n3632), .B0(iwb_adr_o[2]), 
        .B1(n3626), .Y(n3704) );
  INV_X0P5B_A12TR u4374 ( .A(wtblat[2]), .Y(n3575) );
  OAI21_X0P5M_A12TR u4375 ( .A0(n3573), .A1(n3621), .B0(n3705), .Y(n1921) );
  AOI22_X0P5M_A12TR u4376 ( .A0(rpcnxt[0]), .A1(n3632), .B0(iwb_adr_o[1]), 
        .B1(n3626), .Y(n3705) );
  OAI211_X0P5M_A12TR u4377 ( .A0(qfsm[1]), .A1(n3706), .B0(n3054), .C0(qfsm[0]), .Y(n3626) );
  NOR2_X0P5A_A12TR u4378 ( .A(n3624), .B(n3228), .Y(n3632) );
  NAND3_X0P5A_A12TR u4379 ( .A(n3054), .B(n3706), .C(n3460), .Y(n3621) );
  INV_X0P5B_A12TR u4380 ( .A(wtblat[1]), .Y(n3573) );
  AOI221_X0P5M_A12TR u4381 ( .A0(n3707), .A1(n3688), .B0(n3708), .B1(n3074), 
        .C0(n3709), .Y(n1906) );
  MXT4_X0P5M_A12TR u4382 ( .A(n3710), .B(n3711), .C(n3712), .D(n3713), .S0(
        n3714), .S1(rmxskp[1]), .Y(n3707) );
  MXIT2_X0P5M_A12TR u4383 ( .A(n3715), .B(n3155), .S0(n3710), .Y(n3713) );
  NOR2_X0P5A_A12TR u4384 ( .A(n3716), .B(n3710), .Y(n3712) );
  AND2_X0P5M_A12TR u4385 ( .A(n3155), .B(rmxskp[0]), .Y(n3711) );
  NOR2_X0P5A_A12TR u4386 ( .A(n3717), .B(n3718), .Y(n3155) );
  NAND4_X0P5A_A12TR u4387 ( .A(n3067), .B(n3453), .C(n3158), .D(n3458), .Y(
        n3718) );
  NAND4_X0P5A_A12TR u4388 ( .A(n3148), .B(n3466), .C(n3468), .D(n3470), .Y(
        n3717) );
  OAI221_X0P5M_A12TR u4389 ( .A0(n3403), .A1(n3719), .B0(n3720), .B1(n3721), 
        .C0(n3722), .Y(n1904) );
  AOI222_X0P5M_A12TR u4390 ( .A0(n3723), .A1(n3333), .B0(n3724), .B1(rfsr0h[6]), .C0(n3725), .C1(rfsr1h[6]), .Y(n3722) );
  INV_X0P5B_A12TR u4391 ( .A(n1941), .Y(n3333) );
  INV_X0P5B_A12TR u4392 ( .A(rdwbadr[14]), .Y(n3721) );
  OAI22_X0P5M_A12TR u4393 ( .A0(n3726), .A1(n3092), .B0(n3727), .B1(n3728), 
        .Y(n1902) );
  INV_X0P5B_A12TR u4394 ( .A(rsfrstb), .Y(n3728) );
  NAND4_X0P5A_A12TR u4395 ( .A(n3727), .B(n3729), .C(n3730), .D(n3731), .Y(
        n3092) );
  AO21A1AI2_X0P5M_A12TR u4396 ( .A0(dwb_adr_o[5]), .A1(n3732), .B0(n3733), 
        .C0(n3262), .Y(n3731) );
  AO21A1AI2_X0P5M_A12TR u4397 ( .A0(dwb_adr_o[2]), .A1(n3682), .B0(n3678), 
        .C0(n3684), .Y(n3730) );
  OAI31_X0P5M_A12TR u4398 ( .A0(n3684), .A1(dwb_adr_o[2]), .A2(n3678), .B0(
        n3734), .Y(n3729) );
  NOR2_X0P5A_A12TR u4399 ( .A(n3735), .B(n3708), .Y(n3727) );
  OAI221_X0P5M_A12TR u4400 ( .A0(n3736), .A1(n3737), .B0(n3738), .B1(n3739), 
        .C0(n3740), .Y(n1901) );
  AOI221_X0P5M_A12TR u4401 ( .A0(rmask[0]), .A1(n3741), .B0(n3742), .B1(n3743), 
        .C0(n3744), .Y(n3740) );
  NAND4_X0P5A_A12TR u4402 ( .A(n3745), .B(n3746), .C(n3747), .D(n3748), .Y(
        n1899) );
  AOI211_X0P5M_A12TR u4403 ( .A0(n3749), .A1(n3750), .B0(n3751), .C0(n3752), 
        .Y(n3748) );
  OA21A1OI2_X0P5M_A12TR u4404 ( .A0(wneg[0]), .A1(n3753), .B0(n3754), .C0(
        n3739), .Y(n3752) );
  AOI31_X0P5M_A12TR u4405 ( .A0(n3754), .A1(n3755), .A2(n3756), .B0(n4423), 
        .Y(n3751) );
  MXIT2_X0P5M_A12TR u4406 ( .A(n3757), .B(n3758), .S0(n3739), .Y(n3756) );
  INV_X0P5B_A12TR u4407 ( .A(rsrc[0]), .Y(n3739) );
  MXIT2_X0P5M_A12TR u4408 ( .A(n3179), .B(n4430), .S0(n3550), .Y(n3749) );
  AOI22_X0P5M_A12TR u4409 ( .A0(n3759), .A1(rtgt[1]), .B0(n3760), .B1(rtgt[4]), 
        .Y(n3747) );
  AOI222_X0P5M_A12TR u4410 ( .A0(wsubc[0]), .A1(n3761), .B0(wsub[0]), .B1(
        n3762), .C0(wadd[0]), .C1(n3763), .Y(n3746) );
  AOI22_X0P5M_A12TR u4411 ( .A0(waddc[0]), .A1(n3764), .B0(dwb_dat_o[0]), .B1(
        n3765), .Y(n3745) );
  NAND4_X0P5A_A12TR u4412 ( .A(n3766), .B(n3767), .C(n3768), .D(n3769), .Y(
        n1897) );
  AOI211_X0P5M_A12TR u4413 ( .A0(n3770), .A1(n3759), .B0(n3771), .C0(n3772), 
        .Y(n3769) );
  OA21A1OI2_X0P5M_A12TR u4414 ( .A0(rtgt[7]), .A1(n3753), .B0(n3754), .C0(
        n3773), .Y(n3772) );
  AOI21_X0P5M_A12TR u4415 ( .A0(n3774), .A1(n3754), .B0(n4430), .Y(n3771) );
  MXIT2_X0P5M_A12TR u4416 ( .A(n3757), .B(n3758), .S0(n3773), .Y(n3774) );
  MXIT2_X0P5M_A12TR u4417 ( .A(n3179), .B(n4423), .S0(n3550), .Y(n3770) );
  AOI222_X0P5M_A12TR u4418 ( .A0(wsub[7]), .A1(n3762), .B0(n3750), .B1(rtgt[6]), .C0(n3760), .C1(rtgt[3]), .Y(n3768) );
  AOI222_X0P5M_A12TR u4419 ( .A0(wsubc[7]), .A1(n3761), .B0(wneg[7]), .B1(
        n3775), .C0(wadd[7]), .C1(n3763), .Y(n3767) );
  AOI22_X0P5M_A12TR u4420 ( .A0(waddc[7]), .A1(n3764), .B0(dwb_dat_o[7]), .B1(
        n3765), .Y(n3766) );
  OAI222_X0P5M_A12TR u4421 ( .A0(n3470), .A1(n3776), .B0(n3777), .B1(n3778), 
        .C0(qena[3]), .C1(n3779), .Y(n1895) );
  INV_X0P5B_A12TR u4422 ( .A(wpclat[6]), .Y(n3779) );
  OAI221_X0P5M_A12TR u4423 ( .A0(n3780), .A1(n3737), .B0(n3738), .B1(n3773), 
        .C0(n3781), .Y(n1893) );
  AOI221_X0P5M_A12TR u4424 ( .A0(rmask[7]), .A1(n3741), .B0(n3742), .B1(n3782), 
        .C0(n3744), .Y(n3781) );
  INV_X0P5B_A12TR u4425 ( .A(rsrc[7]), .Y(n3773) );
  MXIT2_X0P5M_A12TR u4426 ( .A(n3783), .B(n3716), .S0(n3784), .Y(n1891) );
  MXT4_X0P5M_A12TR u4427 ( .A(n3785), .B(n3786), .C(n3787), .D(n3788), .S0(
        rmxbcc[2]), .S1(rmxbcc[1]), .Y(n3783) );
  XNOR2_X0P5M_A12TR u4428 ( .A(rmxbcc[0]), .B(rn), .Y(n3788) );
  XNOR2_X0P5M_A12TR u4429 ( .A(rmxbcc[0]), .B(wrrc_7_), .Y(n3787) );
  XNOR2_X0P5M_A12TR u4430 ( .A(rmxbcc[0]), .B(rov), .Y(n3786) );
  XNOR2_X0P5M_A12TR u4431 ( .A(rmxbcc[0]), .B(rz), .Y(n3785) );
  OAI211_X0P5M_A12TR u4432 ( .A0(qena[1]), .A1(n3789), .B0(n3790), .C0(n3791), 
        .Y(n1889) );
  AOI222_X0P5M_A12TR u4433 ( .A0(wpcinc[0]), .A1(n3792), .B0(n386), .B1(n3793), 
        .C0(n3794), .C1(wstkw[1]), .Y(n3791) );
  AOI22_X0P5M_A12TR u4434 ( .A0(n366), .A1(n3795), .B0(n3796), .B1(rireg[0]), 
        .Y(n3790) );
  OAI222_X0P5M_A12TR u4435 ( .A0(n3453), .A1(n3776), .B0(n3789), .B1(n3778), 
        .C0(qena[3]), .C1(n3797), .Y(n1887) );
  INV_X0P5B_A12TR u4436 ( .A(wpclat[0]), .Y(n3797) );
  INV_X0P5B_A12TR u4437 ( .A(rpcnxt[0]), .Y(n3789) );
  OAI221_X0P5M_A12TR u4438 ( .A0(n3798), .A1(n3737), .B0(n3738), .B1(n3799), 
        .C0(n3800), .Y(n1885) );
  AOI221_X0P5M_A12TR u4439 ( .A0(rmask[1]), .A1(n3741), .B0(n3742), .B1(n3801), 
        .C0(n3744), .Y(n3800) );
  NAND4_X0P5A_A12TR u4440 ( .A(n3802), .B(n3803), .C(n3804), .D(n3805), .Y(
        n1883) );
  AOI211_X0P5M_A12TR u4441 ( .A0(n3750), .A1(wneg[0]), .B0(n3806), .C0(n3807), 
        .Y(n3805) );
  AOI21_X0P5M_A12TR u4442 ( .A0(n3808), .A1(n3754), .B0(n4424), .Y(n3807) );
  MXIT2_X0P5M_A12TR u4443 ( .A(n3757), .B(n3758), .S0(n3799), .Y(n3808) );
  OA21A1OI2_X0P5M_A12TR u4444 ( .A0(rtgt[1]), .A1(n3753), .B0(n3754), .C0(
        n3799), .Y(n3806) );
  INV_X0P5B_A12TR u4445 ( .A(rsrc[1]), .Y(n3799) );
  AOI222_X0P5M_A12TR u4446 ( .A0(wsub[1]), .A1(n3762), .B0(n3759), .B1(rtgt[2]), .C0(n3760), .C1(rtgt[5]), .Y(n3804) );
  AOI222_X0P5M_A12TR u4447 ( .A0(wsubc[1]), .A1(n3761), .B0(wneg[1]), .B1(
        n3775), .C0(wadd[1]), .C1(n3763), .Y(n3803) );
  AOI22_X0P5M_A12TR u4448 ( .A0(waddc[1]), .A1(n3764), .B0(dwb_dat_o[1]), .B1(
        n3765), .Y(n3802) );
  NAND4_X0P5A_A12TR u4449 ( .A(n3809), .B(n3810), .C(n3811), .D(n3812), .Y(
        n1881) );
  AOI222_X0P5M_A12TR u4450 ( .A0(wfsrplusw1[1]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[1]), .C0(n3815), .C1(wfsrinc2[1]), .Y(n3812) );
  AOI222_X0P5M_A12TR u4451 ( .A0(n3724), .A1(rfsr0l[1]), .B0(wfsrplusw2[1]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[1]), .Y(n3811) );
  AOI222_X0P5M_A12TR u4452 ( .A0(n3723), .A1(rfsr2l[1]), .B0(wfsrplusw0[1]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[1]), .Y(n3810) );
  AOI222_X0P5M_A12TR u4453 ( .A0(dwb_adr_o[1]), .A1(n3819), .B0(n3820), .B1(
        rromlat[1]), .C0(reaptr[1]), .C1(n3821), .Y(n3809) );
  OAI221_X0P5M_A12TR u4454 ( .A0(n3822), .A1(n3737), .B0(n3738), .B1(n3823), 
        .C0(n3824), .Y(n1879) );
  AOI221_X0P5M_A12TR u4455 ( .A0(rmask[4]), .A1(n3741), .B0(n3742), .B1(n3825), 
        .C0(n3744), .Y(n3824) );
  NAND4_X0P5A_A12TR u4456 ( .A(n3826), .B(n3827), .C(n3828), .D(n3829), .Y(
        n1877) );
  AOI211_X0P5M_A12TR u4457 ( .A0(n3750), .A1(rtgt[3]), .B0(n3830), .C0(n3831), 
        .Y(n3829) );
  AOI21_X0P5M_A12TR u4458 ( .A0(n3832), .A1(n3754), .B0(n4427), .Y(n3831) );
  MXIT2_X0P5M_A12TR u4459 ( .A(n3757), .B(n3758), .S0(n3823), .Y(n3832) );
  OA21A1OI2_X0P5M_A12TR u4460 ( .A0(rtgt[4]), .A1(n3753), .B0(n3754), .C0(
        n3823), .Y(n3830) );
  INV_X0P5B_A12TR u4461 ( .A(rsrc[4]), .Y(n3823) );
  AOI222_X0P5M_A12TR u4462 ( .A0(wsub[4]), .A1(n3762), .B0(n3759), .B1(rtgt[5]), .C0(n3760), .C1(wneg[0]), .Y(n3828) );
  AOI222_X0P5M_A12TR u4463 ( .A0(wsubc[4]), .A1(n3761), .B0(wneg[4]), .B1(
        n3775), .C0(wadd[4]), .C1(n3763), .Y(n3827) );
  AOI22_X0P5M_A12TR u4464 ( .A0(waddc[4]), .A1(n3764), .B0(dwb_dat_o[4]), .B1(
        n3765), .Y(n3826) );
  NAND4_X0P5A_A12TR u4465 ( .A(n3833), .B(n3834), .C(n3835), .D(n3836), .Y(
        n1875) );
  AOI222_X0P5M_A12TR u4466 ( .A0(wfsrplusw1[4]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[4]), .C0(n3815), .C1(wfsrinc2[4]), .Y(n3836) );
  AOI222_X0P5M_A12TR u4467 ( .A0(n3724), .A1(rfsr0l[4]), .B0(wfsrplusw2[4]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[4]), .Y(n3835) );
  AOI222_X0P5M_A12TR u4468 ( .A0(n3723), .A1(rfsr2l[4]), .B0(wfsrplusw0[4]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[4]), .Y(n3834) );
  AOI222_X0P5M_A12TR u4469 ( .A0(dwb_adr_o[4]), .A1(n3819), .B0(n3820), .B1(
        rromlat[4]), .C0(reaptr[4]), .C1(n3821), .Y(n3833) );
  INV_X0P5B_A12TR u4470 ( .A(n3837), .Y(n1873) );
  AOI221_X0P5M_A12TR u4471 ( .A0(n3838), .A1(n3839), .B0(n3840), .B1(
        rstkptr_5_), .C0(n3841), .Y(n3837) );
  OAI22_X0P5M_A12TR u4472 ( .A0(n2746), .A1(n3842), .B0(n3843), .B1(n3466), 
        .Y(n3841) );
  INV_X0P5B_A12TR u4473 ( .A(n3844), .Y(n3839) );
  MXIT2_X0P5M_A12TR u4474 ( .A(n3845), .B(n3324), .S0(n3476), .Y(n1872) );
  NAND4_X0P5A_A12TR u4475 ( .A(wstkdec[3]), .B(wstkdec[2]), .C(wstkdec[4]), 
        .D(n3846), .Y(n3845) );
  NOR3_X0P5A_A12TR u4476 ( .A(n3847), .B(n214), .C(n2746), .Y(n3846) );
  INV_X0P5B_A12TR u4477 ( .A(wstkdec[1]), .Y(n3847) );
  OAI21_X0P5M_A12TR u4478 ( .A0(n3067), .A1(n3843), .B0(n3848), .Y(n1871) );
  MXIT2_X0P5M_A12TR u4479 ( .A(n3849), .B(n3840), .S0(n214), .Y(n3848) );
  NAND2_X0P5A_A12TR u4480 ( .A(n3844), .B(n3842), .Y(n3849) );
  MXIT2_X0P5M_A12TR u4481 ( .A(n3850), .B(n3099), .S0(n3476), .Y(n1870) );
  NAND4_X0P5A_A12TR u4482 ( .A(n3838), .B(n3851), .C(n214), .D(n3852), .Y(
        n3850) );
  NOR3_X0P5A_A12TR u4483 ( .A(wstkinc[2]), .B(wstkinc[4]), .C(wstkinc[3]), .Y(
        n3852) );
  XOR2_X0P5M_A12TR u4484 ( .A(rstkptr_5_), .B(add_1310_carry[5]), .Y(n3838) );
  OAI221_X0P5M_A12TR u4485 ( .A0(n3844), .A1(n3853), .B0(n3158), .B1(n3843), 
        .C0(n3854), .Y(n1869) );
  AOI22_X0P5M_A12TR u4486 ( .A0(n216), .A1(n3840), .B0(wstkdec[2]), .B1(n3855), 
        .Y(n3854) );
  OAI221_X0P5M_A12TR u4487 ( .A0(n3856), .A1(n3737), .B0(n3738), .B1(n3857), 
        .C0(n3858), .Y(n1868) );
  AOI221_X0P5M_A12TR u4488 ( .A0(rmask[2]), .A1(n3741), .B0(n3742), .B1(n3859), 
        .C0(n3744), .Y(n3858) );
  NAND4_X0P5A_A12TR u4489 ( .A(n3860), .B(n3861), .C(n3862), .D(n3863), .Y(
        n1866) );
  AOI211_X0P5M_A12TR u4490 ( .A0(n3750), .A1(rtgt[1]), .B0(n3864), .C0(n3865), 
        .Y(n3863) );
  AOI21_X0P5M_A12TR u4491 ( .A0(n3866), .A1(n3754), .B0(n4425), .Y(n3865) );
  MXIT2_X0P5M_A12TR u4492 ( .A(n3757), .B(n3758), .S0(n3857), .Y(n3866) );
  OA21A1OI2_X0P5M_A12TR u4493 ( .A0(rtgt[2]), .A1(n3753), .B0(n3754), .C0(
        n3857), .Y(n3864) );
  INV_X0P5B_A12TR u4494 ( .A(rsrc[2]), .Y(n3857) );
  AOI222_X0P5M_A12TR u4495 ( .A0(wsub[2]), .A1(n3762), .B0(n3759), .B1(rtgt[3]), .C0(n3760), .C1(rtgt[6]), .Y(n3862) );
  AOI222_X0P5M_A12TR u4496 ( .A0(wsubc[2]), .A1(n3761), .B0(wneg[2]), .B1(
        n3775), .C0(wadd[2]), .C1(n3763), .Y(n3861) );
  AOI22_X0P5M_A12TR u4497 ( .A0(waddc[2]), .A1(n3764), .B0(dwb_dat_o[2]), .B1(
        n3765), .Y(n3860) );
  OAI222_X0P5M_A12TR u4498 ( .A0(n3158), .A1(n3776), .B0(n3867), .B1(n3778), 
        .C0(qena[3]), .C1(n3868), .Y(n1864) );
  INV_X0P5B_A12TR u4499 ( .A(wpclat[1]), .Y(n3868) );
  OAI221_X0P5M_A12TR u4500 ( .A0(n3064), .A1(n3869), .B0(n3066), .B1(n3158), 
        .C0(n3870), .Y(n1862) );
  AOI22_X0P5M_A12TR u4501 ( .A0(n2747), .A1(n3069), .B0(n3871), .B1(wpclat[1]), 
        .Y(n3870) );
  INV_X0P5B_A12TR u4502 ( .A(wstkw[2]), .Y(n3869) );
  OAI211_X0P5M_A12TR u4503 ( .A0(qena[1]), .A1(n3867), .B0(n3872), .C0(n3873), 
        .Y(n1861) );
  AOI222_X0P5M_A12TR u4504 ( .A0(wpcinc[1]), .A1(n3792), .B0(n387), .B1(n3793), 
        .C0(n3794), .C1(wstkw[2]), .Y(n3873) );
  AOI22_X0P5M_A12TR u4505 ( .A0(n367), .A1(n3795), .B0(n3796), .B1(rireg[1]), 
        .Y(n3872) );
  INV_X0P5B_A12TR u4506 ( .A(rpcnxt[1]), .Y(n3867) );
  OAI211_X0P5M_A12TR u4507 ( .A0(qena[1]), .A1(n3874), .B0(n3875), .C0(n3876), 
        .Y(n1858) );
  AOI222_X0P5M_A12TR u4508 ( .A0(wpcinc[18]), .A1(n3792), .B0(n404), .B1(n3793), .C0(n3794), .C1(wstkw[19]), .Y(n3876) );
  AOI22_X0P5M_A12TR u4509 ( .A0(n384), .A1(n3795), .B0(n3796), .B1(rromlat[10]), .Y(n3875) );
  OAI222_X0P5M_A12TR u4510 ( .A0(n3877), .A1(n3776), .B0(n3874), .B1(n3778), 
        .C0(qena[3]), .C1(n3878), .Y(n1856) );
  INV_X0P5B_A12TR u4511 ( .A(rpcnxt[18]), .Y(n3874) );
  OAI221_X0P5M_A12TR u4512 ( .A0(n3879), .A1(n3306), .B0(n3458), .B1(n3880), 
        .C0(n3881), .Y(n1854) );
  AOI22_X0P5M_A12TR u4513 ( .A0(n2782), .A1(n3069), .B0(wpclat[18]), .B1(n3871), .Y(n3881) );
  INV_X0P5B_A12TR u4514 ( .A(wstkw[19]), .Y(n3306) );
  OAI221_X0P5M_A12TR u4515 ( .A0(n3882), .A1(n3737), .B0(n3738), .B1(n3883), 
        .C0(n3884), .Y(n1853) );
  AOI221_X0P5M_A12TR u4516 ( .A0(rmask[3]), .A1(n3741), .B0(n3742), .B1(n3885), 
        .C0(n3744), .Y(n3884) );
  NAND4_X0P5A_A12TR u4517 ( .A(n3886), .B(n3887), .C(n3888), .D(n3889), .Y(
        n1851) );
  AOI211_X0P5M_A12TR u4518 ( .A0(n3750), .A1(rtgt[2]), .B0(n3890), .C0(n3891), 
        .Y(n3889) );
  AOI21_X0P5M_A12TR u4519 ( .A0(n3892), .A1(n3754), .B0(n4426), .Y(n3891) );
  MXIT2_X0P5M_A12TR u4520 ( .A(n3757), .B(n3758), .S0(n3883), .Y(n3892) );
  OA21A1OI2_X0P5M_A12TR u4521 ( .A0(rtgt[3]), .A1(n3753), .B0(n3754), .C0(
        n3883), .Y(n3890) );
  INV_X0P5B_A12TR u4522 ( .A(rsrc[3]), .Y(n3883) );
  AOI222_X0P5M_A12TR u4523 ( .A0(wsub[3]), .A1(n3762), .B0(n3759), .B1(rtgt[4]), .C0(n3760), .C1(rtgt[7]), .Y(n3888) );
  AOI222_X0P5M_A12TR u4524 ( .A0(wsubc[3]), .A1(n3761), .B0(wneg[3]), .B1(
        n3775), .C0(wadd[3]), .C1(n3763), .Y(n3887) );
  AOI22_X0P5M_A12TR u4525 ( .A0(waddc[3]), .A1(n3764), .B0(dwb_dat_o[3]), .B1(
        n3765), .Y(n3886) );
  OAI222_X0P5M_A12TR u4526 ( .A0(n3458), .A1(n3776), .B0(n3778), .B1(n3893), 
        .C0(qena[3]), .C1(n3894), .Y(n1849) );
  INV_X0P5B_A12TR u4527 ( .A(wpclat[2]), .Y(n3894) );
  OAI221_X0P5M_A12TR u4528 ( .A0(n3064), .A1(n3895), .B0(n3066), .B1(n3458), 
        .C0(n3896), .Y(n1847) );
  AOI22_X0P5M_A12TR u4529 ( .A0(n2748), .A1(n3069), .B0(n3871), .B1(wpclat[2]), 
        .Y(n3896) );
  INV_X0P5B_A12TR u4530 ( .A(wstkw[3]), .Y(n3895) );
  OAI211_X0P5M_A12TR u4531 ( .A0(qena[1]), .A1(n3893), .B0(n3897), .C0(n3898), 
        .Y(n1846) );
  AOI222_X0P5M_A12TR u4532 ( .A0(wpcinc[2]), .A1(n3792), .B0(n388), .B1(n3793), 
        .C0(n3794), .C1(wstkw[3]), .Y(n3898) );
  AOI22_X0P5M_A12TR u4533 ( .A0(n368), .A1(n3795), .B0(n3796), .B1(rireg[2]), 
        .Y(n3897) );
  INV_X0P5B_A12TR u4534 ( .A(rpcnxt[2]), .Y(n3893) );
  OAI211_X0P5M_A12TR u4535 ( .A0(qena[1]), .A1(n3899), .B0(n3900), .C0(n3901), 
        .Y(n1843) );
  AOI222_X0P5M_A12TR u4536 ( .A0(wpcinc[17]), .A1(n3792), .B0(n403), .B1(n3793), .C0(n3794), .C1(wstkw[18]), .Y(n3901) );
  AOI22_X0P5M_A12TR u4537 ( .A0(n383), .A1(n3795), .B0(n3796), .B1(rromlat[9]), 
        .Y(n3900) );
  OAI211_X0P5M_A12TR u4538 ( .A0(qena[1]), .A1(n3902), .B0(n3903), .C0(n3904), 
        .Y(n1840) );
  AOI222_X0P5M_A12TR u4539 ( .A0(wpcinc[13]), .A1(n3792), .B0(n399), .B1(n3793), .C0(n3794), .C1(wstkw[14]), .Y(n3904) );
  AOI22_X0P5M_A12TR u4540 ( .A0(n379), .A1(n3795), .B0(n3796), .B1(rromlat[5]), 
        .Y(n3903) );
  OAI222_X0P5M_A12TR u4541 ( .A0(n3905), .A1(n3776), .B0(n3902), .B1(n3778), 
        .C0(qena[3]), .C1(n3906), .Y(n1838) );
  INV_X0P5B_A12TR u4542 ( .A(rpcnxt[13]), .Y(n3902) );
  OAI221_X0P5M_A12TR u4543 ( .A0(n3907), .A1(n3908), .B0(n3468), .B1(n3909), 
        .C0(n3910), .Y(n1836) );
  AOI22_X0P5M_A12TR u4544 ( .A0(n2749), .A1(n3069), .B0(wpclat[13]), .B1(n3871), .Y(n3910) );
  INV_X0P5B_A12TR u4545 ( .A(wstkw[14]), .Y(n3908) );
  OAI221_X0P5M_A12TR u4546 ( .A0(n3911), .A1(n3737), .B0(n3738), .B1(n3912), 
        .C0(n3913), .Y(n1835) );
  AOI221_X0P5M_A12TR u4547 ( .A0(rmask[6]), .A1(n3741), .B0(n3742), .B1(n3914), 
        .C0(n3744), .Y(n3913) );
  NAND4_X0P5A_A12TR u4548 ( .A(n3915), .B(n3916), .C(n3917), .D(n3918), .Y(
        n1833) );
  AOI211_X0P5M_A12TR u4549 ( .A0(n3750), .A1(rtgt[5]), .B0(n3919), .C0(n3920), 
        .Y(n3918) );
  AOI21_X0P5M_A12TR u4550 ( .A0(n3921), .A1(n3754), .B0(n4429), .Y(n3920) );
  MXIT2_X0P5M_A12TR u4551 ( .A(n3757), .B(n3758), .S0(n3912), .Y(n3921) );
  OA21A1OI2_X0P5M_A12TR u4552 ( .A0(rtgt[6]), .A1(n3753), .B0(n3754), .C0(
        n3912), .Y(n3919) );
  INV_X0P5B_A12TR u4553 ( .A(rsrc[6]), .Y(n3912) );
  AOI222_X0P5M_A12TR u4554 ( .A0(wsub[6]), .A1(n3762), .B0(n3759), .B1(rtgt[7]), .C0(n3760), .C1(rtgt[2]), .Y(n3917) );
  AOI222_X0P5M_A12TR u4555 ( .A0(wsubc[6]), .A1(n3761), .B0(wneg[6]), .B1(
        n3775), .C0(wadd[6]), .C1(n3763), .Y(n3916) );
  AOI22_X0P5M_A12TR u4556 ( .A0(waddc[6]), .A1(n3764), .B0(dwb_dat_o[6]), .B1(
        n3765), .Y(n3915) );
  NAND4_X0P5A_A12TR u4557 ( .A(n3922), .B(n3923), .C(n3924), .D(n3925), .Y(
        n1831) );
  AOI222_X0P5M_A12TR u4558 ( .A0(wfsrplusw1[5]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[5]), .C0(n3815), .C1(wfsrinc2[5]), .Y(n3925) );
  AOI222_X0P5M_A12TR u4559 ( .A0(n3724), .A1(rfsr0l[5]), .B0(wfsrplusw2[5]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[5]), .Y(n3924) );
  AOI222_X0P5M_A12TR u4560 ( .A0(n3723), .A1(rfsr2l[5]), .B0(wfsrplusw0[5]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[5]), .Y(n3923) );
  AOI222_X0P5M_A12TR u4561 ( .A0(dwb_adr_o[5]), .A1(n3819), .B0(n3820), .B1(
        rromlat[5]), .C0(reaptr[5]), .C1(n3821), .Y(n3922) );
  MXIT2_X0P5M_A12TR u4562 ( .A(n3555), .B(n3067), .S0(n3926), .Y(n1829) );
  AND4_X0P5M_A12TR u4563 ( .A(n3646), .B(n3262), .C(n3263), .D(n3684), .Y(
        n3926) );
  NOR3_X0P5A_A12TR u4564 ( .A(dwb_adr_o[2]), .B(dwb_adr_o[3]), .C(n3734), .Y(
        n3262) );
  INV_X0P5B_A12TR u4565 ( .A(rswdten), .Y(n3555) );
  OAI221_X0P5M_A12TR u4566 ( .A0(n3927), .A1(n3928), .B0(n3242), .B1(n3735), 
        .C0(n3929), .Y(n1809) );
  INV_X0P5B_A12TR u4567 ( .A(dwb_stb_o), .Y(n3735) );
  AOI22_X0P5M_A12TR u4568 ( .A0(rmxsrc[0]), .A1(n3930), .B0(rmxtgt[0]), .B1(
        n3931), .Y(n3927) );
  MXIT2_X0P5M_A12TR u4569 ( .A(n3932), .B(n3074), .S0(n3933), .Y(n1807) );
  MXIT2_X0P5M_A12TR u4570 ( .A(n3074), .B(n3784), .S0(n3933), .Y(n1805) );
  MXIT2_X0P5M_A12TR u4571 ( .A(n3784), .B(n3375), .S0(n3933), .Y(n1803) );
  MXIT2_X0P5M_A12TR u4572 ( .A(n3375), .B(n3932), .S0(n3933), .Y(n1801) );
  XNOR2_X0P5M_A12TR u4573 ( .A(qfsm[0]), .B(n3933), .Y(n1799) );
  NAND2_X0P5A_A12TR u4574 ( .A(n3934), .B(n3238), .Y(n17971) );
  INV_X0P5B_A12TR u4575 ( .A(n3247), .Y(n3238) );
  MXIT2_X0P5M_A12TR u4576 ( .A(n3460), .B(qfsm[1]), .S0(n3933), .Y(n3934) );
  NAND3_X0P5A_A12TR u4577 ( .A(n3935), .B(n3054), .C(n3936), .Y(n3933) );
  XNOR2_X0P5M_A12TR u4578 ( .A(dwb_stb_o), .B(dwb_ack_i), .Y(n3936) );
  XNOR2_X0P5M_A12TR u4579 ( .A(iwb_stb_o), .B(iwb_ack_i), .Y(n3935) );
  OAI22_X0P5M_A12TR u4580 ( .A0(qena[3]), .A1(n3937), .B0(rromlat[11]), .B1(
        n3938), .Y(n17901) );
  MXT2_X0P5M_A12TR u4581 ( .A(rmxbcc[2]), .B(rromlat[10]), .S0(qena[3]), .Y(
        n17871) );
  MXT2_X0P5M_A12TR u4582 ( .A(rmxbcc[1]), .B(rromlat[9]), .S0(qena[3]), .Y(
        n17841) );
  MXT2_X0P5M_A12TR u4583 ( .A(rmask[4]), .B(n3939), .S0(n3940), .Y(n17821) );
  MXIT2_X0P5M_A12TR u4584 ( .A(n3941), .B(n3942), .S0(n3765), .Y(n1780) );
  NAND2_X0P5A_A12TR u4585 ( .A(n3943), .B(n3207), .Y(n3941) );
  MXIT2_X0P5M_A12TR u4586 ( .A(n3944), .B(n3945), .S0(n3765), .Y(n1778) );
  MXT2_X0P5M_A12TR u4587 ( .A(rmask[0]), .B(n3085), .S0(n3940), .Y(n1776) );
  OAI221_X0P5M_A12TR u4588 ( .A0(rromlat[9]), .A1(n3946), .B0(qena[3]), .B1(
        n3947), .C0(n3948), .Y(n1774) );
  AOI31_X0P5M_A12TR u4589 ( .A0(n3949), .A1(n3950), .A2(n3951), .B0(n3952), 
        .Y(n3948) );
  INV_X0P5B_A12TR u4590 ( .A(n3953), .Y(n3952) );
  AO21A1AI2_X0P5M_A12TR u4591 ( .A0(n3211), .A1(rromlat[13]), .B0(n3954), .C0(
        n3955), .Y(n3953) );
  INV_X0P5B_A12TR u4592 ( .A(rmxskp[1]), .Y(n3947) );
  MXT2_X0P5M_A12TR u4593 ( .A(rmask[5]), .B(n3956), .S0(n3940), .Y(n1772) );
  MXIT2_X0P5M_A12TR u4594 ( .A(n3957), .B(n3958), .S0(n3765), .Y(n1770) );
  NAND2_X0P5A_A12TR u4595 ( .A(n3943), .B(rromlat[9]), .Y(n3957) );
  MXIT2_X0P5M_A12TR u4596 ( .A(n3959), .B(n3960), .S0(n3765), .Y(n1768) );
  OAI211_X0P5M_A12TR u4597 ( .A0(n3213), .A1(n3961), .B0(n3946), .C0(n3962), 
        .Y(n1766) );
  AOI21_X0P5M_A12TR u4598 ( .A0(n3963), .A1(n3211), .B0(n3964), .Y(n3962) );
  MXIT2_X0P5M_A12TR u4599 ( .A(n3965), .B(n3710), .S0(n3074), .Y(n3964) );
  INV_X0P5B_A12TR u4600 ( .A(rmxskp[0]), .Y(n3710) );
  AO21A1AI2_X0P5M_A12TR u4601 ( .A0(n3954), .A1(rromlat[12]), .B0(n3966), .C0(
        n3967), .Y(n3965) );
  INV_X0P5B_A12TR u4602 ( .A(n3968), .Y(n3946) );
  INV_X0P5B_A12TR u4603 ( .A(n3969), .Y(n3961) );
  MXT2_X0P5M_A12TR u4604 ( .A(rmxbsr[1]), .B(n3970), .S0(qena[1]), .Y(n1764)
         );
  MXIT2_X0P5M_A12TR u4605 ( .A(n3971), .B(n3972), .S0(n3765), .Y(n1762) );
  NAND3_X0P5A_A12TR u4606 ( .A(n3973), .B(n3944), .C(n3974), .Y(n3971) );
  MXT2_X0P5M_A12TR u4607 ( .A(rmxbcc[0]), .B(rromlat[8]), .S0(qena[3]), .Y(
        n1759) );
  NAND3B_X0P5M_A12TR u4608 ( .AN(n3975), .B(n3976), .C(n3977), .Y(n1757) );
  AOI31_X0P5M_A12TR u4609 ( .A0(n3978), .A1(rromlat[14]), .A2(n3979), .B0(
        n3969), .Y(n3977) );
  MXIT2_X0P5M_A12TR u4610 ( .A(n3980), .B(rmxsrc[1]), .S0(n3074), .Y(n3976) );
  OAI211_X0P5M_A12TR u4611 ( .A0(n3981), .A1(n3982), .B0(n3983), .C0(n3984), 
        .Y(n1755) );
  AOI221_X0P5M_A12TR u4612 ( .A0(n3085), .A1(n3985), .B0(n3986), .B1(n3987), 
        .C0(n3988), .Y(n3984) );
  MXIT2_X0P5M_A12TR u4613 ( .A(n3980), .B(rmxsrc[0]), .S0(n3074), .Y(n3983) );
  NAND4_X0P5A_A12TR u4614 ( .A(n3989), .B(n3990), .C(n3991), .D(n3992), .Y(
        n3980) );
  AO21A1AI2_X0P5M_A12TR u4615 ( .A0(n3993), .A1(n3213), .B0(n3966), .C0(n3950), 
        .Y(n3991) );
  INV_X0P5B_A12TR u4616 ( .A(n3994), .Y(n3966) );
  AO21A1AI2_X0P5M_A12TR u4617 ( .A0(n3995), .A1(n3217), .B0(n3086), .C0(n3967), 
        .Y(n3990) );
  OAI31_X0P5M_A12TR u4618 ( .A0(n3996), .A1(n3939), .A2(n3997), .B0(n3998), 
        .Y(n3989) );
  NOR2_X0P5A_A12TR u4619 ( .A(n3207), .B(n3999), .Y(n3996) );
  OAI221_X0P5M_A12TR u4620 ( .A0(n4000), .A1(n3938), .B0(qena[3]), .B1(n4001), 
        .C0(n4002), .Y(n1753) );
  INV_X0P5B_A12TR u4621 ( .A(n4003), .Y(n4000) );
  MXIT2_X0P5M_A12TR u4622 ( .A(n4004), .B(n3406), .S0(n3375), .Y(n1751) );
  AOI32_X0P5M_A12TR u4623 ( .A0(rromlat[15]), .A1(n3213), .A2(n3993), .B0(
        rromlat[8]), .B1(n3970), .Y(n4004) );
  OAI211_X0P5M_A12TR u4624 ( .A0(rromlat[14]), .A1(n3219), .B0(n4005), .C0(
        n4006), .Y(n3970) );
  AOI211_X0P5M_A12TR u4625 ( .A0(n4007), .A1(n4008), .B0(n3995), .C0(n4009), 
        .Y(n4006) );
  AOI21B_X0P5M_A12TR u4626 ( .A0(n3974), .A1(n3076), .B0N(n3998), .Y(n4009) );
  NOR2_X0P5A_A12TR u4627 ( .A(n4010), .B(n3997), .Y(n3076) );
  OAI211_X0P5M_A12TR u4628 ( .A0(n3974), .A1(n4011), .B0(n4012), .C0(n4013), 
        .Y(n1749) );
  AOI21_X0P5M_A12TR u4629 ( .A0(rmxsta[0]), .A1(n3074), .B0(n4014), .Y(n4013)
         );
  NAND4_X0P5A_A12TR u4630 ( .A(n4012), .B(n4015), .C(n4016), .D(n4017), .Y(
        n1747) );
  AOI222_X0P5M_A12TR u4631 ( .A0(rmxsta[1]), .A1(n3074), .B0(n3978), .B1(n3215), .C0(n4010), .C1(n4018), .Y(n4017) );
  AOI32_X0P5M_A12TR u4632 ( .A0(n3987), .A1(n3219), .A2(n3951), .B0(n4019), 
        .B1(n3997), .Y(n4016) );
  INV_X0P5B_A12TR u4633 ( .A(n3974), .Y(n3987) );
  NAND2_X0P5A_A12TR u4634 ( .A(n3956), .B(n3985), .Y(n4012) );
  INV_X0P5B_A12TR u4635 ( .A(n4020), .Y(n1743) );
  AOI221_X0P5M_A12TR u4636 ( .A0(n3950), .A1(n4018), .B0(n3074), .B1(rmxtgt[1]), .C0(n3988), .Y(n4020) );
  NOR3_X0P5A_A12TR u4637 ( .A(n3213), .B(rromlat[13]), .C(n4021), .Y(n3988) );
  NAND4_X0P5A_A12TR u4638 ( .A(n4022), .B(n4023), .C(n4024), .D(n4025), .Y(
        n1741) );
  AOI221_X0P5M_A12TR u4639 ( .A0(n4018), .A1(n3950), .B0(n3951), .B1(n3213), 
        .C0(n4026), .Y(n4025) );
  AO21A1AI2_X0P5M_A12TR u4640 ( .A0(n3999), .A1(n3959), .B0(n4027), .C0(n4028), 
        .Y(n4026) );
  NOR2_X0P5A_A12TR u4641 ( .A(n3969), .B(n4029), .Y(n4028) );
  AOI21_X0P5M_A12TR u4642 ( .A0(rmxtgt[0]), .A1(n3074), .B0(n3975), .Y(n4024)
         );
  OR6_X0P5M_A12TR u4643 ( .A(n4030), .B(n3968), .C(n3969), .D(n4031), .E(n4032), .F(n4033), .Y(n1739) );
  NAND4_X0P5A_A12TR u4644 ( .A(n4034), .B(n4022), .C(n4035), .D(n4036), .Y(
        n4033) );
  AOI22_X0P5M_A12TR u4645 ( .A0(n4019), .A1(n3956), .B0(n4037), .B1(n4010), 
        .Y(n4036) );
  NOR2_X0P5A_A12TR u4646 ( .A(n3973), .B(n3207), .Y(n3956) );
  AOI22_X0P5M_A12TR u4647 ( .A0(n3997), .A1(n3985), .B0(n4038), .B1(n4018), 
        .Y(n4035) );
  INV_X0P5B_A12TR u4648 ( .A(n3075), .Y(n4018) );
  NOR2B_X0P5M_A12TR u4649 ( .AN(n4039), .B(n4040), .Y(n4022) );
  OAI211_X0P5M_A12TR u4650 ( .A0(n3979), .A1(n4010), .B0(n3219), .C0(n3951), 
        .Y(n4039) );
  AOI22_X0P5M_A12TR u4651 ( .A0(n3993), .A1(n3955), .B0(rmxalu[1]), .B1(n3074), 
        .Y(n4034) );
  AO21A1AI2_X0P5M_A12TR u4652 ( .A0(n4021), .A1(n4041), .B0(n3213), .C0(n4042), 
        .Y(n4032) );
  OA21A1OI2_X0P5M_A12TR u4653 ( .A0(n3986), .A1(n3079), .B0(n3967), .C0(n4043), 
        .Y(n4042) );
  NOR3_X0P5A_A12TR u4654 ( .A(n3999), .B(rromlat[13]), .C(n4044), .Y(n4043) );
  OAI211_X0P5M_A12TR u4655 ( .A0(n3979), .A1(n3950), .B0(qena[3]), .C0(n3954), 
        .Y(n4041) );
  NOR2_X0P5A_A12TR u4656 ( .A(n4021), .B(n3215), .Y(n3969) );
  INV_X0P5B_A12TR u4657 ( .A(n4045), .Y(n4021) );
  NOR2_X0P5A_A12TR u4658 ( .A(n4027), .B(n3974), .Y(n3968) );
  MXT2_X0P5M_A12TR u4659 ( .A(reaptr[7]), .B(rromlat[7]), .S0(n3398), .Y(n1736) );
  MXT2_X0P5M_A12TR u4660 ( .A(reaptr[6]), .B(rromlat[6]), .S0(n3398), .Y(n1733) );
  INV_X0P5B_A12TR u4661 ( .A(n3389), .Y(n3398) );
  MXIT2_X0P5M_A12TR u4662 ( .A(n3201), .B(n4046), .S0(n3389), .Y(n1730) );
  MXIT2_X0P5M_A12TR u4663 ( .A(n3199), .B(n4047), .S0(n3389), .Y(n1727) );
  MXIT2_X0P5M_A12TR u4664 ( .A(n3197), .B(n4048), .S0(n3389), .Y(n1724) );
  OAI21_X0P5M_A12TR u4665 ( .A0(qena[3]), .A1(n3616), .B0(n4049), .Y(n1722) );
  MXIT2_X0P5M_A12TR u4666 ( .A(n3084), .B(n4050), .S0(n3389), .Y(n1719) );
  OAI22_X0P5M_A12TR u4667 ( .A0(qena[3]), .A1(n4051), .B0(n3084), .B1(n4049), 
        .Y(n1717) );
  OAI211_X0P5M_A12TR u4668 ( .A0(qena[3]), .A1(n3714), .B0(n4002), .C0(n4052), 
        .Y(n1715) );
  INV_X0P5B_A12TR u4669 ( .A(rmxskp[2]), .Y(n3714) );
  OAI21_X0P5M_A12TR u4670 ( .A0(qena[3]), .A1(n4053), .B0(n4052), .Y(n1713) );
  AOI222_X0P5M_A12TR u4671 ( .A0(n3079), .A1(n4038), .B0(n4003), .B1(n3963), 
        .C0(qena[3]), .C1(n4054), .Y(n4052) );
  OAI211_X0P5M_A12TR u4672 ( .A0(n3078), .A1(n3205), .B0(n3944), .C0(
        rromlat[11]), .Y(n4003) );
  MXIT2_X0P5M_A12TR u4673 ( .A(n3083), .B(n4055), .S0(n3389), .Y(n1710) );
  OAI22_X0P5M_A12TR u4674 ( .A0(qena[3]), .A1(n3617), .B0(n3083), .B1(n4049), 
        .Y(n1708) );
  MXIT2_X0P5M_A12TR u4675 ( .A(n3192), .B(n4056), .S0(n3389), .Y(n1705) );
  OAI21_X0P5M_A12TR u4676 ( .A0(rmxbsr[1]), .A1(rmxbsr[0]), .B0(qena[2]), .Y(
        n3389) );
  OAI22_X0P5M_A12TR u4677 ( .A0(qena[3]), .A1(n3618), .B0(n3192), .B1(n4049), 
        .Y(n1703) );
  NAND4_X0P5A_A12TR u4678 ( .A(n4057), .B(rromlat[3]), .C(n3079), .D(n3199), 
        .Y(n4049) );
  INV_X0P5B_A12TR u4679 ( .A(n4058), .Y(n1701) );
  AOI211_X0P5M_A12TR u4680 ( .A0(n3074), .A1(rmxsta[2]), .B0(n4059), .C0(n4014), .Y(n4058) );
  NAND4_X0P5A_A12TR u4681 ( .A(n4060), .B(n4061), .C(n4062), .D(n4015), .Y(
        n4014) );
  NAND2_X0P5A_A12TR u4682 ( .A(n4019), .B(n3997), .Y(n4060) );
  NAND4_X0P5A_A12TR u4683 ( .A(n4063), .B(n4064), .C(n4065), .D(n3072), .Y(
        n1699) );
  AOI221_X0P5M_A12TR u4684 ( .A0(n3215), .A1(n4045), .B0(n3950), .B1(n3985), 
        .C0(n3975), .Y(n3072) );
  OAI22_X0P5M_A12TR u4685 ( .A0(rromlat[13]), .A1(n3981), .B0(n4044), .B1(
        n4066), .Y(n3975) );
  NOR3_X0P5A_A12TR u4686 ( .A(n3074), .B(rromlat[14]), .C(n3219), .Y(n4045) );
  AOI21_X0P5M_A12TR u4687 ( .A0(n4019), .A1(n4038), .B0(n4031), .Y(n4065) );
  AND4_X0P5M_A12TR u4688 ( .A(n3997), .B(n3955), .C(rromlat[14]), .D(n3205), 
        .Y(n4031) );
  MXIT2_X0P5M_A12TR u4689 ( .A(n4067), .B(rmxdst[0]), .S0(n3074), .Y(n4063) );
  NOR2_X0P5A_A12TR u4690 ( .A(n4005), .B(n3207), .Y(n4067) );
  INV_X0P5B_A12TR u4691 ( .A(n3073), .Y(n4005) );
  NAND3_X0P5A_A12TR u4692 ( .A(n3992), .B(n3994), .C(n4068), .Y(n3073) );
  OAI211_X0P5M_A12TR u4693 ( .A0(rromlat[12]), .A1(rromlat[14]), .B0(n4066), 
        .C0(n3219), .Y(n4068) );
  OAI211_X0P5M_A12TR u4694 ( .A0(qena[3]), .A1(n4069), .B0(n4070), .C0(n4071), 
        .Y(n1697) );
  OA21A1OI2_X0P5M_A12TR u4695 ( .A0(n3985), .A1(n4019), .B0(n4038), .C0(n4072), 
        .Y(n4071) );
  NOR2_X0P5A_A12TR u4696 ( .A(n3974), .B(n4073), .Y(n4072) );
  NAND4B_X0P5M_A12TR u4697 ( .AN(n4074), .B(n4075), .C(n4076), .D(n4077), .Y(
        n1695) );
  NOR3_X0P5A_A12TR u4698 ( .A(n4030), .B(n4029), .C(n4037), .Y(n4077) );
  INV_X0P5B_A12TR u4699 ( .A(n4015), .Y(n4029) );
  OAI31_X0P5M_A12TR u4700 ( .A0(n4078), .A1(n4079), .A2(n4080), .B0(qena[3]), 
        .Y(n4015) );
  NOR3_X0P5A_A12TR u4701 ( .A(n3982), .B(n4081), .C(n3078), .Y(n4080) );
  INV_X0P5B_A12TR u4702 ( .A(n3992), .Y(n4079) );
  NAND2_X0P5A_A12TR u4703 ( .A(n3943), .B(n4008), .Y(n3992) );
  AO21A1AI2_X0P5M_A12TR u4704 ( .A0(n3974), .A1(n3973), .B0(n3994), .C0(n4082), 
        .Y(n4078) );
  NAND2_X0P5A_A12TR u4705 ( .A(n4038), .B(n3998), .Y(n4082) );
  NOR2_X0P5A_A12TR u4706 ( .A(n3943), .B(n3979), .Y(n3974) );
  INV_X0P5B_A12TR u4707 ( .A(n4062), .Y(n4030) );
  NAND2_X0P5A_A12TR u4708 ( .A(n3939), .B(n3079), .Y(n4062) );
  NOR2_X0P5A_A12TR u4709 ( .A(n3075), .B(rromlat[8]), .Y(n3079) );
  AOI32_X0P5M_A12TR u4710 ( .A0(n4010), .A1(n3219), .A2(n3951), .B0(n3943), 
        .B1(n4083), .Y(n4076) );
  AO21_X0P5M_A12TR u4711 ( .A0(n3207), .A1(n3985), .B0(n3986), .Y(n4083) );
  AOI22_X0P5M_A12TR u4712 ( .A0(n3967), .A1(n4084), .B0(n3979), .B1(n3985), 
        .Y(n4075) );
  NAND2B_X0P5M_A12TR u4713 ( .AN(n4019), .B(n4073), .Y(n4084) );
  AOI21_X0P5M_A12TR u4714 ( .A0(n3949), .A1(n3951), .B0(n4085), .Y(n4073) );
  OAI21_X0P5M_A12TR u4715 ( .A0(n4086), .A1(qena[3]), .B0(n4070), .Y(n4074) );
  AOI31_X0P5M_A12TR u4716 ( .A0(n3997), .A1(n3205), .A2(n3963), .B0(n4087), 
        .Y(n4070) );
  INV_X0P5B_A12TR u4717 ( .A(n4064), .Y(n4087) );
  AOI211_X0P5M_A12TR u4718 ( .A0(n3979), .A1(n4019), .B0(n4059), .C0(n4040), 
        .Y(n4064) );
  NOR2_X0P5A_A12TR u4719 ( .A(n3207), .B(n3078), .Y(n3997) );
  NAND4_X0P5A_A12TR u4720 ( .A(n4088), .B(n4089), .C(n4090), .D(n4091), .Y(
        n1693) );
  NOR3_X0P5A_A12TR u4721 ( .A(n4092), .B(n4040), .C(n4059), .Y(n4091) );
  NOR3_X0P5A_A12TR u4722 ( .A(n4093), .B(n3083), .C(n4094), .Y(n4059) );
  NOR2_X0P5A_A12TR u4723 ( .A(n3959), .B(n3075), .Y(n4040) );
  INV_X0P5B_A12TR u4724 ( .A(n4007), .Y(n3959) );
  NOR2_X0P5A_A12TR u4725 ( .A(n4095), .B(n3207), .Y(n4007) );
  INV_X0P5B_A12TR u4726 ( .A(n4061), .Y(n4092) );
  NAND2_X0P5A_A12TR u4727 ( .A(n3986), .B(n4096), .Y(n4061) );
  NOR2_X0P5A_A12TR u4728 ( .A(n3982), .B(n4044), .Y(n3986) );
  INV_X0P5B_A12TR u4729 ( .A(n3978), .Y(n4044) );
  AOI31_X0P5M_A12TR u4730 ( .A0(n3950), .A1(n3207), .A2(n4019), .B0(n4097), 
        .Y(n4090) );
  NOR3_X0P5A_A12TR u4731 ( .A(n3981), .B(rromlat[14]), .C(rromlat[13]), .Y(
        n4097) );
  NOR2_X0P5A_A12TR u4732 ( .A(n3205), .B(n3075), .Y(n4019) );
  NAND2_X0P5A_A12TR u4733 ( .A(n4008), .B(qena[3]), .Y(n3075) );
  INV_X0P5B_A12TR u4734 ( .A(rromlat[9]), .Y(n3207) );
  NAND2_X0P5A_A12TR u4735 ( .A(n3973), .B(n3078), .Y(n3950) );
  AOI22_X0P5M_A12TR u4736 ( .A0(n4085), .A1(n4096), .B0(n3979), .B1(n4098), 
        .Y(n4089) );
  INV_X0P5B_A12TR u4737 ( .A(n4023), .Y(n4098) );
  AOI21_X0P5M_A12TR u4738 ( .A0(n3217), .A1(n3978), .B0(n4037), .Y(n4023) );
  NOR2_X0P5A_A12TR u4739 ( .A(n3994), .B(n3074), .Y(n4037) );
  NAND2_X0P5A_A12TR u4740 ( .A(n3954), .B(n3949), .Y(n3994) );
  NAND2_X0P5A_A12TR u4741 ( .A(n3973), .B(n3999), .Y(n4096) );
  INV_X0P5B_A12TR u4742 ( .A(n3943), .Y(n3999) );
  NOR2_X0P5A_A12TR u4743 ( .A(n3209), .B(rromlat[11]), .Y(n3943) );
  INV_X0P5B_A12TR u4744 ( .A(n4011), .Y(n4085) );
  NAND2_X0P5A_A12TR u4745 ( .A(n3954), .B(n3978), .Y(n4011) );
  NOR2_X0P5A_A12TR u4746 ( .A(n3074), .B(n4081), .Y(n3978) );
  INV_X0P5B_A12TR u4747 ( .A(n3995), .Y(n4081) );
  NOR2_X0P5A_A12TR u4748 ( .A(n3213), .B(rromlat[15]), .Y(n3995) );
  INV_X0P5B_A12TR u4749 ( .A(rromlat[12]), .Y(n3213) );
  NOR2_X0P5A_A12TR u4750 ( .A(n3215), .B(rromlat[14]), .Y(n3954) );
  AOI22_X0P5M_A12TR u4751 ( .A0(n3939), .A1(n3985), .B0(rmxalu[0]), .B1(n3074), 
        .Y(n4088) );
  INV_X0P5B_A12TR u4752 ( .A(n4027), .Y(n3985) );
  NAND2_X0P5A_A12TR u4753 ( .A(n3998), .B(qena[3]), .Y(n4027) );
  NOR2B_X0P5M_A12TR u4754 ( .AN(n3949), .B(n4066), .Y(n3998) );
  NOR2_X0P5A_A12TR u4755 ( .A(n3973), .B(rromlat[9]), .Y(n3939) );
  INV_X0P5B_A12TR u4756 ( .A(n4010), .Y(n3973) );
  NOR2_X0P5A_A12TR u4757 ( .A(n3211), .B(rromlat[10]), .Y(n4010) );
  OAI31_X0P5M_A12TR u4758 ( .A0(n4099), .A1(n4100), .A2(n4093), .B0(n4101), 
        .Y(n1691) );
  NAND2_X0P5A_A12TR u4759 ( .A(rsleep_), .B(n3074), .Y(n4101) );
  NAND3_X0P5A_A12TR u4760 ( .A(n3084), .B(n3199), .C(rromlat[1]), .Y(n4099) );
  OAI31_X0P5M_A12TR u4761 ( .A0(n3944), .A1(n3205), .A2(n3938), .B0(n4102), 
        .Y(n1684) );
  MXIT2_X0P5M_A12TR u4762 ( .A(n4103), .B(rmxsha[1]), .S0(n3074), .Y(n4102) );
  AOI31_X0P5M_A12TR u4763 ( .A0(n4038), .A1(rromlat[15]), .A2(n4104), .B0(
        n4105), .Y(n4103) );
  NOR2_X0P5A_A12TR u4764 ( .A(rromlat[12]), .B(n4066), .Y(n4104) );
  INV_X0P5B_A12TR u4765 ( .A(n3963), .Y(n3938) );
  INV_X0P5B_A12TR u4766 ( .A(n4038), .Y(n3944) );
  OAI31_X0P5M_A12TR u4767 ( .A0(n4093), .A1(n4106), .A2(n3624), .B0(n4107), 
        .Y(n1682) );
  NAND2_X0P5A_A12TR u4768 ( .A(rmxsha[0]), .B(n3074), .Y(n4107) );
  INV_X0P5B_A12TR u4769 ( .A(n4054), .Y(n4106) );
  INV_X0P5B_A12TR u4770 ( .A(n4108), .Y(n4093) );
  MXT2_X0P5M_A12TR u4771 ( .A(rmxstk[0]), .B(n4109), .S0(qena[3]), .Y(n1680)
         );
  AO21A1AI2_X0P5M_A12TR u4772 ( .A0(n4110), .A1(n4111), .B0(n4109), .C0(n4112), 
        .Y(n1678) );
  NAND2_X0P5A_A12TR u4773 ( .A(rmxstk[1]), .B(n3074), .Y(n4112) );
  OAI31_X0P5M_A12TR u4774 ( .A0(n4094), .A1(rromlat[0]), .A2(n3083), .B0(n4113), .Y(n4109) );
  AOI21_X0P5M_A12TR u4775 ( .A0(n4038), .A1(n3086), .B0(n4054), .Y(n4113) );
  NOR3_X0P5A_A12TR u4776 ( .A(n3199), .B(rromlat[2]), .C(n4100), .Y(n4054) );
  INV_X0P5B_A12TR u4777 ( .A(rromlat[4]), .Y(n3199) );
  INV_X0P5B_A12TR u4778 ( .A(n4114), .Y(n4094) );
  AOI32_X0P5M_A12TR u4779 ( .A0(n4108), .A1(n3083), .A2(n4114), .B0(n4115), 
        .B1(rromlat[11]), .Y(n4111) );
  INV_X0P5B_A12TR u4780 ( .A(n4002), .Y(n4115) );
  NAND3_X0P5A_A12TR u4781 ( .A(rromlat[15]), .B(rromlat[12]), .C(n3951), .Y(
        n4002) );
  NOR2_X0P5A_A12TR u4782 ( .A(n3982), .B(n3074), .Y(n3951) );
  INV_X0P5B_A12TR u4783 ( .A(n3993), .Y(n3982) );
  NOR2_X0P5A_A12TR u4784 ( .A(n3217), .B(rromlat[13]), .Y(n3993) );
  NOR2_X0P5A_A12TR u4785 ( .A(n3192), .B(n3074), .Y(n4108) );
  AOI22_X0P5M_A12TR u4786 ( .A0(qena[3]), .A1(n3624), .B0(n4038), .B1(n3963), 
        .Y(n4110) );
  NOR2_X0P5A_A12TR u4787 ( .A(n3981), .B(n4066), .Y(n3963) );
  NAND2_X0P5A_A12TR u4788 ( .A(rromlat[14]), .B(rromlat[13]), .Y(n4066) );
  INV_X0P5B_A12TR u4789 ( .A(n3955), .Y(n3981) );
  NOR3_X0P5A_A12TR u4790 ( .A(n3074), .B(rromlat[12]), .C(n3219), .Y(n3955) );
  INV_X0P5B_A12TR u4791 ( .A(rromlat[15]), .Y(n3219) );
  NOR2_X0P5A_A12TR u4792 ( .A(n3078), .B(rromlat[9]), .Y(n4038) );
  INV_X0P5B_A12TR u4793 ( .A(n3967), .Y(n3078) );
  NOR2_X0P5A_A12TR u4794 ( .A(n3211), .B(n3209), .Y(n3967) );
  INV_X0P5B_A12TR u4795 ( .A(rromlat[10]), .Y(n3209) );
  INV_X0P5B_A12TR u4796 ( .A(rromlat[11]), .Y(n3211) );
  INV_X0P5B_A12TR u4797 ( .A(n4105), .Y(n3624) );
  XNOR2_X0P5M_A12TR u4798 ( .A(rintf[0]), .B(rintf[1]), .Y(n4105) );
  MXIT2_X0P5M_A12TR u4799 ( .A(n4116), .B(n4117), .S0(n3074), .Y(n1676) );
  NAND3_X0P5A_A12TR u4800 ( .A(n3192), .B(n3083), .C(n4114), .Y(n4116) );
  NOR3_X0P5A_A12TR u4801 ( .A(n3084), .B(rromlat[4]), .C(n4100), .Y(n4114) );
  NAND3_X0P5A_A12TR u4802 ( .A(n3086), .B(n3197), .C(n4057), .Y(n4100) );
  AND4_X0P5M_A12TR u4803 ( .A(n3085), .B(n3201), .C(n3088), .D(n3089), .Y(
        n4057) );
  INV_X0P5B_A12TR u4804 ( .A(rromlat[7]), .Y(n3089) );
  INV_X0P5B_A12TR u4805 ( .A(rromlat[6]), .Y(n3088) );
  INV_X0P5B_A12TR u4806 ( .A(rromlat[5]), .Y(n3201) );
  NOR2_X0P5A_A12TR u4807 ( .A(n4095), .B(rromlat[9]), .Y(n3085) );
  INV_X0P5B_A12TR u4808 ( .A(n3979), .Y(n4095) );
  NOR2_X0P5A_A12TR u4809 ( .A(rromlat[10]), .B(rromlat[11]), .Y(n3979) );
  INV_X0P5B_A12TR u4810 ( .A(rromlat[3]), .Y(n3197) );
  AND2_X0P5M_A12TR u4811 ( .A(n4008), .B(n3205), .Y(n3086) );
  INV_X0P5B_A12TR u4812 ( .A(rromlat[8]), .Y(n3205) );
  AND3_X0P5M_A12TR u4813 ( .A(n3215), .B(n3217), .C(n3949), .Y(n4008) );
  NOR2_X0P5A_A12TR u4814 ( .A(rromlat[12]), .B(rromlat[15]), .Y(n3949) );
  INV_X0P5B_A12TR u4815 ( .A(rromlat[14]), .Y(n3217) );
  INV_X0P5B_A12TR u4816 ( .A(rromlat[13]), .Y(n3215) );
  INV_X0P5B_A12TR u4817 ( .A(rromlat[2]), .Y(n3084) );
  INV_X0P5B_A12TR u4818 ( .A(rromlat[1]), .Y(n3083) );
  INV_X0P5B_A12TR u4819 ( .A(rromlat[0]), .Y(n3192) );
  OAI21_X0P5M_A12TR u4820 ( .A0(n3242), .A1(n4118), .B0(n3929), .Y(n1662) );
  NAND4_X0P5A_A12TR u4821 ( .A(rmxdst[0]), .B(n3247), .C(rmxdst[1]), .D(n3242), 
        .Y(n3929) );
  NOR2_X0P5A_A12TR u4822 ( .A(n4119), .B(qfsm[0]), .Y(n3247) );
  AO1B2_X0P5M_A12TR u4823 ( .B0(iwb_we_o), .B1(n3221), .A0N(n4120), .Y(n1660)
         );
  NAND4_X0P5A_A12TR u4824 ( .A(rmxtbl[2]), .B(rmxtbl[3]), .C(n3460), .D(n3242), 
        .Y(n4120) );
  MXIT2_X0P5M_A12TR u4825 ( .A(n4121), .B(n4122), .S0(n3054), .Y(n1658) );
  AOI31_X0P5M_A12TR u4826 ( .A0(rnskp), .A1(n3706), .A2(qfsm[0]), .B0(n3472), 
        .Y(n4122) );
  NAND4_X0P5A_A12TR u4827 ( .A(n3618), .B(n3617), .C(n4051), .D(n3616), .Y(
        n3706) );
  INV_X0P5B_A12TR u4828 ( .A(rmxtbl[3]), .Y(n3616) );
  INV_X0P5B_A12TR u4829 ( .A(rmxtbl[1]), .Y(n3617) );
  INV_X0P5B_A12TR u4830 ( .A(rmxtbl[0]), .Y(n3618) );
  INV_X0P5B_A12TR u4831 ( .A(iwb_stb_o), .Y(n4121) );
  MXIT2_X0P5M_A12TR u4832 ( .A(n214), .B(n3381), .S0(n3784), .Y(n1656) );
  INV_X0P5B_A12TR u4833 ( .A(rstkptr_[0]), .Y(n3381) );
  MXIT2_X0P5M_A12TR u4834 ( .A(n3851), .B(n3382), .S0(n3784), .Y(n1655) );
  INV_X0P5B_A12TR u4835 ( .A(rstkptr_[1]), .Y(n3382) );
  MXIT2_X0P5M_A12TR u4836 ( .A(n3853), .B(n3383), .S0(n3784), .Y(n1654) );
  INV_X0P5B_A12TR u4837 ( .A(rstkptr_[2]), .Y(n3383) );
  INV_X0P5B_A12TR u4838 ( .A(wstkinc[2]), .Y(n3853) );
  MXIT2_X0P5M_A12TR u4839 ( .A(n4123), .B(n3377), .S0(n3784), .Y(n1653) );
  INV_X0P5B_A12TR u4840 ( .A(rstkptr_[3]), .Y(n3377) );
  MXIT2_X0P5M_A12TR u4841 ( .A(n4124), .B(n3379), .S0(n3784), .Y(n1652) );
  INV_X0P5B_A12TR u4842 ( .A(qena[0]), .Y(n3784) );
  INV_X0P5B_A12TR u4843 ( .A(rstkptr_[4]), .Y(n3379) );
  OAI221_X0P5M_A12TR u4844 ( .A0(n3844), .A1(n4123), .B0(n3458), .B1(n3843), 
        .C0(n4125), .Y(n1651) );
  AOI22_X0P5M_A12TR u4845 ( .A0(n217), .A1(n3840), .B0(wstkdec[3]), .B1(n3855), 
        .Y(n4125) );
  INV_X0P5B_A12TR u4846 ( .A(wstkinc[3]), .Y(n4123) );
  OAI221_X0P5M_A12TR u4847 ( .A0(n3844), .A1(n4124), .B0(n3148), .B1(n3843), 
        .C0(n4126), .Y(n1650) );
  AOI22_X0P5M_A12TR u4848 ( .A0(n218), .A1(n3840), .B0(wstkdec[4]), .B1(n3855), 
        .Y(n4126) );
  INV_X0P5B_A12TR u4849 ( .A(wstkinc[4]), .Y(n4124) );
  OAI22_X0P5M_A12TR u4850 ( .A0(n3148), .A1(n3880), .B0(n3879), .B1(n3167), 
        .Y(n1649) );
  INV_X0P5B_A12TR u4851 ( .A(rtosu[4]), .Y(n3167) );
  OAI22_X0P5M_A12TR u4852 ( .A0(n3468), .A1(n3880), .B0(n3879), .B1(n3323), 
        .Y(n1648) );
  INV_X0P5B_A12TR u4853 ( .A(rtosu[6]), .Y(n3323) );
  OAI22_X0P5M_A12TR u4854 ( .A0(n3470), .A1(n3880), .B0(n3879), .B1(n3097), 
        .Y(n1647) );
  INV_X0P5B_A12TR u4855 ( .A(rtosu[7]), .Y(n3097) );
  MXIT2_X0P5M_A12TR u4856 ( .A(n3182), .B(n3179), .S0(n4127), .Y(n1646) );
  INV_X0P5B_A12TR u4857 ( .A(wrrc_7_), .Y(n3179) );
  INV_X0P5B_A12TR u4858 ( .A(rstatus_[0]), .Y(n3182) );
  MXT2_X0P5M_A12TR u4859 ( .A(rstatus_[3]), .B(rov), .S0(n4127), .Y(n1645) );
  MXT2_X0P5M_A12TR u4860 ( .A(rmxstal[2]), .B(rmxsta[2]), .S0(qena[3]), .Y(
        n1644) );
  MXT2_X0P5M_A12TR u4861 ( .A(rmxstal[0]), .B(rmxsta[0]), .S0(qena[3]), .Y(
        n1642) );
  MXT2_X0P5M_A12TR u4862 ( .A(rmxstal[1]), .B(rmxsta[1]), .S0(qena[3]), .Y(
        n1640) );
  OAI222_X0P5M_A12TR u4863 ( .A0(n3466), .A1(n3776), .B0(n4128), .B1(n3778), 
        .C0(qena[3]), .C1(n3663), .Y(n1638) );
  INV_X0P5B_A12TR u4864 ( .A(wpclat[4]), .Y(n3663) );
  INV_X0P5B_A12TR u4865 ( .A(rpcnxt[4]), .Y(n4128) );
  OAI221_X0P5M_A12TR u4866 ( .A0(n4129), .A1(n3737), .B0(n3738), .B1(n4130), 
        .C0(n4131), .Y(n1636) );
  AOI221_X0P5M_A12TR u4867 ( .A0(rmask[5]), .A1(n3741), .B0(n3742), .B1(n4132), 
        .C0(n3744), .Y(n4131) );
  AND2_X0P5M_A12TR u4868 ( .A(n3742), .B(rmxsrc[1]), .Y(n3744) );
  AND2_X0P5M_A12TR u4869 ( .A(rmxsrc[0]), .B(n3738), .Y(n3742) );
  AND2_X0P5M_A12TR u4870 ( .A(n3738), .B(rmxsrc[1]), .Y(n3741) );
  NAND3B_X0P5M_A12TR u4871 ( .AN(rmxsrc[0]), .B(n3930), .C(n3738), .Y(n3737)
         );
  INV_X0P5B_A12TR u4872 ( .A(rmxsrc[1]), .Y(n3930) );
  NAND4_X0P5A_A12TR u4873 ( .A(n4133), .B(n4134), .C(n4135), .D(n4136), .Y(
        n1634) );
  AOI211_X0P5M_A12TR u4874 ( .A0(n3750), .A1(rtgt[4]), .B0(n4137), .C0(n4138), 
        .Y(n4136) );
  AOI21_X0P5M_A12TR u4875 ( .A0(n4139), .A1(n3754), .B0(n4428), .Y(n4138) );
  MXIT2_X0P5M_A12TR u4876 ( .A(n3757), .B(n3758), .S0(n4130), .Y(n4139) );
  INV_X0P5B_A12TR u4877 ( .A(n3753), .Y(n3758) );
  AND3_X0P5M_A12TR u4878 ( .A(n3550), .B(n4086), .C(n4140), .Y(n3757) );
  OA21A1OI2_X0P5M_A12TR u4879 ( .A0(rtgt[5]), .A1(n3753), .B0(n3754), .C0(
        n4130), .Y(n4137) );
  INV_X0P5B_A12TR u4880 ( .A(rsrc[5]), .Y(n4130) );
  NAND4_X0P5A_A12TR u4881 ( .A(n4141), .B(rmxalu[0]), .C(n4142), .D(n4086), 
        .Y(n3754) );
  NAND3_X0P5A_A12TR u4882 ( .A(n3940), .B(n4143), .C(n4144), .Y(n3753) );
  MXIT2_X0P5M_A12TR u4883 ( .A(n4086), .B(n4145), .S0(n4069), .Y(n4144) );
  NAND2_X0P5A_A12TR u4884 ( .A(n4142), .B(n3550), .Y(n4145) );
  AOI222_X0P5M_A12TR u4885 ( .A0(wsub[5]), .A1(n3762), .B0(n3759), .B1(rtgt[6]), .C0(n3760), .C1(rtgt[1]), .Y(n4135) );
  AND3_X0P5M_A12TR u4886 ( .A(rmxalu[0]), .B(n4086), .C(n4140), .Y(n3760) );
  INV_X0P5B_A12TR u4887 ( .A(n4146), .Y(n3762) );
  AOI222_X0P5M_A12TR u4888 ( .A0(wsubc[5]), .A1(n3761), .B0(wneg[5]), .B1(
        n3775), .C0(wadd[5]), .C1(n3763), .Y(n4134) );
  INV_X0P5B_A12TR u4889 ( .A(n4147), .Y(n3761) );
  AOI22_X0P5M_A12TR u4890 ( .A0(waddc[5]), .A1(n3764), .B0(dwb_dat_o[5]), .B1(
        n3765), .Y(n4133) );
  OAI22_X0P5M_A12TR u4891 ( .A0(n3466), .A1(n3880), .B0(n3879), .B1(n3664), 
        .Y(n1632) );
  INV_X0P5B_A12TR u4892 ( .A(rtosu[5]), .Y(n3664) );
  NAND4_X0P5A_A12TR u4893 ( .A(n4148), .B(n4149), .C(n4150), .D(n4151), .Y(
        n1631) );
  AOI222_X0P5M_A12TR u4894 ( .A0(wfsrplusw1[3]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[3]), .C0(n3815), .C1(wfsrinc2[3]), .Y(n4151) );
  AOI222_X0P5M_A12TR u4895 ( .A0(n3724), .A1(rfsr0l[3]), .B0(wfsrplusw2[3]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[3]), .Y(n4150) );
  AOI222_X0P5M_A12TR u4896 ( .A0(n3723), .A1(rfsr2l[3]), .B0(wfsrplusw0[3]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[3]), .Y(n4149) );
  AOI222_X0P5M_A12TR u4897 ( .A0(dwb_adr_o[3]), .A1(n3819), .B0(n3820), .B1(
        rromlat[3]), .C0(reaptr[3]), .C1(n3821), .Y(n4148) );
  OAI221_X0P5M_A12TR u4898 ( .A0(n3235), .A1(n4152), .B0(n3404), .B1(n4153), 
        .C0(n4154), .Y(n1629) );
  AOI22_X0P5M_A12TR u4899 ( .A0(rbsr_[7]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[7]), .Y(n4154) );
  INV_X0P5B_A12TR u4900 ( .A(wfilebsr[15]), .Y(n3404) );
  INV_X0P5B_A12TR u4901 ( .A(rireg[7]), .Y(n3235) );
  MXT2_X0P5M_A12TR u4902 ( .A(rbsr_[7]), .B(wfilebsr[15]), .S0(n4127), .Y(
        n1628) );
  OAI221_X0P5M_A12TR u4903 ( .A0(n3234), .A1(n4152), .B0(n3402), .B1(n4153), 
        .C0(n4157), .Y(n1626) );
  AOI22_X0P5M_A12TR u4904 ( .A0(rbsr_[6]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[6]), .Y(n4157) );
  INV_X0P5B_A12TR u4905 ( .A(wfilebsr[14]), .Y(n3402) );
  INV_X0P5B_A12TR u4906 ( .A(rireg[6]), .Y(n3234) );
  MXT2_X0P5M_A12TR u4907 ( .A(rbsr_[6]), .B(wfilebsr[14]), .S0(n4127), .Y(
        n1625) );
  OAI221_X0P5M_A12TR u4908 ( .A0(n3233), .A1(n4152), .B0(n3400), .B1(n4153), 
        .C0(n4158), .Y(n1623) );
  AOI22_X0P5M_A12TR u4909 ( .A0(rbsr_[5]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[5]), .Y(n4158) );
  INV_X0P5B_A12TR u4910 ( .A(wfilebsr[13]), .Y(n3400) );
  INV_X0P5B_A12TR u4911 ( .A(rireg[5]), .Y(n3233) );
  MXT2_X0P5M_A12TR u4912 ( .A(rbsr_[5]), .B(wfilebsr[13]), .S0(n4127), .Y(
        n1622) );
  OAI221_X0P5M_A12TR u4913 ( .A0(n3232), .A1(n4152), .B0(n3397), .B1(n4153), 
        .C0(n4159), .Y(n1620) );
  AOI22_X0P5M_A12TR u4914 ( .A0(rbsr_[4]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[4]), .Y(n4159) );
  INV_X0P5B_A12TR u4915 ( .A(wfilebsr[12]), .Y(n3397) );
  INV_X0P5B_A12TR u4916 ( .A(rireg[4]), .Y(n3232) );
  MXT2_X0P5M_A12TR u4917 ( .A(rbsr_[4]), .B(wfilebsr[12]), .S0(n4127), .Y(
        n1619) );
  OAI221_X0P5M_A12TR u4918 ( .A0(n3231), .A1(n4152), .B0(n3394), .B1(n4153), 
        .C0(n4160), .Y(n1617) );
  AOI22_X0P5M_A12TR u4919 ( .A0(rbsr_[3]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[3]), .Y(n4160) );
  INV_X0P5B_A12TR u4920 ( .A(wfilebsr[11]), .Y(n3394) );
  INV_X0P5B_A12TR u4921 ( .A(rireg[3]), .Y(n3231) );
  MXT2_X0P5M_A12TR u4922 ( .A(rbsr_[3]), .B(wfilebsr[11]), .S0(n4127), .Y(
        n1616) );
  OAI221_X0P5M_A12TR u4923 ( .A0(n3230), .A1(n4152), .B0(n3392), .B1(n4153), 
        .C0(n4161), .Y(n1614) );
  AOI22_X0P5M_A12TR u4924 ( .A0(rbsr_[2]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[2]), .Y(n4161) );
  INV_X0P5B_A12TR u4925 ( .A(wfilebsr[10]), .Y(n3392) );
  INV_X0P5B_A12TR u4926 ( .A(rireg[2]), .Y(n3230) );
  MXT2_X0P5M_A12TR u4927 ( .A(rbsr_[2]), .B(wfilebsr[10]), .S0(n4127), .Y(
        n1613) );
  OAI221_X0P5M_A12TR u4928 ( .A0(n3229), .A1(n4152), .B0(n3390), .B1(n4153), 
        .C0(n4162), .Y(n1611) );
  AOI22_X0P5M_A12TR u4929 ( .A0(rbsr_[1]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[1]), .Y(n4162) );
  INV_X0P5B_A12TR u4930 ( .A(wfilebsr[9]), .Y(n3390) );
  INV_X0P5B_A12TR u4931 ( .A(rireg[1]), .Y(n3229) );
  MXT2_X0P5M_A12TR u4932 ( .A(rbsr_[1]), .B(wfilebsr[9]), .S0(n4127), .Y(n1610) );
  OAI221_X0P5M_A12TR u4933 ( .A0(n3227), .A1(n4152), .B0(n3384), .B1(n4153), 
        .C0(n4163), .Y(n1608) );
  AOI22_X0P5M_A12TR u4934 ( .A0(rbsr_[0]), .A1(n4155), .B0(n4156), .B1(
        dwb_dat_o[0]), .Y(n4163) );
  INV_X0P5B_A12TR u4935 ( .A(n4164), .Y(n4156) );
  AOI211_X0P5M_A12TR u4936 ( .A0(n4165), .A1(n3424), .B0(n3476), .C0(n3239), 
        .Y(n4155) );
  INV_X0P5B_A12TR u4937 ( .A(n3473), .Y(n3424) );
  NOR2_X0P5A_A12TR u4938 ( .A(n3423), .B(n3645), .Y(n3473) );
  OR2_X0P5M_A12TR u4939 ( .A(n3111), .B(n3423), .Y(n4165) );
  NAND3_X0P5A_A12TR u4940 ( .A(n4152), .B(n4164), .C(n4166), .Y(n4153) );
  NAND3_X0P5A_A12TR u4941 ( .A(n4167), .B(n3242), .C(n3472), .Y(n4166) );
  NAND3_X0P5A_A12TR u4942 ( .A(n3111), .B(n3242), .C(n3422), .Y(n4164) );
  NOR2_X0P5A_A12TR u4943 ( .A(n3423), .B(n3597), .Y(n3422) );
  NOR2B_X0P5M_A12TR u4944 ( .AN(n3680), .B(n3682), .Y(n3111) );
  NAND2_X0P5A_A12TR u4945 ( .A(n3317), .B(n3679), .Y(n3682) );
  INV_X0P5B_A12TR u4946 ( .A(wfilebsr[8]), .Y(n3384) );
  NAND4_X0P5A_A12TR u4947 ( .A(n3423), .B(n3551), .C(n3242), .D(n4168), .Y(
        n4152) );
  AND3_X0P5M_A12TR u4948 ( .A(n4169), .B(rmxalu[3]), .C(rmxdst[0]), .Y(n4168)
         );
  INV_X0P5B_A12TR u4949 ( .A(rireg[0]), .Y(n3227) );
  MXT2_X0P5M_A12TR u4950 ( .A(rbsr_[0]), .B(wfilebsr[8]), .S0(n4127), .Y(n1607) );
  OAI211_X0P5M_A12TR u4951 ( .A0(qena[3]), .A1(n3528), .B0(n4170), .C0(n4171), 
        .Y(n1605) );
  AOI211_X0P5M_A12TR u4952 ( .A0(n4172), .A1(n4048), .B0(n4173), .C0(n4174), 
        .Y(n4171) );
  MXT2_X0P5M_A12TR u4953 ( .A(n4175), .B(n4176), .S0(reaptr[1]), .Y(n4170) );
  OAI211_X0P5M_A12TR u4954 ( .A0(qena[3]), .A1(n3479), .B0(n4176), .C0(n4177), 
        .Y(n1603) );
  AOI21_X0P5M_A12TR u4955 ( .A0(n4178), .A1(reaptr[1]), .B0(n4174), .Y(n4177)
         );
  AOI21_X0P5M_A12TR u4956 ( .A0(reaptr[0]), .A1(n4178), .B0(n4179), .Y(n4176)
         );
  OAI221_X0P5M_A12TR u4957 ( .A0(n4055), .A1(n4175), .B0(qena[3]), .B1(n3483), 
        .C0(n4180), .Y(n1601) );
  OA21A1OI2_X0P5M_A12TR u4958 ( .A0(n4173), .A1(n4172), .B0(n4048), .C0(n4179), 
        .Y(n4180) );
  INV_X0P5B_A12TR u4959 ( .A(n4181), .Y(n4179) );
  AND3_X0P5M_A12TR u4960 ( .A(n4056), .B(n4055), .C(n4182), .Y(n4173) );
  OAI211_X0P5M_A12TR u4961 ( .A0(qena[3]), .A1(n3543), .B0(n4183), .C0(n4184), 
        .Y(n1599) );
  AOI21_X0P5M_A12TR u4962 ( .A0(n4172), .A1(reaptr[3]), .B0(n4174), .Y(n4184)
         );
  AND2_X0P5M_A12TR u4963 ( .A(n4185), .B(n4186), .Y(n4174) );
  AND3_X0P5M_A12TR u4964 ( .A(reaptr[5]), .B(n4047), .C(n4185), .Y(n4172) );
  AND3_X0P5M_A12TR u4965 ( .A(n4187), .B(n4188), .C(n4189), .Y(n4185) );
  NOR3_X0P5A_A12TR u4966 ( .A(n4056), .B(reaptr[2]), .C(n4055), .Y(n4189) );
  INV_X0P5B_A12TR u4967 ( .A(reaptr[1]), .Y(n4055) );
  MXIT2_X0P5M_A12TR u4968 ( .A(n4190), .B(n4178), .S0(n4056), .Y(n4183) );
  INV_X0P5B_A12TR u4969 ( .A(reaptr[0]), .Y(n4056) );
  NOR2B_X0P5M_A12TR u4970 ( .AN(n4182), .B(reaptr[3]), .Y(n4178) );
  NAND2_X0P5A_A12TR u4971 ( .A(n4181), .B(n4175), .Y(n4190) );
  NAND2_X0P5A_A12TR u4972 ( .A(n4182), .B(reaptr[3]), .Y(n4175) );
  AND3_X0P5M_A12TR u4973 ( .A(n4187), .B(n4188), .C(n4191), .Y(n4182) );
  NOR3_X0P5A_A12TR u4974 ( .A(n4050), .B(reaptr[4]), .C(n4046), .Y(n4191) );
  INV_X0P5B_A12TR u4975 ( .A(reaptr[5]), .Y(n4046) );
  INV_X0P5B_A12TR u4976 ( .A(reaptr[2]), .Y(n4050) );
  NAND4_X0P5A_A12TR u4977 ( .A(n4186), .B(n4187), .C(n4188), .D(reaptr[2]), 
        .Y(n4181) );
  AND4_X0P5M_A12TR u4978 ( .A(reaptr[8]), .B(qena[3]), .C(reaptr[9]), .D(n4192), .Y(n4188) );
  AND3_X0P5M_A12TR u4979 ( .A(reaptr[6]), .B(reaptr[11]), .C(reaptr[7]), .Y(
        n4192) );
  AND2_X0P5M_A12TR u4980 ( .A(n4193), .B(reaptr[10]), .Y(n4187) );
  MXIT2_X0P5M_A12TR u4981 ( .A(n4194), .B(n4195), .S0(n3399), .Y(n4193) );
  NAND3_X0P5A_A12TR u4982 ( .A(n3403), .B(n3405), .C(n3401), .Y(n4195) );
  INV_X0P5B_A12TR u4983 ( .A(reaptr[14]), .Y(n3403) );
  NAND3_X0P5A_A12TR u4984 ( .A(reaptr[14]), .B(reaptr[13]), .C(reaptr[15]), 
        .Y(n4194) );
  NOR3_X0P5A_A12TR u4985 ( .A(n4047), .B(reaptr[5]), .C(n4048), .Y(n4186) );
  INV_X0P5B_A12TR u4986 ( .A(reaptr[3]), .Y(n4048) );
  INV_X0P5B_A12TR u4987 ( .A(reaptr[4]), .Y(n4047) );
  NAND4_X0P5A_A12TR u4988 ( .A(n4196), .B(n4197), .C(n4198), .D(n4199), .Y(
        n1597) );
  AOI222_X0P5M_A12TR u4989 ( .A0(wfsrplusw1[0]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[0]), .C0(n3815), .C1(wfsrinc2[0]), .Y(n4199) );
  AOI222_X0P5M_A12TR u4990 ( .A0(n3724), .A1(rfsr0l[0]), .B0(wfsrplusw2[0]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[0]), .Y(n4198) );
  AOI222_X0P5M_A12TR u4991 ( .A0(n3723), .A1(rfsr2l[0]), .B0(wfsrplusw0[0]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[0]), .Y(n4197) );
  AOI222_X0P5M_A12TR u4992 ( .A0(dwb_adr_o[0]), .A1(n3819), .B0(n3820), .B1(
        rromlat[0]), .C0(reaptr[0]), .C1(n3821), .Y(n4196) );
  OAI221_X0P5M_A12TR u4993 ( .A0(n3064), .A1(n4200), .B0(n3066), .B1(n3470), 
        .C0(n4201), .Y(n1595) );
  AOI22_X0P5M_A12TR u4994 ( .A0(n2750), .A1(n3069), .B0(n3871), .B1(wpclat[6]), 
        .Y(n4201) );
  INV_X0P5B_A12TR u4995 ( .A(wstkw[7]), .Y(n4200) );
  OAI211_X0P5M_A12TR u4996 ( .A0(qena[1]), .A1(n3777), .B0(n4202), .C0(n4203), 
        .Y(n1594) );
  AOI222_X0P5M_A12TR u4997 ( .A0(wpcinc[6]), .A1(n3792), .B0(n392), .B1(n3793), 
        .C0(n3794), .C1(wstkw[7]), .Y(n4203) );
  AOI22_X0P5M_A12TR u4998 ( .A0(n372), .A1(n3795), .B0(n3796), .B1(rireg[6]), 
        .Y(n4202) );
  INV_X0P5B_A12TR u4999 ( .A(rpcnxt[6]), .Y(n3777) );
  OAI221_X0P5M_A12TR u5000 ( .A0(n3064), .A1(n3669), .B0(n3066), .B1(n3466), 
        .C0(n4204), .Y(n1592) );
  AOI22_X0P5M_A12TR u5001 ( .A0(n2784), .A1(n3069), .B0(n3871), .B1(wpclat[4]), 
        .Y(n4204) );
  INV_X0P5B_A12TR u5002 ( .A(wstkw[5]), .Y(n3669) );
  NAND4_X0P5A_A12TR u5003 ( .A(n4205), .B(n4206), .C(n4207), .D(n4208), .Y(
        n1591) );
  AOI222_X0P5M_A12TR u5004 ( .A0(rpcnxt[4]), .A1(n3375), .B0(wpcinc[4]), .B1(
        n3792), .C0(n3796), .C1(rireg[4]), .Y(n4208) );
  AOI22_X0P5M_A12TR u5005 ( .A0(n390), .A1(n3793), .B0(n3794), .B1(wstkw[5]), 
        .Y(n4207) );
  NAND4_X0P5A_A12TR u5006 ( .A(n370), .B(n4209), .C(n3738), .D(rbcc), .Y(n4205) );
  OAI221_X0P5M_A12TR u5007 ( .A0(n3064), .A1(n4210), .B0(n3066), .B1(n3453), 
        .C0(n4211), .Y(n1589) );
  AOI22_X0P5M_A12TR u5008 ( .A0(n2751), .A1(n3069), .B0(n3871), .B1(wpclat[0]), 
        .Y(n4211) );
  INV_X0P5B_A12TR u5009 ( .A(wstkw[1]), .Y(n4210) );
  OAI222_X0P5M_A12TR u5010 ( .A0(n3470), .A1(n4212), .B0(n3780), .B1(n4213), 
        .C0(n4214), .C1(n4215), .Y(n1588) );
  MXIT2_X0P5M_A12TR u5011 ( .A(n4215), .B(n3780), .S0(n4127), .Y(n1587) );
  INV_X0P5B_A12TR u5012 ( .A(rwreg_[7]), .Y(n4215) );
  OAI221_X0P5M_A12TR u5013 ( .A0(n3780), .A1(n4216), .B0(n4430), .B1(n3738), 
        .C0(n4217), .Y(n1586) );
  AOI222_X0P5M_A12TR u5014 ( .A0(n4218), .A1(n3972), .B0(n4219), .B1(n3782), 
        .C0(n4220), .C1(rireg[7]), .Y(n4217) );
  MXT2_X0P5M_A12TR u5015 ( .A(dwb_dat_i[7]), .B(rsfrdat[7]), .S0(rsfrstb), .Y(
        n3782) );
  INV_X0P5B_A12TR u5016 ( .A(rmask[7]), .Y(n3972) );
  INV_X0P5B_A12TR u5017 ( .A(rtgt[7]), .Y(n4430) );
  INV_X0P5B_A12TR u5018 ( .A(rwreg[7]), .Y(n3780) );
  OAI222_X0P5M_A12TR u5019 ( .A0(n3468), .A1(n4212), .B0(n3911), .B1(n4213), 
        .C0(n4214), .C1(n4221), .Y(n1584) );
  MXIT2_X0P5M_A12TR u5020 ( .A(n4221), .B(n3911), .S0(n4127), .Y(n1583) );
  INV_X0P5B_A12TR u5021 ( .A(rwreg_[6]), .Y(n4221) );
  OAI221_X0P5M_A12TR u5022 ( .A0(n3911), .A1(n4216), .B0(n4429), .B1(n3738), 
        .C0(n4222), .Y(n1582) );
  AOI222_X0P5M_A12TR u5023 ( .A0(n4218), .A1(n3945), .B0(n4219), .B1(n3914), 
        .C0(n4220), .C1(rireg[6]), .Y(n4222) );
  MXT2_X0P5M_A12TR u5024 ( .A(dwb_dat_i[6]), .B(rsfrdat[6]), .S0(rsfrstb), .Y(
        n3914) );
  INV_X0P5B_A12TR u5025 ( .A(rmask[6]), .Y(n3945) );
  INV_X0P5B_A12TR u5026 ( .A(rtgt[6]), .Y(n4429) );
  INV_X0P5B_A12TR u5027 ( .A(rwreg[6]), .Y(n3911) );
  OAI222_X0P5M_A12TR u5028 ( .A0(n3466), .A1(n4212), .B0(n4129), .B1(n4213), 
        .C0(n4214), .C1(n4223), .Y(n1580) );
  MXIT2_X0P5M_A12TR u5029 ( .A(n4223), .B(n4129), .S0(n4127), .Y(n1579) );
  INV_X0P5B_A12TR u5030 ( .A(rwreg_[5]), .Y(n4223) );
  OAI221_X0P5M_A12TR u5031 ( .A0(n4129), .A1(n4216), .B0(n4428), .B1(n3738), 
        .C0(n4224), .Y(n1578) );
  AOI222_X0P5M_A12TR u5032 ( .A0(n4218), .A1(n4225), .B0(n4219), .B1(n4132), 
        .C0(n4220), .C1(rireg[5]), .Y(n4224) );
  MXT2_X0P5M_A12TR u5033 ( .A(dwb_dat_i[5]), .B(rsfrdat[5]), .S0(rsfrstb), .Y(
        n4132) );
  INV_X0P5B_A12TR u5034 ( .A(rmask[5]), .Y(n4225) );
  INV_X0P5B_A12TR u5035 ( .A(rtgt[5]), .Y(n4428) );
  INV_X0P5B_A12TR u5036 ( .A(rwreg[5]), .Y(n4129) );
  OAI222_X0P5M_A12TR u5037 ( .A0(n3148), .A1(n4212), .B0(n3822), .B1(n4213), 
        .C0(n4214), .C1(n4226), .Y(n1576) );
  MXIT2_X0P5M_A12TR u5038 ( .A(n4226), .B(n3822), .S0(n4127), .Y(n1575) );
  INV_X0P5B_A12TR u5039 ( .A(rwreg_[4]), .Y(n4226) );
  OAI221_X0P5M_A12TR u5040 ( .A0(n3822), .A1(n4216), .B0(n4427), .B1(n3738), 
        .C0(n4227), .Y(n1574) );
  AOI222_X0P5M_A12TR u5041 ( .A0(n4218), .A1(n4228), .B0(n4219), .B1(n3825), 
        .C0(n4220), .C1(rireg[4]), .Y(n4227) );
  MXT2_X0P5M_A12TR u5042 ( .A(dwb_dat_i[4]), .B(rsfrdat[4]), .S0(rsfrstb), .Y(
        n3825) );
  INV_X0P5B_A12TR u5043 ( .A(rmask[4]), .Y(n4228) );
  INV_X0P5B_A12TR u5044 ( .A(rtgt[4]), .Y(n4427) );
  INV_X0P5B_A12TR u5045 ( .A(rwreg[4]), .Y(n3822) );
  OAI222_X0P5M_A12TR u5046 ( .A0(n3458), .A1(n4212), .B0(n3882), .B1(n4213), 
        .C0(n4214), .C1(n4229), .Y(n1572) );
  MXIT2_X0P5M_A12TR u5047 ( .A(n4229), .B(n3882), .S0(n4127), .Y(n1571) );
  INV_X0P5B_A12TR u5048 ( .A(rwreg_[3]), .Y(n4229) );
  OAI221_X0P5M_A12TR u5049 ( .A0(n3882), .A1(n4216), .B0(n4426), .B1(n3738), 
        .C0(n4230), .Y(n1570) );
  AOI222_X0P5M_A12TR u5050 ( .A0(n4218), .A1(n3958), .B0(n4219), .B1(n3885), 
        .C0(n4220), .C1(rireg[3]), .Y(n4230) );
  MXT2_X0P5M_A12TR u5051 ( .A(dwb_dat_i[3]), .B(rsfrdat[3]), .S0(rsfrstb), .Y(
        n3885) );
  INV_X0P5B_A12TR u5052 ( .A(rmask[3]), .Y(n3958) );
  INV_X0P5B_A12TR u5053 ( .A(rtgt[3]), .Y(n4426) );
  INV_X0P5B_A12TR u5054 ( .A(rwreg[3]), .Y(n3882) );
  OAI222_X0P5M_A12TR u5055 ( .A0(n3158), .A1(n4212), .B0(n3856), .B1(n4213), 
        .C0(n4214), .C1(n4231), .Y(n1568) );
  MXIT2_X0P5M_A12TR u5056 ( .A(n4231), .B(n3856), .S0(n4127), .Y(n1567) );
  INV_X0P5B_A12TR u5057 ( .A(rwreg_[2]), .Y(n4231) );
  OAI221_X0P5M_A12TR u5058 ( .A0(n3856), .A1(n4216), .B0(n4425), .B1(n3738), 
        .C0(n4232), .Y(n1566) );
  AOI222_X0P5M_A12TR u5059 ( .A0(n4218), .A1(n3942), .B0(n4219), .B1(n3859), 
        .C0(n4220), .C1(rireg[2]), .Y(n4232) );
  MXT2_X0P5M_A12TR u5060 ( .A(dwb_dat_i[2]), .B(rsfrdat[2]), .S0(rsfrstb), .Y(
        n3859) );
  INV_X0P5B_A12TR u5061 ( .A(rmask[2]), .Y(n3942) );
  INV_X0P5B_A12TR u5062 ( .A(rtgt[2]), .Y(n4425) );
  INV_X0P5B_A12TR u5063 ( .A(rwreg[2]), .Y(n3856) );
  OAI222_X0P5M_A12TR u5064 ( .A0(n3453), .A1(n4212), .B0(n3798), .B1(n4213), 
        .C0(n4214), .C1(n4233), .Y(n1564) );
  MXIT2_X0P5M_A12TR u5065 ( .A(n4233), .B(n3798), .S0(n4127), .Y(n1563) );
  INV_X0P5B_A12TR u5066 ( .A(rwreg_[1]), .Y(n4233) );
  OAI221_X0P5M_A12TR u5067 ( .A0(n3798), .A1(n4216), .B0(n4424), .B1(n3738), 
        .C0(n4234), .Y(n1562) );
  AOI222_X0P5M_A12TR u5068 ( .A0(n4218), .A1(n3960), .B0(n4219), .B1(n3801), 
        .C0(n4220), .C1(rireg[1]), .Y(n4234) );
  MXT2_X0P5M_A12TR u5069 ( .A(dwb_dat_i[1]), .B(rsfrdat[1]), .S0(rsfrstb), .Y(
        n3801) );
  INV_X0P5B_A12TR u5070 ( .A(rmask[1]), .Y(n3960) );
  INV_X0P5B_A12TR u5071 ( .A(rtgt[1]), .Y(n4424) );
  INV_X0P5B_A12TR u5072 ( .A(rwreg[1]), .Y(n3798) );
  OAI222_X0P5M_A12TR u5073 ( .A0(n3067), .A1(n4212), .B0(n3736), .B1(n4213), 
        .C0(n4214), .C1(n4235), .Y(n1560) );
  NAND3B_X0P5M_A12TR u5074 ( .AN(n4236), .B(n3688), .C(n4167), .Y(n4214) );
  OAI21_X0P5M_A12TR u5075 ( .A0(n3239), .A1(n4237), .B0(n4212), .Y(n4213) );
  INV_X0P5B_A12TR u5076 ( .A(n4167), .Y(n3239) );
  NOR2_X0P5A_A12TR u5077 ( .A(n4238), .B(rmxsha[1]), .Y(n4167) );
  NAND2_X0P5A_A12TR u5078 ( .A(n3688), .B(n4236), .Y(n4212) );
  OAI22_X0P5M_A12TR u5079 ( .A0(rmxdst[0]), .A1(n3551), .B0(n3597), .B1(n3671), 
        .Y(n4236) );
  NAND3_X0P5A_A12TR u5080 ( .A(n3317), .B(dwb_adr_o[3]), .C(n3680), .Y(n3671)
         );
  NOR3_X0P5A_A12TR u5081 ( .A(dwb_adr_o[2]), .B(dwb_adr_o[4]), .C(n3684), .Y(
        n3680) );
  INV_X0P5B_A12TR u5082 ( .A(rmxdst[1]), .Y(n3551) );
  MXIT2_X0P5M_A12TR u5083 ( .A(n4235), .B(n3736), .S0(n4127), .Y(n1559) );
  INV_X0P5B_A12TR u5084 ( .A(rwreg_[0]), .Y(n4235) );
  NAND4_X0P5A_A12TR u5085 ( .A(n4239), .B(n4240), .C(n4241), .D(n4242), .Y(
        n1558) );
  AOI222_X0P5M_A12TR u5086 ( .A0(wfsrplusw1[2]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[2]), .C0(n3815), .C1(wfsrinc2[2]), .Y(n4242) );
  AOI222_X0P5M_A12TR u5087 ( .A0(n3724), .A1(rfsr0l[2]), .B0(wfsrplusw2[2]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[2]), .Y(n4241) );
  AOI222_X0P5M_A12TR u5088 ( .A0(n3723), .A1(rfsr2l[2]), .B0(wfsrplusw0[2]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[2]), .Y(n4240) );
  AOI222_X0P5M_A12TR u5089 ( .A0(dwb_adr_o[2]), .A1(n3819), .B0(n3820), .B1(
        rromlat[2]), .C0(reaptr[2]), .C1(n3821), .Y(n4239) );
  MXIT2_X0P5M_A12TR u5090 ( .A(n3157), .B(n3153), .S0(n4127), .Y(n1556) );
  INV_X0P5B_A12TR u5091 ( .A(rz), .Y(n3153) );
  INV_X0P5B_A12TR u5092 ( .A(rstatus_[2]), .Y(n3157) );
  OAI222_X0P5M_A12TR u5093 ( .A0(n3148), .A1(n3776), .B0(n3628), .B1(n3778), 
        .C0(qena[3]), .C1(n4243), .Y(n1555) );
  INV_X0P5B_A12TR u5094 ( .A(wpclat[3]), .Y(n4243) );
  OAI221_X0P5M_A12TR u5095 ( .A0(n3064), .A1(n4244), .B0(n3066), .B1(n3148), 
        .C0(n4245), .Y(n1553) );
  AOI22_X0P5M_A12TR u5096 ( .A0(n2783), .A1(n3069), .B0(n3871), .B1(wpclat[3]), 
        .Y(n4245) );
  OAI211_X0P5M_A12TR u5097 ( .A0(qena[1]), .A1(n3628), .B0(n4246), .C0(n4247), 
        .Y(n1552) );
  AOI211_X0P5M_A12TR u5098 ( .A0(n389), .A1(n3793), .B0(n4248), .C0(n4249), 
        .Y(n4247) );
  NOR3_X0P5A_A12TR u5099 ( .A(n3937), .B(n4250), .C(n4053), .Y(n4249) );
  AOI32_X0P5M_A12TR u5100 ( .A0(n3738), .A1(rbcc), .A2(n369), .B0(qena[1]), 
        .B1(n4001), .Y(n4250) );
  OAI31_X0P5M_A12TR u5101 ( .A0(n4251), .A1(rmxnpc[1]), .A2(n4244), .B0(n4206), 
        .Y(n4248) );
  NAND3_X0P5A_A12TR u5102 ( .A(qena[1]), .B(n4053), .C(n4209), .Y(n4206) );
  INV_X0P5B_A12TR u5103 ( .A(wstkw[4]), .Y(n4244) );
  AOI22_X0P5M_A12TR u5104 ( .A0(wpcinc[3]), .A1(n3792), .B0(n3796), .B1(
        rireg[3]), .Y(n4246) );
  INV_X0P5B_A12TR u5105 ( .A(rpcnxt[3]), .Y(n3628) );
  AO22_X0P5M_A12TR u5106 ( .A0(n3074), .A1(rpcl_0_), .B0(dwb_dat_o[0]), .B1(
        n3709), .Y(n1550) );
  OAI222_X0P5M_A12TR u5107 ( .A0(n3468), .A1(n4252), .B0(n3905), .B1(n4253), 
        .C0(n3906), .C1(n4254), .Y(n1548) );
  INV_X0P5B_A12TR u5108 ( .A(wpclat[13]), .Y(n3906) );
  INV_X0P5B_A12TR u5109 ( .A(rpclath[6]), .Y(n3905) );
  OAI222_X0P5M_A12TR u5110 ( .A0(n3466), .A1(n4252), .B0(n4255), .B1(n4253), 
        .C0(n4254), .C1(n4256), .Y(n1547) );
  OAI222_X0P5M_A12TR u5111 ( .A0(n4255), .A1(n3776), .B0(n4257), .B1(n3778), 
        .C0(qena[3]), .C1(n4256), .Y(n1546) );
  INV_X0P5B_A12TR u5112 ( .A(wpclat[12]), .Y(n4256) );
  INV_X0P5B_A12TR u5113 ( .A(rpclath[5]), .Y(n4255) );
  OAI221_X0P5M_A12TR u5114 ( .A0(n3907), .A1(n4258), .B0(n3466), .B1(n3909), 
        .C0(n4259), .Y(n1544) );
  AOI22_X0P5M_A12TR u5115 ( .A0(n2752), .A1(n3069), .B0(wpclat[12]), .B1(n3871), .Y(n4259) );
  INV_X0P5B_A12TR u5116 ( .A(wstkw[13]), .Y(n4258) );
  OAI211_X0P5M_A12TR u5117 ( .A0(qena[1]), .A1(n4257), .B0(n4260), .C0(n4261), 
        .Y(n1543) );
  AOI222_X0P5M_A12TR u5118 ( .A0(wpcinc[12]), .A1(n3792), .B0(n398), .B1(n3793), .C0(n3794), .C1(wstkw[13]), .Y(n4261) );
  AOI22_X0P5M_A12TR u5119 ( .A0(n378), .A1(n3795), .B0(n3796), .B1(rromlat[4]), 
        .Y(n4260) );
  INV_X0P5B_A12TR u5120 ( .A(rpcnxt[12]), .Y(n4257) );
  OAI222_X0P5M_A12TR u5121 ( .A0(n3148), .A1(n4252), .B0(n4262), .B1(n4253), 
        .C0(n4254), .C1(n4263), .Y(n1541) );
  OAI222_X0P5M_A12TR u5122 ( .A0(n4262), .A1(n3776), .B0(n4264), .B1(n3778), 
        .C0(qena[3]), .C1(n4263), .Y(n1540) );
  INV_X0P5B_A12TR u5123 ( .A(wpclat[11]), .Y(n4263) );
  INV_X0P5B_A12TR u5124 ( .A(rpclath[4]), .Y(n4262) );
  OAI221_X0P5M_A12TR u5125 ( .A0(n3907), .A1(n4265), .B0(n3148), .B1(n3909), 
        .C0(n4266), .Y(n1538) );
  AOI22_X0P5M_A12TR u5126 ( .A0(n2753), .A1(n3069), .B0(wpclat[11]), .B1(n3871), .Y(n4266) );
  INV_X0P5B_A12TR u5127 ( .A(wstkw[12]), .Y(n4265) );
  OAI211_X0P5M_A12TR u5128 ( .A0(qena[1]), .A1(n4264), .B0(n4267), .C0(n4268), 
        .Y(n1537) );
  AOI222_X0P5M_A12TR u5129 ( .A0(wpcinc[11]), .A1(n3792), .B0(n397), .B1(n3793), .C0(n3794), .C1(wstkw[12]), .Y(n4268) );
  AOI22_X0P5M_A12TR u5130 ( .A0(n377), .A1(n3795), .B0(n3796), .B1(rromlat[3]), 
        .Y(n4267) );
  INV_X0P5B_A12TR u5131 ( .A(rpcnxt[11]), .Y(n4264) );
  OAI222_X0P5M_A12TR u5132 ( .A0(n3458), .A1(n4252), .B0(n4269), .B1(n4253), 
        .C0(n4254), .C1(n4270), .Y(n1535) );
  OAI222_X0P5M_A12TR u5133 ( .A0(n4269), .A1(n3776), .B0(n4271), .B1(n3778), 
        .C0(qena[3]), .C1(n4270), .Y(n1534) );
  INV_X0P5B_A12TR u5134 ( .A(wpclat[10]), .Y(n4270) );
  INV_X0P5B_A12TR u5135 ( .A(rpclath[3]), .Y(n4269) );
  OAI221_X0P5M_A12TR u5136 ( .A0(n3907), .A1(n4272), .B0(n3458), .B1(n3909), 
        .C0(n4273), .Y(n1532) );
  AOI22_X0P5M_A12TR u5137 ( .A0(n2754), .A1(n3069), .B0(wpclat[10]), .B1(n3871), .Y(n4273) );
  INV_X0P5B_A12TR u5138 ( .A(wstkw[11]), .Y(n4272) );
  OAI211_X0P5M_A12TR u5139 ( .A0(qena[1]), .A1(n4271), .B0(n4274), .C0(n4275), 
        .Y(n1531) );
  AOI222_X0P5M_A12TR u5140 ( .A0(wpcinc[10]), .A1(n3792), .B0(n396), .B1(n3793), .C0(n3794), .C1(wstkw[11]), .Y(n4275) );
  AOI22_X0P5M_A12TR u5141 ( .A0(n376), .A1(n3795), .B0(n3796), .B1(rromlat[2]), 
        .Y(n4274) );
  INV_X0P5B_A12TR u5142 ( .A(rpcnxt[10]), .Y(n4271) );
  OAI222_X0P5M_A12TR u5143 ( .A0(n3158), .A1(n4252), .B0(n4276), .B1(n4253), 
        .C0(n4254), .C1(n4277), .Y(n1529) );
  OAI222_X0P5M_A12TR u5144 ( .A0(n4276), .A1(n3776), .B0(n4278), .B1(n3778), 
        .C0(qena[3]), .C1(n4277), .Y(n1528) );
  INV_X0P5B_A12TR u5145 ( .A(wpclat[9]), .Y(n4277) );
  INV_X0P5B_A12TR u5146 ( .A(rpclath[2]), .Y(n4276) );
  OAI221_X0P5M_A12TR u5147 ( .A0(n3907), .A1(n4279), .B0(n3158), .B1(n3909), 
        .C0(n4280), .Y(n1526) );
  AOI22_X0P5M_A12TR u5148 ( .A0(n2755), .A1(n3069), .B0(wpclat[9]), .B1(n3871), 
        .Y(n4280) );
  INV_X0P5B_A12TR u5149 ( .A(wstkw[10]), .Y(n4279) );
  OAI211_X0P5M_A12TR u5150 ( .A0(qena[1]), .A1(n4278), .B0(n4281), .C0(n4282), 
        .Y(n1525) );
  AOI222_X0P5M_A12TR u5151 ( .A0(wpcinc[9]), .A1(n3792), .B0(n395), .B1(n3793), 
        .C0(n3794), .C1(wstkw[10]), .Y(n4282) );
  AOI22_X0P5M_A12TR u5152 ( .A0(n375), .A1(n3795), .B0(n3796), .B1(rromlat[1]), 
        .Y(n4281) );
  INV_X0P5B_A12TR u5153 ( .A(rpcnxt[9]), .Y(n4278) );
  OAI222_X0P5M_A12TR u5154 ( .A0(n3453), .A1(n4252), .B0(n4283), .B1(n4253), 
        .C0(n4254), .C1(n4284), .Y(n1523) );
  OAI222_X0P5M_A12TR u5155 ( .A0(n4283), .A1(n3776), .B0(n4285), .B1(n3778), 
        .C0(qena[3]), .C1(n4284), .Y(n1522) );
  INV_X0P5B_A12TR u5156 ( .A(wpclat[8]), .Y(n4284) );
  INV_X0P5B_A12TR u5157 ( .A(rpclath[1]), .Y(n4283) );
  OAI221_X0P5M_A12TR u5158 ( .A0(n3907), .A1(n4286), .B0(n3453), .B1(n3909), 
        .C0(n4287), .Y(n1520) );
  AOI22_X0P5M_A12TR u5159 ( .A0(n2756), .A1(n3069), .B0(wpclat[8]), .B1(n3871), 
        .Y(n4287) );
  INV_X0P5B_A12TR u5160 ( .A(wstkw[9]), .Y(n4286) );
  OAI211_X0P5M_A12TR u5161 ( .A0(qena[1]), .A1(n4285), .B0(n4288), .C0(n4289), 
        .Y(n1519) );
  AOI222_X0P5M_A12TR u5162 ( .A0(wpcinc[8]), .A1(n3792), .B0(n394), .B1(n3793), 
        .C0(n3794), .C1(wstkw[9]), .Y(n4289) );
  AOI22_X0P5M_A12TR u5163 ( .A0(n374), .A1(n3795), .B0(n3796), .B1(rromlat[0]), 
        .Y(n4288) );
  INV_X0P5B_A12TR u5164 ( .A(rpcnxt[8]), .Y(n4285) );
  OAI222_X0P5M_A12TR u5165 ( .A0(n3067), .A1(n4252), .B0(n4290), .B1(n4253), 
        .C0(n4254), .C1(n4291), .Y(n1517) );
  OAI222_X0P5M_A12TR u5166 ( .A0(n4290), .A1(n3776), .B0(n4292), .B1(n3778), 
        .C0(qena[3]), .C1(n4291), .Y(n1516) );
  INV_X0P5B_A12TR u5167 ( .A(wpclat[7]), .Y(n4291) );
  INV_X0P5B_A12TR u5168 ( .A(rpclath[0]), .Y(n4290) );
  OAI221_X0P5M_A12TR u5169 ( .A0(n3907), .A1(n4293), .B0(n3067), .B1(n3909), 
        .C0(n4294), .Y(n1514) );
  AOI22_X0P5M_A12TR u5170 ( .A0(n2757), .A1(n3069), .B0(wpclat[7]), .B1(n3871), 
        .Y(n4294) );
  INV_X0P5B_A12TR u5171 ( .A(wstkw[8]), .Y(n4293) );
  OAI211_X0P5M_A12TR u5172 ( .A0(qena[1]), .A1(n4292), .B0(n4295), .C0(n4296), 
        .Y(n1513) );
  AOI222_X0P5M_A12TR u5173 ( .A0(wpcinc[7]), .A1(n3792), .B0(n393), .B1(n3793), 
        .C0(n3794), .C1(wstkw[8]), .Y(n4296) );
  AOI22_X0P5M_A12TR u5174 ( .A0(n373), .A1(n3795), .B0(n3796), .B1(rireg[7]), 
        .Y(n4295) );
  INV_X0P5B_A12TR u5175 ( .A(rpcnxt[7]), .Y(n4292) );
  OAI22_X0P5M_A12TR u5176 ( .A0(n3470), .A1(n4297), .B0(n4298), .B1(n4299), 
        .Y(n1511) );
  INV_X0P5B_A12TR u5177 ( .A(rpclatu[7]), .Y(n4298) );
  OAI22_X0P5M_A12TR u5178 ( .A0(n3468), .A1(n4297), .B0(n4300), .B1(n4299), 
        .Y(n1510) );
  INV_X0P5B_A12TR u5179 ( .A(rpclatu[6]), .Y(n4300) );
  OAI22_X0P5M_A12TR u5180 ( .A0(n3466), .A1(n4297), .B0(n4301), .B1(n4299), 
        .Y(n1509) );
  INV_X0P5B_A12TR u5181 ( .A(rpclatu[5]), .Y(n4301) );
  OAI222_X0P5M_A12TR u5182 ( .A0(n3458), .A1(n4297), .B0(n3877), .B1(n4299), 
        .C0(n3878), .C1(n4254), .Y(n1508) );
  INV_X0P5B_A12TR u5183 ( .A(wpclat[18]), .Y(n3878) );
  INV_X0P5B_A12TR u5184 ( .A(rpclatu[3]), .Y(n3877) );
  OAI22_X0P5M_A12TR u5185 ( .A0(n4302), .A1(n3105), .B0(n3470), .B1(n4303), 
        .Y(n1507) );
  INV_X0P5B_A12TR u5186 ( .A(rtblptru[7]), .Y(n3105) );
  OAI22_X0P5M_A12TR u5187 ( .A0(n4302), .A1(n3326), .B0(n3468), .B1(n4303), 
        .Y(n1506) );
  INV_X0P5B_A12TR u5188 ( .A(rtblptru[6]), .Y(n3326) );
  OAI22_X0P5M_A12TR u5189 ( .A0(n4302), .A1(n4304), .B0(n3466), .B1(n4303), 
        .Y(n1505) );
  INV_X0P5B_A12TR u5190 ( .A(rtblptru[5]), .Y(n4304) );
  OAI22_X0P5M_A12TR u5191 ( .A0(n4302), .A1(n3170), .B0(n3148), .B1(n4303), 
        .Y(n1504) );
  NAND3_X0P5A_A12TR u5192 ( .A(n3240), .B(n3242), .C(n3268), .Y(n4303) );
  INV_X0P5B_A12TR u5193 ( .A(n3104), .Y(n3268) );
  INV_X0P5B_A12TR u5194 ( .A(rtblptru[4]), .Y(n3170) );
  AOI211_X0P5M_A12TR u5195 ( .A0(n3104), .A1(qfsm[0]), .B0(n3248), .C0(n3476), 
        .Y(n4302) );
  NOR2_X0P5A_A12TR u5196 ( .A(n4305), .B(n3645), .Y(n3248) );
  NAND2_X0P5A_A12TR u5197 ( .A(n4306), .B(n3317), .Y(n3104) );
  OAI221_X0P5M_A12TR u5198 ( .A0(n3405), .A1(n3719), .B0(n3720), .B1(n4307), 
        .C0(n4308), .Y(n1503) );
  AOI222_X0P5M_A12TR u5199 ( .A0(n3723), .A1(n3125), .B0(n3724), .B1(rfsr0h[7]), .C0(n3725), .C1(rfsr1h[7]), .Y(n4308) );
  INV_X0P5B_A12TR u5200 ( .A(n1940), .Y(n3125) );
  INV_X0P5B_A12TR u5201 ( .A(rdwbadr[15]), .Y(n4307) );
  INV_X0P5B_A12TR u5202 ( .A(reaptr[15]), .Y(n3405) );
  OAI221_X0P5M_A12TR u5203 ( .A0(n3401), .A1(n3719), .B0(n3720), .B1(n4309), 
        .C0(n4310), .Y(n1501) );
  AOI222_X0P5M_A12TR u5204 ( .A0(n3723), .A1(n3681), .B0(n3724), .B1(rfsr0h[5]), .C0(n3725), .C1(rfsr1h[5]), .Y(n4310) );
  INV_X0P5B_A12TR u5205 ( .A(n1942), .Y(n3681) );
  INV_X0P5B_A12TR u5206 ( .A(rdwbadr[13]), .Y(n4309) );
  INV_X0P5B_A12TR u5207 ( .A(reaptr[13]), .Y(n3401) );
  OAI221_X0P5M_A12TR u5208 ( .A0(n3399), .A1(n3719), .B0(n3720), .B1(n4311), 
        .C0(n4312), .Y(n1499) );
  AOI222_X0P5M_A12TR u5209 ( .A0(n3723), .A1(rfsr2h[4]), .B0(n3724), .B1(
        rfsr0h[4]), .C0(n3725), .C1(rfsr1h[4]), .Y(n4312) );
  INV_X0P5B_A12TR u5210 ( .A(rdwbadr[12]), .Y(n4311) );
  INV_X0P5B_A12TR u5211 ( .A(n3819), .Y(n3720) );
  INV_X0P5B_A12TR u5212 ( .A(reaptr[12]), .Y(n3399) );
  OAI221_X0P5M_A12TR u5213 ( .A0(n3736), .A1(n4216), .B0(n4423), .B1(n3738), 
        .C0(n4313), .Y(n1497) );
  AOI222_X0P5M_A12TR u5214 ( .A0(n4218), .A1(n4314), .B0(n4219), .B1(n3743), 
        .C0(n4220), .C1(rireg[0]), .Y(n4313) );
  AND3_X0P5M_A12TR u5215 ( .A(rmxtgt[0]), .B(n3738), .C(rmxtgt[1]), .Y(n4220)
         );
  MXT2_X0P5M_A12TR u5216 ( .A(dwb_dat_i[0]), .B(rsfrdat[0]), .S0(rsfrstb), .Y(
        n3743) );
  AND3_X0P5M_A12TR u5217 ( .A(n3738), .B(n3931), .C(rmxtgt[0]), .Y(n4219) );
  INV_X0P5B_A12TR u5218 ( .A(rmask[0]), .Y(n4314) );
  AND3_X0P5M_A12TR u5219 ( .A(n3738), .B(n4315), .C(rmxtgt[1]), .Y(n4218) );
  INV_X0P5B_A12TR u5220 ( .A(wneg[0]), .Y(n4423) );
  NAND3_X0P5A_A12TR u5221 ( .A(n4315), .B(n3931), .C(n3738), .Y(n4216) );
  INV_X0P5B_A12TR u5222 ( .A(rmxtgt[1]), .Y(n3931) );
  INV_X0P5B_A12TR u5223 ( .A(rmxtgt[0]), .Y(n4315) );
  INV_X0P5B_A12TR u5224 ( .A(rwreg[0]), .Y(n3736) );
  NAND2_X0P5A_A12TR u5225 ( .A(n4316), .B(n4317), .Y(n1495) );
  AOI211_X0P5M_A12TR u5226 ( .A0(wadd[8]), .A1(n3763), .B0(n4318), .C0(n4319), 
        .Y(n4317) );
  NOR2_X0P5A_A12TR u5227 ( .A(n2779), .B(n3755), .Y(n4319) );
  INV_X0P5B_A12TR u5228 ( .A(n3775), .Y(n3755) );
  NOR3_X0P5A_A12TR u5229 ( .A(n3765), .B(n4069), .C(n4143), .Y(n3775) );
  INV_X0P5B_A12TR u5230 ( .A(n4169), .Y(n4143) );
  OAI22_X0P5M_A12TR u5231 ( .A0(wsub[8]), .A1(n4146), .B0(n4320), .B1(n3550), 
        .Y(n4318) );
  AOI22_X0P5M_A12TR u5232 ( .A0(n3750), .A1(rtgt[7]), .B0(n3759), .B1(wneg[0]), 
        .Y(n4320) );
  AND2_X0P5M_A12TR u5233 ( .A(n4321), .B(rmxalu[1]), .Y(n3759) );
  AND2_X0P5M_A12TR u5234 ( .A(n4321), .B(n4142), .Y(n3750) );
  NOR3_X0P5A_A12TR u5235 ( .A(n4069), .B(rmxalu[2]), .C(n3765), .Y(n4321) );
  INV_X0P5B_A12TR u5236 ( .A(rmxalu[3]), .Y(n4069) );
  NAND3_X0P5A_A12TR u5237 ( .A(rmxalu[2]), .B(n3550), .C(n4140), .Y(n4146) );
  AND2_X0P5M_A12TR u5238 ( .A(n4141), .B(rmxalu[1]), .Y(n4140) );
  INV_X0P5B_A12TR u5239 ( .A(rmxalu[0]), .Y(n3550) );
  AND2_X0P5M_A12TR u5240 ( .A(n4141), .B(n4169), .Y(n3763) );
  NOR3_X0P5A_A12TR u5241 ( .A(rmxalu[0]), .B(rmxalu[1]), .C(n4086), .Y(n4169)
         );
  INV_X0P5B_A12TR u5242 ( .A(rmxalu[2]), .Y(n4086) );
  AOI211_X0P5M_A12TR u5243 ( .A0(waddc[8]), .A1(n3764), .B0(n4322), .C0(n4323), 
        .Y(n4316) );
  NOR2_X0P5A_A12TR u5244 ( .A(wsubc[8]), .B(n4147), .Y(n4323) );
  NAND2_X0P5A_A12TR u5245 ( .A(n4324), .B(rmxalu[1]), .Y(n4147) );
  MXIT2_X0P5M_A12TR u5246 ( .A(n4325), .B(n3715), .S0(n3765), .Y(n4322) );
  INV_X0P5B_A12TR u5247 ( .A(rc_), .Y(n3715) );
  NAND2_X0P5A_A12TR u5248 ( .A(wrrc_7_), .B(n4326), .Y(n4325) );
  AO21A1AI2_X0P5M_A12TR u5249 ( .A0(rmxalu[0]), .A1(rmxalu[3]), .B0(rmxalu[2]), 
        .C0(n4327), .Y(n4326) );
  OAI211_X0P5M_A12TR u5250 ( .A0(rmxalu[1]), .A1(rmxalu[0]), .B0(rmxalu[2]), 
        .C0(rmxalu[3]), .Y(n4327) );
  AND2_X0P5M_A12TR u5251 ( .A(n4324), .B(n4142), .Y(n3764) );
  INV_X0P5B_A12TR u5252 ( .A(rmxalu[1]), .Y(n4142) );
  AND3_X0P5M_A12TR u5253 ( .A(rmxalu[0]), .B(rmxalu[2]), .C(n4141), .Y(n4324)
         );
  NOR2_X0P5A_A12TR u5254 ( .A(n3765), .B(rmxalu[3]), .Y(n4141) );
  INV_X0P5B_A12TR u5255 ( .A(n3940), .Y(n3765) );
  NOR2_X0P5A_A12TR u5256 ( .A(n3932), .B(n3708), .Y(n3940) );
  INV_X0P5B_A12TR u5257 ( .A(qena[2]), .Y(n3932) );
  NAND2_X0P5A_A12TR u5258 ( .A(n4328), .B(n3228), .Y(n1481) );
  MXIT2_X0P5M_A12TR u5259 ( .A(iwb_sel_o[1]), .B(n4329), .S0(n3054), .Y(n4328)
         );
  NOR2_X0P5A_A12TR u5260 ( .A(n4305), .B(n3558), .Y(n4329) );
  INV_X0P5B_A12TR u5261 ( .A(wtblat[0]), .Y(n3558) );
  NAND2_X0P5A_A12TR u5262 ( .A(n4330), .B(n3228), .Y(n1471) );
  INV_X0P5B_A12TR u5263 ( .A(n3625), .Y(n3228) );
  NOR2_X0P5A_A12TR u5264 ( .A(n3423), .B(n3221), .Y(n3625) );
  INV_X0P5B_A12TR u5265 ( .A(n3472), .Y(n3423) );
  NOR2_X0P5A_A12TR u5266 ( .A(n4305), .B(n4119), .Y(n3472) );
  MXIT2_X0P5M_A12TR u5267 ( .A(iwb_sel_o[0]), .B(n4331), .S0(n3054), .Y(n4330)
         );
  INV_X0P5B_A12TR u5268 ( .A(n3221), .Y(n3054) );
  NOR2_X0P5A_A12TR u5269 ( .A(wtblat[0]), .B(n4305), .Y(n4331) );
  OAI222_X0P5M_A12TR u5270 ( .A0(n3572), .A1(n4332), .B0(n4333), .B1(n4334), 
        .C0(n3470), .C1(n4335), .Y(n1469) );
  INV_X0P5B_A12TR u5271 ( .A(iwb_dat_o[15]), .Y(n4334) );
  INV_X0P5B_A12TR u5272 ( .A(rilat[7]), .Y(n3572) );
  OAI222_X0P5M_A12TR u5273 ( .A0(n3571), .A1(n4332), .B0(n4333), .B1(n4336), 
        .C0(n3468), .C1(n4335), .Y(n1468) );
  INV_X0P5B_A12TR u5274 ( .A(iwb_dat_o[14]), .Y(n4336) );
  INV_X0P5B_A12TR u5275 ( .A(rilat[6]), .Y(n3571) );
  OAI222_X0P5M_A12TR u5276 ( .A0(n3570), .A1(n4332), .B0(n4333), .B1(n3667), 
        .C0(n3466), .C1(n4335), .Y(n1467) );
  INV_X0P5B_A12TR u5277 ( .A(dwb_dat_o[5]), .Y(n3466) );
  INV_X0P5B_A12TR u5278 ( .A(iwb_dat_o[13]), .Y(n3667) );
  INV_X0P5B_A12TR u5279 ( .A(rilat[5]), .Y(n3570) );
  OAI222_X0P5M_A12TR u5280 ( .A0(n3569), .A1(n4332), .B0(n4333), .B1(n4337), 
        .C0(n3148), .C1(n4335), .Y(n1466) );
  INV_X0P5B_A12TR u5281 ( .A(iwb_dat_o[12]), .Y(n4337) );
  INV_X0P5B_A12TR u5282 ( .A(rilat[4]), .Y(n3569) );
  OAI222_X0P5M_A12TR u5283 ( .A0(n3568), .A1(n4332), .B0(n4333), .B1(n4338), 
        .C0(n3458), .C1(n4335), .Y(n1465) );
  INV_X0P5B_A12TR u5284 ( .A(dwb_dat_o[3]), .Y(n3458) );
  INV_X0P5B_A12TR u5285 ( .A(iwb_dat_o[11]), .Y(n4338) );
  INV_X0P5B_A12TR u5286 ( .A(rilat[3]), .Y(n3568) );
  OAI222_X0P5M_A12TR u5287 ( .A0(n3567), .A1(n4332), .B0(n4333), .B1(n4339), 
        .C0(n3158), .C1(n4335), .Y(n1464) );
  INV_X0P5B_A12TR u5288 ( .A(iwb_dat_o[10]), .Y(n4339) );
  INV_X0P5B_A12TR u5289 ( .A(rilat[2]), .Y(n3567) );
  OAI222_X0P5M_A12TR u5290 ( .A0(n3566), .A1(n4332), .B0(n4333), .B1(n4340), 
        .C0(n3453), .C1(n4335), .Y(n1463) );
  INV_X0P5B_A12TR u5291 ( .A(iwb_dat_o[9]), .Y(n4340) );
  INV_X0P5B_A12TR u5292 ( .A(rilat[1]), .Y(n3566) );
  OAI222_X0P5M_A12TR u5293 ( .A0(n3565), .A1(n4332), .B0(n4333), .B1(n4341), 
        .C0(n3067), .C1(n4335), .Y(n1462) );
  NAND3_X0P5A_A12TR u5294 ( .A(n3109), .B(n4342), .C(n3646), .Y(n4335) );
  INV_X0P5B_A12TR u5295 ( .A(n3666), .Y(n3109) );
  INV_X0P5B_A12TR u5296 ( .A(iwb_dat_o[8]), .Y(n4341) );
  OA21A1OI2_X0P5M_A12TR u5297 ( .A0(n3666), .A1(n3597), .B0(n4342), .C0(n4237), 
        .Y(n4333) );
  NAND2_X0P5A_A12TR u5298 ( .A(n3677), .B(n3263), .Y(n3666) );
  AND3_X0P5M_A12TR u5299 ( .A(n4343), .B(n3679), .C(dwb_adr_o[2]), .Y(n3677)
         );
  INV_X0P5B_A12TR u5300 ( .A(dwb_adr_o[3]), .Y(n3679) );
  OR2_X0P5M_A12TR u5301 ( .A(n4342), .B(n4237), .Y(n4332) );
  NAND2_X0P5A_A12TR u5302 ( .A(rmxtbl[3]), .B(n4051), .Y(n4342) );
  INV_X0P5B_A12TR u5303 ( .A(rmxtbl[2]), .Y(n4051) );
  INV_X0P5B_A12TR u5304 ( .A(rilat[0]), .Y(n3565) );
  OAI22_X0P5M_A12TR u5305 ( .A0(qena[3]), .A1(n4344), .B0(n4345), .B1(n3776), 
        .Y(n1461) );
  OAI222_X0P5M_A12TR u5306 ( .A0(n3148), .A1(n4297), .B0(n4345), .B1(n4299), 
        .C0(n4254), .C1(n4344), .Y(n1459) );
  INV_X0P5B_A12TR u5307 ( .A(rpcu_4_), .Y(n4344) );
  INV_X0P5B_A12TR u5308 ( .A(rpclatu[4]), .Y(n4345) );
  INV_X0P5B_A12TR u5309 ( .A(dwb_dat_o[4]), .Y(n3148) );
  NAND4_X0P5A_A12TR u5310 ( .A(n4346), .B(n4347), .C(n4348), .D(n4349), .Y(
        n1458) );
  AOI222_X0P5M_A12TR u5311 ( .A0(wfsrplusw1[7]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[7]), .C0(n3815), .C1(wfsrinc2[7]), .Y(n4349) );
  AOI222_X0P5M_A12TR u5312 ( .A0(n3724), .A1(rfsr0l[7]), .B0(wfsrplusw2[7]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[7]), .Y(n4348) );
  AOI222_X0P5M_A12TR u5313 ( .A0(n3723), .A1(rfsr2l[7]), .B0(wfsrplusw0[7]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[7]), .Y(n4347) );
  AOI222_X0P5M_A12TR u5314 ( .A0(dwb_adr_o[7]), .A1(n3819), .B0(n3820), .B1(
        rromlat[7]), .C0(reaptr[7]), .C1(n3821), .Y(n4346) );
  NAND4_X0P5A_A12TR u5315 ( .A(n4350), .B(n4351), .C(n4352), .D(n4353), .Y(
        n1456) );
  AOI222_X0P5M_A12TR u5316 ( .A0(wfsrplusw1[8]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[8]), .C0(n3815), .C1(wfsrinc2[8]), .Y(n4353) );
  AOI222_X0P5M_A12TR u5317 ( .A0(n3724), .A1(rfsr0h[0]), .B0(wfsrplusw2[8]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[8]), .Y(n4352) );
  AOI222_X0P5M_A12TR u5318 ( .A0(n3723), .A1(rfsr2h[0]), .B0(wfsrplusw0[8]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1h[0]), .Y(n4351) );
  AOI222_X0P5M_A12TR u5319 ( .A0(dwb_adr_o[8]), .A1(n3819), .B0(n3820), .B1(
        rromlat[8]), .C0(n3821), .C1(reaptr[8]), .Y(n4350) );
  NAND4_X0P5A_A12TR u5320 ( .A(n4354), .B(n4355), .C(n4356), .D(n4357), .Y(
        n1454) );
  AOI222_X0P5M_A12TR u5321 ( .A0(wfsrplusw1[9]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[9]), .C0(n3815), .C1(wfsrinc2[9]), .Y(n4357) );
  AOI222_X0P5M_A12TR u5322 ( .A0(n3724), .A1(rfsr0h[1]), .B0(wfsrplusw2[9]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[9]), .Y(n4356) );
  AOI222_X0P5M_A12TR u5323 ( .A0(n3723), .A1(rfsr2h[1]), .B0(wfsrplusw0[9]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1h[1]), .Y(n4355) );
  AOI222_X0P5M_A12TR u5324 ( .A0(dwb_adr_o[9]), .A1(n3819), .B0(n3820), .B1(
        rromlat[9]), .C0(n3821), .C1(reaptr[9]), .Y(n4354) );
  NAND4_X0P5A_A12TR u5325 ( .A(n4358), .B(n4359), .C(n4360), .D(n4361), .Y(
        n1452) );
  AOI222_X0P5M_A12TR u5326 ( .A0(wfsrplusw1[10]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[10]), .C0(n3815), .C1(wfsrinc2[10]), .Y(n4361) );
  AOI222_X0P5M_A12TR u5327 ( .A0(n3724), .A1(rfsr0h[2]), .B0(wfsrplusw2[10]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[10]), .Y(n4360) );
  AOI222_X0P5M_A12TR u5328 ( .A0(n3723), .A1(rfsr2h[2]), .B0(wfsrplusw0[10]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1h[2]), .Y(n4359) );
  AOI222_X0P5M_A12TR u5329 ( .A0(dwb_adr_o[10]), .A1(n3819), .B0(n3820), .B1(
        rromlat[10]), .C0(n3821), .C1(reaptr[10]), .Y(n4358) );
  NAND4_X0P5A_A12TR u5330 ( .A(n4362), .B(n4363), .C(n4364), .D(n4365), .Y(
        n1450) );
  AOI222_X0P5M_A12TR u5331 ( .A0(wfsrplusw1[11]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[11]), .C0(n3815), .C1(wfsrinc2[11]), .Y(n4365) );
  AOI222_X0P5M_A12TR u5332 ( .A0(n3724), .A1(rfsr0h[3]), .B0(wfsrplusw2[11]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[11]), .Y(n4364) );
  AOI222_X0P5M_A12TR u5333 ( .A0(n3723), .A1(rfsr2h[3]), .B0(wfsrplusw0[11]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1h[3]), .Y(n4363) );
  AOI222_X0P5M_A12TR u5334 ( .A0(dwb_adr_o[11]), .A1(n3819), .B0(n3820), .B1(
        rromlat[11]), .C0(n3821), .C1(reaptr[11]), .Y(n4362) );
  NAND4_X0P5A_A12TR u5335 ( .A(n4366), .B(n4367), .C(n4368), .D(n4369), .Y(
        n1448) );
  AOI222_X0P5M_A12TR u5336 ( .A0(wfsrplusw1[6]), .A1(n3813), .B0(n3814), .B1(
        wfsrinc0[6]), .C0(n3815), .C1(wfsrinc2[6]), .Y(n4369) );
  AND3_X0P5M_A12TR u5337 ( .A(n3463), .B(n3554), .C(n4370), .Y(n3815) );
  AND2_X0P5M_A12TR u5338 ( .A(n4371), .B(n3484), .Y(n3814) );
  AND3_X0P5M_A12TR u5339 ( .A(n3484), .B(rmxfsr[2]), .C(n4370), .Y(n3813) );
  NOR3_X0P5A_A12TR u5340 ( .A(rmxfsr[0]), .B(rmxfsr[3]), .C(n3528), .Y(n3484)
         );
  AOI222_X0P5M_A12TR u5341 ( .A0(n3724), .A1(rfsr0l[6]), .B0(wfsrplusw2[6]), 
        .B1(n3816), .C0(n3817), .C1(wfsrinc1[6]), .Y(n4368) );
  INV_X0P5B_A12TR u5342 ( .A(n3527), .Y(n3817) );
  NAND4_X0P5A_A12TR u5343 ( .A(n4370), .B(n3462), .C(rmxfsr[2]), .D(n3479), 
        .Y(n3527) );
  AND3_X0P5M_A12TR u5344 ( .A(n3462), .B(rmxfsr[3]), .C(n4371), .Y(n3816) );
  AND3_X0P5M_A12TR u5345 ( .A(n4370), .B(n3479), .C(n4372), .Y(n3724) );
  MXIT2_X0P5M_A12TR u5346 ( .A(rmxfsr[1]), .B(n3482), .S0(n3483), .Y(n4372) );
  AOI222_X0P5M_A12TR u5347 ( .A0(n3723), .A1(rfsr2l[6]), .B0(wfsrplusw0[6]), 
        .B1(n3818), .C0(n3725), .C1(rfsr1l[6]), .Y(n4367) );
  AND3_X0P5M_A12TR u5348 ( .A(rmxfsr[3]), .B(n3482), .C(n4371), .Y(n3725) );
  INV_X0P5B_A12TR u5349 ( .A(n3462), .Y(n3482) );
  NOR2_X0P5A_A12TR u5350 ( .A(n3528), .B(n3543), .Y(n3462) );
  INV_X0P5B_A12TR u5351 ( .A(rmxfsr[0]), .Y(n3543) );
  AND4_X0P5M_A12TR u5352 ( .A(n4371), .B(rmxfsr[0]), .C(n3528), .D(n3479), .Y(
        n3818) );
  INV_X0P5B_A12TR u5353 ( .A(rmxfsr[1]), .Y(n3528) );
  AND3_X0P5M_A12TR u5354 ( .A(n3554), .B(n3481), .C(n4370), .Y(n3723) );
  INV_X0P5B_A12TR u5355 ( .A(n3463), .Y(n3481) );
  NOR2_X0P5A_A12TR u5356 ( .A(n3479), .B(n3483), .Y(n3554) );
  INV_X0P5B_A12TR u5357 ( .A(rmxfsr[2]), .Y(n3483) );
  AOI222_X0P5M_A12TR u5358 ( .A0(dwb_adr_o[6]), .A1(n3819), .B0(n3820), .B1(
        rromlat[6]), .C0(reaptr[6]), .C1(n3821), .Y(n4366) );
  INV_X0P5B_A12TR u5359 ( .A(n3719), .Y(n3821) );
  NAND3_X0P5A_A12TR u5360 ( .A(n3463), .B(n3479), .C(n4371), .Y(n3719) );
  NOR2_X0P5A_A12TR u5361 ( .A(n3928), .B(rmxfsr[2]), .Y(n4371) );
  INV_X0P5B_A12TR u5362 ( .A(n4370), .Y(n3928) );
  NOR2_X0P5A_A12TR u5363 ( .A(n3138), .B(n3476), .Y(n4370) );
  INV_X0P5B_A12TR u5364 ( .A(n3143), .Y(n3138) );
  NOR2_X0P5A_A12TR u5365 ( .A(qfsm[0]), .B(qfsm[1]), .Y(n3143) );
  INV_X0P5B_A12TR u5366 ( .A(rmxfsr[3]), .Y(n3479) );
  NOR2_X0P5A_A12TR u5367 ( .A(rmxfsr[0]), .B(rmxfsr[1]), .Y(n3463) );
  AND4_X0P5M_A12TR u5368 ( .A(n4373), .B(rmxbsr[0]), .C(n3460), .D(n3242), .Y(
        n3820) );
  NOR2_X0P5A_A12TR u5369 ( .A(n4305), .B(qfsm[1]), .Y(n3460) );
  INV_X0P5B_A12TR u5370 ( .A(rmxbsr[1]), .Y(n4373) );
  NAND2_X0P5A_A12TR u5371 ( .A(n4374), .B(n3242), .Y(n3819) );
  OA21A1OI2_X0P5M_A12TR u5372 ( .A0(rmxbsr[1]), .A1(n3406), .B0(qfsm[0]), .C0(
        qfsm[1]), .Y(n4374) );
  INV_X0P5B_A12TR u5373 ( .A(rmxbsr[0]), .Y(n3406) );
  OAI222_X0P5M_A12TR u5374 ( .A0(n3468), .A1(n3776), .B0(n4375), .B1(n3778), 
        .C0(qena[3]), .C1(n4376), .Y(n1446) );
  INV_X0P5B_A12TR u5375 ( .A(wpclat[5]), .Y(n4376) );
  OAI221_X0P5M_A12TR u5376 ( .A0(n3064), .A1(n4377), .B0(n3066), .B1(n3468), 
        .C0(n4378), .Y(n1444) );
  AOI22_X0P5M_A12TR u5377 ( .A0(n2758), .A1(n3069), .B0(n3871), .B1(wpclat[5]), 
        .Y(n4378) );
  INV_X0P5B_A12TR u5378 ( .A(dwb_dat_o[6]), .Y(n3468) );
  NAND2_X0P5A_A12TR u5379 ( .A(n3110), .B(n4379), .Y(n3066) );
  INV_X0P5B_A12TR u5380 ( .A(n3668), .Y(n3110) );
  INV_X0P5B_A12TR u5381 ( .A(wstkw[6]), .Y(n4377) );
  AOI21_X0P5M_A12TR u5382 ( .A0(n3668), .A1(n4380), .B0(n4381), .Y(n3064) );
  NAND2_X0P5A_A12TR u5383 ( .A(n4382), .B(n3263), .Y(n3668) );
  OAI211_X0P5M_A12TR u5384 ( .A0(qena[1]), .A1(n4375), .B0(n4383), .C0(n4384), 
        .Y(n1443) );
  AOI222_X0P5M_A12TR u5385 ( .A0(wpcinc[5]), .A1(n3792), .B0(n391), .B1(n3793), 
        .C0(n3794), .C1(wstkw[6]), .Y(n4384) );
  AOI22_X0P5M_A12TR u5386 ( .A0(n371), .A1(n3795), .B0(n3796), .B1(rireg[5]), 
        .Y(n4383) );
  INV_X0P5B_A12TR u5387 ( .A(rpcnxt[5]), .Y(n4375) );
  OAI211_X0P5M_A12TR u5388 ( .A0(qena[1]), .A1(n4385), .B0(n4386), .C0(n4387), 
        .Y(n1440) );
  AOI222_X0P5M_A12TR u5389 ( .A0(wpcinc[14]), .A1(n3792), .B0(n400), .B1(n3793), .C0(n3794), .C1(wstkw[15]), .Y(n4387) );
  AOI22_X0P5M_A12TR u5390 ( .A0(n380), .A1(n3795), .B0(n3796), .B1(rromlat[6]), 
        .Y(n4386) );
  OAI222_X0P5M_A12TR u5391 ( .A0(n4388), .A1(n3776), .B0(n4385), .B1(n3778), 
        .C0(qena[3]), .C1(n4389), .Y(n1437) );
  INV_X0P5B_A12TR u5392 ( .A(rpcnxt[14]), .Y(n4385) );
  OAI222_X0P5M_A12TR u5393 ( .A0(n3470), .A1(n4252), .B0(n4388), .B1(n4253), 
        .C0(n4254), .C1(n4389), .Y(n1435) );
  INV_X0P5B_A12TR u5394 ( .A(wpclat[14]), .Y(n4389) );
  NAND2_X0P5A_A12TR u5395 ( .A(n4254), .B(n4252), .Y(n4253) );
  INV_X0P5B_A12TR u5396 ( .A(rpclath[7]), .Y(n4388) );
  NAND2_X0P5A_A12TR u5397 ( .A(n3646), .B(n3108), .Y(n4252) );
  AND2_X0P5M_A12TR u5398 ( .A(n4306), .B(n3676), .Y(n3108) );
  OAI221_X0P5M_A12TR u5399 ( .A0(n3907), .A1(n4390), .B0(n3470), .B1(n3909), 
        .C0(n4391), .Y(n1434) );
  AOI22_X0P5M_A12TR u5400 ( .A0(n2759), .A1(n3069), .B0(wpclat[14]), .B1(n3871), .Y(n4391) );
  NAND2_X0P5A_A12TR u5401 ( .A(n3102), .B(n4379), .Y(n3909) );
  INV_X0P5B_A12TR u5402 ( .A(n4392), .Y(n3102) );
  INV_X0P5B_A12TR u5403 ( .A(dwb_dat_o[7]), .Y(n3470) );
  INV_X0P5B_A12TR u5404 ( .A(wstkw[15]), .Y(n4390) );
  AOI21_X0P5M_A12TR u5405 ( .A0(n4392), .A1(n4380), .B0(n4381), .Y(n3907) );
  NAND2_X0P5A_A12TR u5406 ( .A(n3676), .B(n4382), .Y(n4392) );
  NOR2_X0P5A_A12TR u5407 ( .A(n3732), .B(dwb_adr_o[0]), .Y(n3676) );
  OAI211_X0P5M_A12TR u5408 ( .A0(qena[1]), .A1(n4393), .B0(n4394), .C0(n4395), 
        .Y(n1433) );
  AOI222_X0P5M_A12TR u5409 ( .A0(wpcinc[15]), .A1(n3792), .B0(n401), .B1(n3793), .C0(n3794), .C1(wstkw[16]), .Y(n4395) );
  AOI22_X0P5M_A12TR u5410 ( .A0(n381), .A1(n3795), .B0(n3796), .B1(rromlat[7]), 
        .Y(n4394) );
  OAI222_X0P5M_A12TR u5411 ( .A0(n4396), .A1(n3776), .B0(n4393), .B1(n3778), 
        .C0(qena[3]), .C1(n4397), .Y(n1430) );
  INV_X0P5B_A12TR u5412 ( .A(rpcnxt[15]), .Y(n4393) );
  OAI222_X0P5M_A12TR u5413 ( .A0(n3067), .A1(n4297), .B0(n4396), .B1(n4299), 
        .C0(n4254), .C1(n4397), .Y(n1428) );
  INV_X0P5B_A12TR u5414 ( .A(wpclat[15]), .Y(n4397) );
  INV_X0P5B_A12TR u5415 ( .A(rpclatu[0]), .Y(n4396) );
  OAI221_X0P5M_A12TR u5416 ( .A0(n3879), .A1(n4398), .B0(n3067), .B1(n3880), 
        .C0(n4399), .Y(n1427) );
  AOI22_X0P5M_A12TR u5417 ( .A0(n2760), .A1(n3069), .B0(wpclat[15]), .B1(n3871), .Y(n4399) );
  INV_X0P5B_A12TR u5418 ( .A(dwb_dat_o[0]), .Y(n3067) );
  INV_X0P5B_A12TR u5419 ( .A(wstkw[16]), .Y(n4398) );
  OAI211_X0P5M_A12TR u5420 ( .A0(qena[1]), .A1(n4400), .B0(n4401), .C0(n4402), 
        .Y(n1426) );
  AOI222_X0P5M_A12TR u5421 ( .A0(wpcinc[16]), .A1(n3792), .B0(n402), .B1(n3793), .C0(n3794), .C1(wstkw[17]), .Y(n4402) );
  NOR3_X0P5A_A12TR u5422 ( .A(rmxnpc[1]), .B(rmxnpc[2]), .C(n4251), .Y(n3794)
         );
  AND4_X0P5M_A12TR u5423 ( .A(rmxnpc[1]), .B(n3738), .C(n4053), .D(n3937), .Y(
        n3793) );
  INV_X0P5B_A12TR u5424 ( .A(rmxnpc[2]), .Y(n3937) );
  OA21_X0P5M_A12TR u5425 ( .A0(n4403), .A1(n4404), .B0(qena[1]), .Y(n3792) );
  MXIT2_X0P5M_A12TR u5426 ( .A(n4405), .B(rmxnpc[1]), .S0(n4053), .Y(n4404) );
  NAND2_X0P5A_A12TR u5427 ( .A(n4209), .B(n3716), .Y(n4405) );
  INV_X0P5B_A12TR u5428 ( .A(n4406), .Y(n4209) );
  OA21A1OI2_X0P5M_A12TR u5429 ( .A0(n4001), .A1(n4053), .B0(rmxnpc[2]), .C0(
        rnskp), .Y(n4403) );
  INV_X0P5B_A12TR u5430 ( .A(rmxnpc[0]), .Y(n4053) );
  AOI22_X0P5M_A12TR u5431 ( .A0(n382), .A1(n3795), .B0(n3796), .B1(rromlat[8]), 
        .Y(n4401) );
  NOR3_X0P5A_A12TR u5432 ( .A(n4001), .B(rmxnpc[2]), .C(n4251), .Y(n3796) );
  INV_X0P5B_A12TR u5433 ( .A(rmxnpc[1]), .Y(n4001) );
  NOR3_X0P5A_A12TR u5434 ( .A(n4251), .B(n3716), .C(n4406), .Y(n3795) );
  NAND2_X0P5A_A12TR u5435 ( .A(rmxnpc[2]), .B(rmxnpc[1]), .Y(n4406) );
  INV_X0P5B_A12TR u5436 ( .A(rbcc), .Y(n3716) );
  NAND2_X0P5A_A12TR u5437 ( .A(rmxnpc[0]), .B(n3738), .Y(n4251) );
  NOR2_X0P5A_A12TR u5438 ( .A(n3375), .B(n3708), .Y(n3738) );
  INV_X0P5B_A12TR u5439 ( .A(qena[1]), .Y(n3375) );
  OAI222_X0P5M_A12TR u5440 ( .A0(n4407), .A1(n3776), .B0(n4400), .B1(n3778), 
        .C0(qena[3]), .C1(n4408), .Y(n1423) );
  INV_X0P5B_A12TR u5441 ( .A(rpcnxt[16]), .Y(n4400) );
  OAI222_X0P5M_A12TR u5442 ( .A0(n3453), .A1(n4297), .B0(n4407), .B1(n4299), 
        .C0(n4254), .C1(n4408), .Y(n1421) );
  INV_X0P5B_A12TR u5443 ( .A(wpclat[16]), .Y(n4408) );
  INV_X0P5B_A12TR u5444 ( .A(rpclatu[1]), .Y(n4407) );
  OAI221_X0P5M_A12TR u5445 ( .A0(n3879), .A1(n3276), .B0(n3453), .B1(n3880), 
        .C0(n4409), .Y(n1420) );
  AOI22_X0P5M_A12TR u5446 ( .A0(n2781), .A1(n3069), .B0(wpclat[16]), .B1(n3871), .Y(n4409) );
  INV_X0P5B_A12TR u5447 ( .A(wstkw[17]), .Y(n3276) );
  OAI222_X0P5M_A12TR u5448 ( .A0(n4410), .A1(n3776), .B0(n3899), .B1(n3778), 
        .C0(qena[3]), .C1(n4411), .Y(n1419) );
  OAI21_X0P5M_A12TR u5449 ( .A0(n3597), .A1(n3662), .B0(qena[3]), .Y(n3778) );
  INV_X0P5B_A12TR u5450 ( .A(rpcnxt[17]), .Y(n3899) );
  INV_X0P5B_A12TR u5451 ( .A(n3709), .Y(n3776) );
  NOR3_X0P5A_A12TR u5452 ( .A(n3074), .B(n3597), .C(n3662), .Y(n3709) );
  OAI222_X0P5M_A12TR u5453 ( .A0(n3158), .A1(n4297), .B0(n4410), .B1(n4299), 
        .C0(n4254), .C1(n4411), .Y(n1417) );
  INV_X0P5B_A12TR u5454 ( .A(wpclat[17]), .Y(n4411) );
  NAND2_X0P5A_A12TR u5455 ( .A(n4254), .B(n4297), .Y(n4299) );
  NAND4B_X0P5M_A12TR u5456 ( .AN(n3726), .B(n3688), .C(n3101), .D(n4118), .Y(
        n4254) );
  INV_X0P5B_A12TR u5457 ( .A(n3662), .Y(n3101) );
  NAND2_X0P5A_A12TR u5458 ( .A(n4306), .B(n3263), .Y(n3662) );
  NOR2_X0P5A_A12TR u5459 ( .A(n3733), .B(dwb_adr_o[1]), .Y(n3263) );
  INV_X0P5B_A12TR u5460 ( .A(rpclatu[2]), .Y(n4410) );
  NAND2_X0P5A_A12TR u5461 ( .A(n3646), .B(n3103), .Y(n4297) );
  AND2_X0P5M_A12TR u5462 ( .A(n4306), .B(n3678), .Y(n3103) );
  AND3_X0P5M_A12TR u5463 ( .A(n4343), .B(n3683), .C(dwb_adr_o[3]), .Y(n4306)
         );
  INV_X0P5B_A12TR u5464 ( .A(dwb_adr_o[2]), .Y(n3683) );
  NOR2_X0P5A_A12TR u5465 ( .A(n4237), .B(n3597), .Y(n3646) );
  OAI221_X0P5M_A12TR u5466 ( .A0(n3879), .A1(n3291), .B0(n3158), .B1(n3880), 
        .C0(n4412), .Y(n1416) );
  AOI22_X0P5M_A12TR u5467 ( .A0(n2780), .A1(n3069), .B0(wpclat[17]), .B1(n3871), .Y(n4412) );
  NAND2_X0P5A_A12TR u5468 ( .A(n3270), .B(n4379), .Y(n3880) );
  INV_X0P5B_A12TR u5469 ( .A(n3096), .Y(n3270) );
  INV_X0P5B_A12TR u5470 ( .A(dwb_dat_o[2]), .Y(n3158) );
  INV_X0P5B_A12TR u5471 ( .A(wstkw[18]), .Y(n3291) );
  AOI21_X0P5M_A12TR u5472 ( .A0(n3096), .A1(n4380), .B0(n4381), .Y(n3879) );
  OAI21_X0P5M_A12TR u5473 ( .A0(n3240), .A1(n4413), .B0(n4414), .Y(n4381) );
  INV_X0P5B_A12TR u5474 ( .A(n4413), .Y(n4380) );
  NAND2_X0P5A_A12TR u5475 ( .A(n4415), .B(n4416), .Y(n4413) );
  NAND2_X0P5A_A12TR u5476 ( .A(n3678), .B(n4382), .Y(n3096) );
  NOR2_X0P5A_A12TR u5477 ( .A(n3732), .B(n3733), .Y(n3678) );
  INV_X0P5B_A12TR u5478 ( .A(dwb_adr_o[0]), .Y(n3733) );
  INV_X0P5B_A12TR u5479 ( .A(dwb_adr_o[1]), .Y(n3732) );
  OAI221_X0P5M_A12TR u5480 ( .A0(n3844), .A1(n3851), .B0(n3453), .B1(n3843), 
        .C0(n4417), .Y(n1415) );
  AOI22_X0P5M_A12TR u5481 ( .A0(n215), .A1(n3840), .B0(wstkdec[1]), .B1(n3855), 
        .Y(n4417) );
  INV_X0P5B_A12TR u5482 ( .A(n3842), .Y(n3855) );
  NAND2_X0P5A_A12TR u5483 ( .A(n3069), .B(n3324), .Y(n3842) );
  INV_X0P5B_A12TR u5484 ( .A(rstkunf), .Y(n3324) );
  NOR2B_X0P5M_A12TR u5485 ( .AN(n4414), .B(n4416), .Y(n3069) );
  AO21A1AI2_X0P5M_A12TR u5486 ( .A0(n3269), .A1(n3240), .B0(n4418), .C0(n4414), 
        .Y(n3840) );
  OAI22_X0P5M_A12TR u5487 ( .A0(rstkful), .A1(n4415), .B0(rstkunf), .B1(n4416), 
        .Y(n4418) );
  NAND3B_X0P5M_A12TR u5488 ( .AN(rmxstk[1]), .B(n4305), .C(rmxstk[0]), .Y(
        n4416) );
  NAND2_X0P5A_A12TR u5489 ( .A(n3269), .B(n4379), .Y(n3843) );
  AND2_X0P5M_A12TR u5490 ( .A(n3240), .B(n4414), .Y(n4379) );
  NOR2_X0P5A_A12TR u5491 ( .A(n4305), .B(n3597), .Y(n3240) );
  INV_X0P5B_A12TR u5492 ( .A(n3645), .Y(n3597) );
  NOR2_X0P5A_A12TR u5493 ( .A(n4118), .B(n3726), .Y(n3645) );
  NAND4B_X0P5M_A12TR u5494 ( .AN(n4419), .B(rdwbadr[15]), .C(rdwbadr[14]), .D(
        n4420), .Y(n3726) );
  AND3_X0P5M_A12TR u5495 ( .A(rdwbadr[13]), .B(dwb_adr_o[9]), .C(rdwbadr[12]), 
        .Y(n4420) );
  NAND3B_X0P5M_A12TR u5496 ( .AN(n4421), .B(dwb_adr_o[7]), .C(dwb_adr_o[8]), 
        .Y(n4419) );
  NAND3_X0P5A_A12TR u5497 ( .A(dwb_adr_o[11]), .B(dwb_adr_o[10]), .C(
        dwb_adr_o[6]), .Y(n4421) );
  INV_X0P5B_A12TR u5498 ( .A(dwb_we_o), .Y(n4118) );
  INV_X0P5B_A12TR u5499 ( .A(n3098), .Y(n3269) );
  NAND2_X0P5A_A12TR u5500 ( .A(n3317), .B(n4382), .Y(n3098) );
  AND3_X0P5M_A12TR u5501 ( .A(dwb_adr_o[2]), .B(n4343), .C(dwb_adr_o[3]), .Y(
        n4382) );
  NOR2_X0P5A_A12TR u5502 ( .A(n3684), .B(n3734), .Y(n4343) );
  INV_X0P5B_A12TR u5503 ( .A(dwb_adr_o[4]), .Y(n3734) );
  INV_X0P5B_A12TR u5504 ( .A(dwb_adr_o[5]), .Y(n3684) );
  NOR2_X0P5A_A12TR u5505 ( .A(dwb_adr_o[0]), .B(dwb_adr_o[1]), .Y(n3317) );
  INV_X0P5B_A12TR u5506 ( .A(dwb_dat_o[1]), .Y(n3453) );
  INV_X0P5B_A12TR u5507 ( .A(wstkinc[1]), .Y(n3851) );
  NAND2_X0P5A_A12TR u5508 ( .A(n3871), .B(n3099), .Y(n3844) );
  INV_X0P5B_A12TR u5509 ( .A(rstkful), .Y(n3099) );
  NOR2B_X0P5M_A12TR u5510 ( .AN(n4414), .B(n4415), .Y(n3871) );
  NAND3B_X0P5M_A12TR u5511 ( .AN(rmxstk[0]), .B(n4305), .C(rmxstk[1]), .Y(
        n4415) );
  INV_X0P5B_A12TR u5512 ( .A(qfsm[0]), .Y(n4305) );
  NOR2_X0P5A_A12TR u5513 ( .A(n4119), .B(n3476), .Y(n4414) );
  INV_X0P5B_A12TR u5514 ( .A(n3242), .Y(n3476) );
  NOR2_X0P5A_A12TR u5515 ( .A(n3708), .B(n3221), .Y(n3242) );
  NOR2_X0P5A_A12TR u5516 ( .A(n3223), .B(n3226), .Y(n3221) );
  INV_X0P5B_A12TR u5517 ( .A(rfsm[0]), .Y(n3226) );
  INV_X0P5B_A12TR u5518 ( .A(rfsm[1]), .Y(n3223) );
  INV_X0P5B_A12TR u5519 ( .A(qfsm[1]), .Y(n4119) );
  MXIT2_X0P5M_A12TR u5520 ( .A(n3146), .B(n3141), .S0(n4127), .Y(n1414) );
  INV_X0P5B_A12TR u5521 ( .A(rn), .Y(n3141) );
  INV_X0P5B_A12TR u5522 ( .A(rstatus_[4]), .Y(n3146) );
  MXT2_X0P5M_A12TR u5523 ( .A(rstatus_[1]), .B(rdc), .S0(n4127), .Y(n1413) );
  AND3_X0P5M_A12TR u5524 ( .A(n3688), .B(n4238), .C(rmxsha[1]), .Y(n4127) );
  INV_X0P5B_A12TR u5525 ( .A(rmxsha[0]), .Y(n4238) );
  AND2_X0P5M_A12TR u5526 ( .A(rsleep_), .B(n3688), .Y(n846) );
  NOR2_X0P5A_A12TR u5527 ( .A(n4237), .B(n4117), .Y(n845) );
  INV_X0P5B_A12TR u5528 ( .A(rclrwdt_), .Y(n4117) );
  INV_X0P5B_A12TR u5529 ( .A(n3688), .Y(n4237) );
  NOR2_X0P5A_A12TR u5530 ( .A(n3074), .B(n3708), .Y(n3688) );
  INV_X0P5B_A12TR u5531 ( .A(rnskp), .Y(n3708) );
  INV_X0P5B_A12TR u5532 ( .A(qena[3]), .Y(n3074) );
  XOR3_X0P5M_A12TR u5533 ( .A(rprng[4]), .B(n4422), .C(rprng[3]), .Y(n262) );
  XOR2_X0P5M_A12TR u5534 ( .A(rprng[7]), .B(rprng[5]), .Y(n4422) );
  OR2_X1M_A12TR sub_1479_u22 ( .A(sub_1479_n2), .B(rfsr2h[2]), .Y(sub_1479_n10) );
  OR2_X1M_A12TR sub_1479_u21 ( .A(sub_1479_n7), .B(rfsr2l[3]), .Y(sub_1479_n9)
         );
  OR2_X1M_A12TR sub_1479_u20 ( .A(sub_1479_n3), .B(rfsr2l[5]), .Y(sub_1479_n8)
         );
  OR2_X1M_A12TR sub_1479_u19 ( .A(sub_1479_n6), .B(rfsr2l[2]), .Y(sub_1479_n7)
         );
  OR2_X1M_A12TR sub_1479_u18 ( .A(rfsr2l[0]), .B(rfsr2l[1]), .Y(sub_1479_n6)
         );
  OR2_X1M_A12TR sub_1479_u17 ( .A(sub_1479_n8), .B(rfsr2l[6]), .Y(sub_1479_n5)
         );
  OR2_X1M_A12TR sub_1479_u16 ( .A(sub_1479_n5), .B(rfsr2l[7]), .Y(sub_1479_n4)
         );
  OR2_X1M_A12TR sub_1479_u15 ( .A(sub_1479_n9), .B(rfsr2l[4]), .Y(sub_1479_n3)
         );
  OR2_X1M_A12TR sub_1479_u14 ( .A(sub_1479_n1), .B(rfsr2h[1]), .Y(sub_1479_n2)
         );
  OR2_X1M_A12TR sub_1479_u13 ( .A(sub_1479_n4), .B(rfsr2h[0]), .Y(sub_1479_n1)
         );
  XNOR2_X1M_A12TR sub_1479_u12 ( .A(rfsr2l[1]), .B(rfsr2l[0]), .Y(wfsrdec2[1])
         );
  XNOR2_X1M_A12TR sub_1479_u11 ( .A(rfsr2l[4]), .B(sub_1479_n9), .Y(
        wfsrdec2[4]) );
  XNOR2_X1M_A12TR sub_1479_u10 ( .A(rfsr2l[6]), .B(sub_1479_n8), .Y(
        wfsrdec2[6]) );
  XNOR2_X1M_A12TR sub_1479_u9 ( .A(rfsr2l[3]), .B(sub_1479_n7), .Y(wfsrdec2[3]) );
  XNOR2_X1M_A12TR sub_1479_u8 ( .A(rfsr2l[2]), .B(sub_1479_n6), .Y(wfsrdec2[2]) );
  INV_X1M_A12TR sub_1479_u7 ( .A(rfsr2l[0]), .Y(wfsrdec2[0]) );
  XNOR2_X1M_A12TR sub_1479_u6 ( .A(rfsr2l[7]), .B(sub_1479_n5), .Y(wfsrdec2[7]) );
  XNOR2_X1M_A12TR sub_1479_u5 ( .A(rfsr2l[5]), .B(sub_1479_n3), .Y(wfsrdec2[5]) );
  XNOR2_X1M_A12TR sub_1479_u4 ( .A(rfsr2h[3]), .B(sub_1479_n10), .Y(
        wfsrdec2[11]) );
  XNOR2_X1M_A12TR sub_1479_u3 ( .A(rfsr2h[2]), .B(sub_1479_n2), .Y(
        wfsrdec2[10]) );
  XNOR2_X1M_A12TR sub_1479_u2 ( .A(rfsr2h[1]), .B(sub_1479_n1), .Y(wfsrdec2[9]) );
  XNOR2_X1M_A12TR sub_1479_u1 ( .A(rfsr2h[0]), .B(sub_1479_n4), .Y(wfsrdec2[8]) );
  OR2_X1M_A12TR sub_1552_u38 ( .A(sub_1552_n17), .B(wtblat[18]), .Y(
        sub_1552_n18) );
  OR2_X1M_A12TR sub_1552_u37 ( .A(sub_1552_n15), .B(wtblat[17]), .Y(
        sub_1552_n17) );
  OR2_X1M_A12TR sub_1552_u36 ( .A(sub_1552_n4), .B(wtblat[8]), .Y(sub_1552_n16) );
  OR2_X1M_A12TR sub_1552_u35 ( .A(sub_1552_n14), .B(wtblat[16]), .Y(
        sub_1552_n15) );
  OR2_X1M_A12TR sub_1552_u34 ( .A(sub_1552_n13), .B(wtblat[15]), .Y(
        sub_1552_n14) );
  OR2_X1M_A12TR sub_1552_u33 ( .A(sub_1552_n12), .B(wtblat[14]), .Y(
        sub_1552_n13) );
  OR2_X1M_A12TR sub_1552_u32 ( .A(sub_1552_n8), .B(wtblat[13]), .Y(
        sub_1552_n12) );
  OR2_X1M_A12TR sub_1552_u31 ( .A(sub_1552_n10), .B(wtblat[3]), .Y(
        sub_1552_n11) );
  OR2_X1M_A12TR sub_1552_u30 ( .A(sub_1552_n9), .B(wtblat[2]), .Y(sub_1552_n10) );
  OR2_X1M_A12TR sub_1552_u29 ( .A(wtblat[0]), .B(wtblat[1]), .Y(sub_1552_n9)
         );
  OR2_X1M_A12TR sub_1552_u28 ( .A(sub_1552_n7), .B(wtblat[12]), .Y(sub_1552_n8) );
  OR2_X1M_A12TR sub_1552_u27 ( .A(sub_1552_n6), .B(wtblat[11]), .Y(sub_1552_n7) );
  OR2_X1M_A12TR sub_1552_u26 ( .A(sub_1552_n5), .B(wtblat[10]), .Y(sub_1552_n6) );
  OR2_X1M_A12TR sub_1552_u25 ( .A(sub_1552_n16), .B(wtblat[9]), .Y(sub_1552_n5) );
  OR2_X1M_A12TR sub_1552_u24 ( .A(sub_1552_n3), .B(wtblat[7]), .Y(sub_1552_n4)
         );
  OR2_X1M_A12TR sub_1552_u23 ( .A(sub_1552_n2), .B(wtblat[6]), .Y(sub_1552_n3)
         );
  OR2_X1M_A12TR sub_1552_u22 ( .A(sub_1552_n1), .B(wtblat[5]), .Y(sub_1552_n2)
         );
  OR2_X1M_A12TR sub_1552_u21 ( .A(sub_1552_n11), .B(wtblat[4]), .Y(sub_1552_n1) );
  XNOR2_X1M_A12TR sub_1552_u20 ( .A(wtblat[17]), .B(sub_1552_n15), .Y(
        wtbldec[17]) );
  XNOR2_X1M_A12TR sub_1552_u19 ( .A(wtblat[19]), .B(sub_1552_n18), .Y(
        wtbldec[19]) );
  XNOR2_X1M_A12TR sub_1552_u18 ( .A(wtblat[18]), .B(sub_1552_n17), .Y(
        wtbldec[18]) );
  XNOR2_X1M_A12TR sub_1552_u17 ( .A(wtblat[16]), .B(sub_1552_n14), .Y(
        wtbldec[16]) );
  INV_X1M_A12TR sub_1552_u16 ( .A(wtblat[0]), .Y(wtbldec[0]) );
  XNOR2_X1M_A12TR sub_1552_u15 ( .A(wtblat[1]), .B(wtblat[0]), .Y(wtbldec[1])
         );
  XNOR2_X1M_A12TR sub_1552_u14 ( .A(wtblat[2]), .B(sub_1552_n9), .Y(wtbldec[2]) );
  XNOR2_X1M_A12TR sub_1552_u13 ( .A(wtblat[3]), .B(sub_1552_n10), .Y(
        wtbldec[3]) );
  XNOR2_X1M_A12TR sub_1552_u12 ( .A(wtblat[4]), .B(sub_1552_n11), .Y(
        wtbldec[4]) );
  XNOR2_X1M_A12TR sub_1552_u11 ( .A(wtblat[5]), .B(sub_1552_n1), .Y(wtbldec[5]) );
  XNOR2_X1M_A12TR sub_1552_u10 ( .A(wtblat[6]), .B(sub_1552_n2), .Y(wtbldec[6]) );
  XNOR2_X1M_A12TR sub_1552_u9 ( .A(wtblat[7]), .B(sub_1552_n3), .Y(wtbldec[7])
         );
  XNOR2_X1M_A12TR sub_1552_u8 ( .A(wtblat[8]), .B(sub_1552_n4), .Y(wtbldec[8])
         );
  XNOR2_X1M_A12TR sub_1552_u7 ( .A(wtblat[9]), .B(sub_1552_n16), .Y(wtbldec[9]) );
  XNOR2_X1M_A12TR sub_1552_u6 ( .A(wtblat[10]), .B(sub_1552_n5), .Y(
        wtbldec[10]) );
  XNOR2_X1M_A12TR sub_1552_u5 ( .A(wtblat[11]), .B(sub_1552_n6), .Y(
        wtbldec[11]) );
  XNOR2_X1M_A12TR sub_1552_u4 ( .A(wtblat[12]), .B(sub_1552_n7), .Y(
        wtbldec[12]) );
  XNOR2_X1M_A12TR sub_1552_u3 ( .A(wtblat[13]), .B(sub_1552_n8), .Y(
        wtbldec[13]) );
  XNOR2_X1M_A12TR sub_1552_u2 ( .A(wtblat[14]), .B(sub_1552_n12), .Y(
        wtbldec[14]) );
  XNOR2_X1M_A12TR sub_1552_u1 ( .A(wtblat[15]), .B(sub_1552_n13), .Y(
        wtbldec[15]) );
  OR2_X1M_A12TR sub_1478_u22 ( .A(sub_1478_n2), .B(rfsr1h[2]), .Y(sub_1478_n10) );
  OR2_X1M_A12TR sub_1478_u21 ( .A(sub_1478_n7), .B(rfsr1l[7]), .Y(sub_1478_n9)
         );
  OR2_X1M_A12TR sub_1478_u20 ( .A(sub_1478_n3), .B(rfsr1l[5]), .Y(sub_1478_n8)
         );
  OR2_X1M_A12TR sub_1478_u19 ( .A(sub_1478_n8), .B(rfsr1l[6]), .Y(sub_1478_n7)
         );
  OR2_X1M_A12TR sub_1478_u18 ( .A(rfsr1l[0]), .B(rfsr1l[1]), .Y(sub_1478_n6)
         );
  OR2_X1M_A12TR sub_1478_u17 ( .A(sub_1478_n6), .B(rfsr1l[2]), .Y(sub_1478_n5)
         );
  OR2_X1M_A12TR sub_1478_u16 ( .A(sub_1478_n5), .B(rfsr1l[3]), .Y(sub_1478_n4)
         );
  OR2_X1M_A12TR sub_1478_u15 ( .A(sub_1478_n4), .B(rfsr1l[4]), .Y(sub_1478_n3)
         );
  OR2_X1M_A12TR sub_1478_u14 ( .A(sub_1478_n1), .B(rfsr1h[1]), .Y(sub_1478_n2)
         );
  OR2_X1M_A12TR sub_1478_u13 ( .A(sub_1478_n9), .B(rfsr1h[0]), .Y(sub_1478_n1)
         );
  XNOR2_X1M_A12TR sub_1478_u12 ( .A(rfsr1h[1]), .B(sub_1478_n1), .Y(
        wfsrdec1[9]) );
  XNOR2_X1M_A12TR sub_1478_u11 ( .A(rfsr1h[3]), .B(sub_1478_n10), .Y(
        wfsrdec1[11]) );
  XNOR2_X1M_A12TR sub_1478_u10 ( .A(rfsr1h[2]), .B(sub_1478_n2), .Y(
        wfsrdec1[10]) );
  XNOR2_X1M_A12TR sub_1478_u9 ( .A(rfsr1h[0]), .B(sub_1478_n9), .Y(wfsrdec1[8]) );
  INV_X1M_A12TR sub_1478_u8 ( .A(rfsr1l[0]), .Y(wfsrdec1[0]) );
  XNOR2_X1M_A12TR sub_1478_u7 ( .A(rfsr1l[1]), .B(rfsr1l[0]), .Y(wfsrdec1[1])
         );
  XNOR2_X1M_A12TR sub_1478_u6 ( .A(rfsr1l[2]), .B(sub_1478_n6), .Y(wfsrdec1[2]) );
  XNOR2_X1M_A12TR sub_1478_u5 ( .A(rfsr1l[3]), .B(sub_1478_n5), .Y(wfsrdec1[3]) );
  XNOR2_X1M_A12TR sub_1478_u4 ( .A(rfsr1l[4]), .B(sub_1478_n4), .Y(wfsrdec1[4]) );
  XNOR2_X1M_A12TR sub_1478_u3 ( .A(rfsr1l[5]), .B(sub_1478_n3), .Y(wfsrdec1[5]) );
  XNOR2_X1M_A12TR sub_1478_u2 ( .A(rfsr1l[6]), .B(sub_1478_n8), .Y(wfsrdec1[6]) );
  XNOR2_X1M_A12TR sub_1478_u1 ( .A(rfsr1l[7]), .B(sub_1478_n7), .Y(wfsrdec1[7]) );
  XOR2_X0P5M_A12TR add_1550_u2 ( .A(add_1550_carry[19]), .B(wtblat[19]), .Y(
        wtblinc[19]) );
  INV_X1M_A12TR add_1550_u1 ( .A(wtblat[0]), .Y(wtblinc[0]) );
  ADDH_X1M_A12TR add_1550_u1_1_1 ( .A(wtblat[1]), .B(wtblat[0]), .CO(
        add_1550_carry[2]), .S(wtblinc[1]) );
  ADDH_X1M_A12TR add_1550_u1_1_4 ( .A(wtblat[4]), .B(add_1550_carry[4]), .CO(
        add_1550_carry[5]), .S(wtblinc[4]) );
  ADDH_X1M_A12TR add_1550_u1_1_2 ( .A(wtblat[2]), .B(add_1550_carry[2]), .CO(
        add_1550_carry[3]), .S(wtblinc[2]) );
  ADDH_X1M_A12TR add_1550_u1_1_3 ( .A(wtblat[3]), .B(add_1550_carry[3]), .CO(
        add_1550_carry[4]), .S(wtblinc[3]) );
  ADDH_X1M_A12TR add_1550_u1_1_5 ( .A(wtblat[5]), .B(add_1550_carry[5]), .CO(
        add_1550_carry[6]), .S(wtblinc[5]) );
  ADDH_X1M_A12TR add_1550_u1_1_6 ( .A(wtblat[6]), .B(add_1550_carry[6]), .CO(
        add_1550_carry[7]), .S(wtblinc[6]) );
  ADDH_X1M_A12TR add_1550_u1_1_7 ( .A(wtblat[7]), .B(add_1550_carry[7]), .CO(
        add_1550_carry[8]), .S(wtblinc[7]) );
  ADDH_X1M_A12TR add_1550_u1_1_9 ( .A(wtblat[9]), .B(add_1550_carry[9]), .CO(
        add_1550_carry[10]), .S(wtblinc[9]) );
  ADDH_X1M_A12TR add_1550_u1_1_10 ( .A(wtblat[10]), .B(add_1550_carry[10]), 
        .CO(add_1550_carry[11]), .S(wtblinc[10]) );
  ADDH_X1M_A12TR add_1550_u1_1_11 ( .A(wtblat[11]), .B(add_1550_carry[11]), 
        .CO(add_1550_carry[12]), .S(wtblinc[11]) );
  ADDH_X1M_A12TR add_1550_u1_1_12 ( .A(wtblat[12]), .B(add_1550_carry[12]), 
        .CO(add_1550_carry[13]), .S(wtblinc[12]) );
  ADDH_X1M_A12TR add_1550_u1_1_13 ( .A(wtblat[13]), .B(add_1550_carry[13]), 
        .CO(add_1550_carry[14]), .S(wtblinc[13]) );
  ADDH_X1M_A12TR add_1550_u1_1_14 ( .A(wtblat[14]), .B(add_1550_carry[14]), 
        .CO(add_1550_carry[15]), .S(wtblinc[14]) );
  ADDH_X1M_A12TR add_1550_u1_1_15 ( .A(wtblat[15]), .B(add_1550_carry[15]), 
        .CO(add_1550_carry[16]), .S(wtblinc[15]) );
  ADDH_X1M_A12TR add_1550_u1_1_16 ( .A(wtblat[16]), .B(add_1550_carry[16]), 
        .CO(add_1550_carry[17]), .S(wtblinc[16]) );
  ADDH_X1M_A12TR add_1550_u1_1_8 ( .A(wtblat[8]), .B(add_1550_carry[8]), .CO(
        add_1550_carry[9]), .S(wtblinc[8]) );
  ADDH_X1M_A12TR add_1550_u1_1_17 ( .A(wtblat[17]), .B(add_1550_carry[17]), 
        .CO(add_1550_carry[18]), .S(wtblinc[17]) );
  ADDH_X1M_A12TR add_1550_u1_1_18 ( .A(wtblat[18]), .B(add_1550_carry[18]), 
        .CO(add_1550_carry[19]), .S(wtblinc[18]) );
  AND2_X1M_A12TR add_1151_u9 ( .A(rfsr1h[1]), .B(add_1151_n2), .Y(add_1151_n3)
         );
  AND2_X1M_A12TR add_1151_u8 ( .A(rfsr1h[0]), .B(add_1151_carry_8_), .Y(
        add_1151_n2) );
  AND2_X1M_A12TR add_1151_u7 ( .A(rwreg[0]), .B(rfsr1l[0]), .Y(add_1151_n1) );
  XOR2_X1M_A12TR add_1151_u6 ( .A(rfsr1h[1]), .B(add_1151_n2), .Y(
        wfsrplusw1[9]) );
  XOR2_X1M_A12TR add_1151_u5 ( .A(rfsr1h[2]), .B(add_1151_n3), .Y(
        wfsrplusw1[10]) );
  NAND2_X1M_A12TR add_1151_u4 ( .A(rfsr1h[2]), .B(add_1151_n3), .Y(add_1151_n4) );
  XNOR2_X1M_A12TR add_1151_u3 ( .A(rfsr1h[3]), .B(add_1151_n4), .Y(
        wfsrplusw1[11]) );
  XOR2_X1M_A12TR add_1151_u2 ( .A(rwreg[0]), .B(rfsr1l[0]), .Y(wfsrplusw1[0])
         );
  XOR2_X1M_A12TR add_1151_u1 ( .A(rfsr1h[0]), .B(add_1151_carry_8_), .Y(
        wfsrplusw1[8]) );
  ADDF_X1M_A12TR add_1151_u1_1 ( .A(rfsr1l[1]), .B(rwreg[1]), .CI(add_1151_n1), 
        .CO(add_1151_carry_2_), .S(wfsrplusw1[1]) );
  ADDF_X1M_A12TR add_1151_u1_2 ( .A(rfsr1l[2]), .B(rwreg[2]), .CI(
        add_1151_carry_2_), .CO(add_1151_carry_3_), .S(wfsrplusw1[2]) );
  ADDF_X1M_A12TR add_1151_u1_3 ( .A(rfsr1l[3]), .B(rwreg[3]), .CI(
        add_1151_carry_3_), .CO(add_1151_carry_4_), .S(wfsrplusw1[3]) );
  ADDF_X1M_A12TR add_1151_u1_4 ( .A(rfsr1l[4]), .B(rwreg[4]), .CI(
        add_1151_carry_4_), .CO(add_1151_carry_5_), .S(wfsrplusw1[4]) );
  ADDF_X1M_A12TR add_1151_u1_5 ( .A(rfsr1l[5]), .B(rwreg[5]), .CI(
        add_1151_carry_5_), .CO(add_1151_carry_6_), .S(wfsrplusw1[5]) );
  ADDF_X1M_A12TR add_1151_u1_6 ( .A(rfsr1l[6]), .B(rwreg[6]), .CI(
        add_1151_carry_6_), .CO(add_1151_carry_7_), .S(wfsrplusw1[6]) );
  ADDF_X1M_A12TR add_1151_u1_7 ( .A(rfsr1l[7]), .B(rwreg[7]), .CI(
        add_1151_carry_7_), .CO(add_1151_carry_8_), .S(wfsrplusw1[7]) );
  AND2_X1M_A12TR add_1150_u9 ( .A(rfsr0h[1]), .B(add_1150_n2), .Y(add_1150_n3)
         );
  AND2_X1M_A12TR add_1150_u8 ( .A(rfsr0h[0]), .B(add_1150_carry_8_), .Y(
        add_1150_n2) );
  AND2_X1M_A12TR add_1150_u7 ( .A(rwreg[0]), .B(rfsr0l[0]), .Y(add_1150_n1) );
  XOR2_X1M_A12TR add_1150_u6 ( .A(rfsr0h[1]), .B(add_1150_n2), .Y(
        wfsrplusw0[9]) );
  XOR2_X1M_A12TR add_1150_u5 ( .A(rfsr0h[2]), .B(add_1150_n3), .Y(
        wfsrplusw0[10]) );
  NAND2_X1M_A12TR add_1150_u4 ( .A(rfsr0h[2]), .B(add_1150_n3), .Y(add_1150_n4) );
  XNOR2_X1M_A12TR add_1150_u3 ( .A(rfsr0h[3]), .B(add_1150_n4), .Y(
        wfsrplusw0[11]) );
  XOR2_X1M_A12TR add_1150_u2 ( .A(rwreg[0]), .B(rfsr0l[0]), .Y(wfsrplusw0[0])
         );
  XOR2_X1M_A12TR add_1150_u1 ( .A(rfsr0h[0]), .B(add_1150_carry_8_), .Y(
        wfsrplusw0[8]) );
  ADDF_X1M_A12TR add_1150_u1_1 ( .A(rfsr0l[1]), .B(rwreg[1]), .CI(add_1150_n1), 
        .CO(add_1150_carry_2_), .S(wfsrplusw0[1]) );
  ADDF_X1M_A12TR add_1150_u1_2 ( .A(rfsr0l[2]), .B(rwreg[2]), .CI(
        add_1150_carry_2_), .CO(add_1150_carry_3_), .S(wfsrplusw0[2]) );
  ADDF_X1M_A12TR add_1150_u1_3 ( .A(rfsr0l[3]), .B(rwreg[3]), .CI(
        add_1150_carry_3_), .CO(add_1150_carry_4_), .S(wfsrplusw0[3]) );
  ADDF_X1M_A12TR add_1150_u1_4 ( .A(rfsr0l[4]), .B(rwreg[4]), .CI(
        add_1150_carry_4_), .CO(add_1150_carry_5_), .S(wfsrplusw0[4]) );
  ADDF_X1M_A12TR add_1150_u1_5 ( .A(rfsr0l[5]), .B(rwreg[5]), .CI(
        add_1150_carry_5_), .CO(add_1150_carry_6_), .S(wfsrplusw0[5]) );
  ADDF_X1M_A12TR add_1150_u1_6 ( .A(rfsr0l[6]), .B(rwreg[6]), .CI(
        add_1150_carry_6_), .CO(add_1150_carry_7_), .S(wfsrplusw0[6]) );
  ADDF_X1M_A12TR add_1150_u1_7 ( .A(rfsr0l[7]), .B(rwreg[7]), .CI(
        add_1150_carry_7_), .CO(add_1150_carry_8_), .S(wfsrplusw0[7]) );
  XOR2_X0P5M_A12TR add_1149_u2 ( .A(add_1149_carry[11]), .B(rfsr2h[3]), .Y(
        wfsrinc2[11]) );
  INV_X1M_A12TR add_1149_u1 ( .A(rfsr2l[0]), .Y(wfsrinc2[0]) );
  ADDH_X1M_A12TR add_1149_u1_1_1 ( .A(rfsr2l[1]), .B(rfsr2l[0]), .CO(
        add_1149_carry[2]), .S(wfsrinc2[1]) );
  ADDH_X1M_A12TR add_1149_u1_1_9 ( .A(rfsr2h[1]), .B(add_1149_carry[9]), .CO(
        add_1149_carry[10]), .S(wfsrinc2[9]) );
  ADDH_X1M_A12TR add_1149_u1_1_8 ( .A(rfsr2h[0]), .B(add_1149_carry[8]), .CO(
        add_1149_carry[9]), .S(wfsrinc2[8]) );
  ADDH_X1M_A12TR add_1149_u1_1_6 ( .A(rfsr2l[6]), .B(add_1149_carry[6]), .CO(
        add_1149_carry[7]), .S(wfsrinc2[6]) );
  ADDH_X1M_A12TR add_1149_u1_1_7 ( .A(rfsr2l[7]), .B(add_1149_carry[7]), .CO(
        add_1149_carry[8]), .S(wfsrinc2[7]) );
  ADDH_X1M_A12TR add_1149_u1_1_2 ( .A(rfsr2l[2]), .B(add_1149_carry[2]), .CO(
        add_1149_carry[3]), .S(wfsrinc2[2]) );
  ADDH_X1M_A12TR add_1149_u1_1_3 ( .A(rfsr2l[3]), .B(add_1149_carry[3]), .CO(
        add_1149_carry[4]), .S(wfsrinc2[3]) );
  ADDH_X1M_A12TR add_1149_u1_1_5 ( .A(rfsr2l[5]), .B(add_1149_carry[5]), .CO(
        add_1149_carry[6]), .S(wfsrinc2[5]) );
  ADDH_X1M_A12TR add_1149_u1_1_4 ( .A(rfsr2l[4]), .B(add_1149_carry[4]), .CO(
        add_1149_carry[5]), .S(wfsrinc2[4]) );
  ADDH_X1M_A12TR add_1149_u1_1_10 ( .A(rfsr2h[2]), .B(add_1149_carry[10]), 
        .CO(add_1149_carry[11]), .S(wfsrinc2[10]) );
  XOR2_X0P5M_A12TR add_1148_u2 ( .A(add_1148_carry[11]), .B(rfsr1h[3]), .Y(
        wfsrinc1[11]) );
  INV_X1M_A12TR add_1148_u1 ( .A(rfsr1l[0]), .Y(wfsrinc1[0]) );
  ADDH_X1M_A12TR add_1148_u1_1_1 ( .A(rfsr1l[1]), .B(rfsr1l[0]), .CO(
        add_1148_carry[2]), .S(wfsrinc1[1]) );
  ADDH_X1M_A12TR add_1148_u1_1_8 ( .A(rfsr1h[0]), .B(add_1148_carry[8]), .CO(
        add_1148_carry[9]), .S(wfsrinc1[8]) );
  ADDH_X1M_A12TR add_1148_u1_1_9 ( .A(rfsr1h[1]), .B(add_1148_carry[9]), .CO(
        add_1148_carry[10]), .S(wfsrinc1[9]) );
  ADDH_X1M_A12TR add_1148_u1_1_2 ( .A(rfsr1l[2]), .B(add_1148_carry[2]), .CO(
        add_1148_carry[3]), .S(wfsrinc1[2]) );
  ADDH_X1M_A12TR add_1148_u1_1_3 ( .A(rfsr1l[3]), .B(add_1148_carry[3]), .CO(
        add_1148_carry[4]), .S(wfsrinc1[3]) );
  ADDH_X1M_A12TR add_1148_u1_1_4 ( .A(rfsr1l[4]), .B(add_1148_carry[4]), .CO(
        add_1148_carry[5]), .S(wfsrinc1[4]) );
  ADDH_X1M_A12TR add_1148_u1_1_6 ( .A(rfsr1l[6]), .B(add_1148_carry[6]), .CO(
        add_1148_carry[7]), .S(wfsrinc1[6]) );
  ADDH_X1M_A12TR add_1148_u1_1_7 ( .A(rfsr1l[7]), .B(add_1148_carry[7]), .CO(
        add_1148_carry[8]), .S(wfsrinc1[7]) );
  ADDH_X1M_A12TR add_1148_u1_1_5 ( .A(rfsr1l[5]), .B(add_1148_carry[5]), .CO(
        add_1148_carry[6]), .S(wfsrinc1[5]) );
  ADDH_X1M_A12TR add_1148_u1_1_10 ( .A(rfsr1h[2]), .B(add_1148_carry[10]), 
        .CO(add_1148_carry[11]), .S(wfsrinc1[10]) );
  XOR2_X0P5M_A12TR add_1147_u2 ( .A(add_1147_carry[11]), .B(rfsr0h[3]), .Y(
        wfsrinc0[11]) );
  INV_X1M_A12TR add_1147_u1 ( .A(rfsr0l[0]), .Y(wfsrinc0[0]) );
  ADDH_X1M_A12TR add_1147_u1_1_1 ( .A(rfsr0l[1]), .B(rfsr0l[0]), .CO(
        add_1147_carry[2]), .S(wfsrinc0[1]) );
  ADDH_X1M_A12TR add_1147_u1_1_9 ( .A(rfsr0h[1]), .B(add_1147_carry[9]), .CO(
        add_1147_carry[10]), .S(wfsrinc0[9]) );
  ADDH_X1M_A12TR add_1147_u1_1_8 ( .A(rfsr0h[0]), .B(add_1147_carry[8]), .CO(
        add_1147_carry[9]), .S(wfsrinc0[8]) );
  ADDH_X1M_A12TR add_1147_u1_1_6 ( .A(rfsr0l[6]), .B(add_1147_carry[6]), .CO(
        add_1147_carry[7]), .S(wfsrinc0[6]) );
  ADDH_X1M_A12TR add_1147_u1_1_7 ( .A(rfsr0l[7]), .B(add_1147_carry[7]), .CO(
        add_1147_carry[8]), .S(wfsrinc0[7]) );
  ADDH_X1M_A12TR add_1147_u1_1_5 ( .A(rfsr0l[5]), .B(add_1147_carry[5]), .CO(
        add_1147_carry[6]), .S(wfsrinc0[5]) );
  ADDH_X1M_A12TR add_1147_u1_1_2 ( .A(rfsr0l[2]), .B(add_1147_carry[2]), .CO(
        add_1147_carry[3]), .S(wfsrinc0[2]) );
  ADDH_X1M_A12TR add_1147_u1_1_3 ( .A(rfsr0l[3]), .B(add_1147_carry[3]), .CO(
        add_1147_carry[4]), .S(wfsrinc0[3]) );
  ADDH_X1M_A12TR add_1147_u1_1_4 ( .A(rfsr0l[4]), .B(add_1147_carry[4]), .CO(
        add_1147_carry[5]), .S(wfsrinc0[4]) );
  ADDH_X1M_A12TR add_1147_u1_1_10 ( .A(rfsr0h[2]), .B(add_1147_carry[10]), 
        .CO(add_1147_carry[11]), .S(wfsrinc0[10]) );
  INV_X1M_A12TR sub_1006_u11 ( .A(rsrc[0]), .Y(sub_1006_n3) );
  INV_X1M_A12TR sub_1006_u10 ( .A(rsrc[6]), .Y(sub_1006_n9) );
  INV_X1M_A12TR sub_1006_u9 ( .A(rsrc[2]), .Y(sub_1006_n7) );
  INV_X1M_A12TR sub_1006_u8 ( .A(rsrc[3]), .Y(sub_1006_n8) );
  INV_X1M_A12TR sub_1006_u7 ( .A(rsrc[5]), .Y(sub_1006_n10) );
  OR2_X1M_A12TR sub_1006_u6 ( .A(wneg[0]), .B(sub_1006_n3), .Y(sub_1006_n1) );
  INV_X1M_A12TR sub_1006_u5 ( .A(rsrc[4]), .Y(sub_1006_n6) );
  INV_X1M_A12TR sub_1006_u4 ( .A(rsrc[7]), .Y(sub_1006_n4) );
  XNOR2_X1M_A12TR sub_1006_u3 ( .A(sub_1006_n3), .B(wneg[0]), .Y(wsub[0]) );
  INV_X1M_A12TR sub_1006_u2 ( .A(sub_1006_carry[8]), .Y(wsub[8]) );
  INV_X1M_A12TR sub_1006_u1 ( .A(rsrc[1]), .Y(sub_1006_n5) );
  ADDF_X1M_A12TR sub_1006_u2_1 ( .A(rtgt[1]), .B(sub_1006_n5), .CI(sub_1006_n1), .CO(sub_1006_carry[2]), .S(wsub[1]) );
  ADDF_X1M_A12TR sub_1006_u2_2 ( .A(rtgt[2]), .B(sub_1006_n7), .CI(
        sub_1006_carry[2]), .CO(sub_1006_carry[3]), .S(wsub[2]) );
  ADDF_X1M_A12TR sub_1006_u2_3 ( .A(rtgt[3]), .B(sub_1006_n8), .CI(
        sub_1006_carry[3]), .CO(sub_1006_carry[4]), .S(wsub[3]) );
  ADDF_X1M_A12TR sub_1006_u2_4 ( .A(rtgt[4]), .B(sub_1006_n6), .CI(
        sub_1006_carry[4]), .CO(sub_1006_carry[5]), .S(wsub[4]) );
  ADDF_X1M_A12TR sub_1006_u2_5 ( .A(rtgt[5]), .B(sub_1006_n10), .CI(
        sub_1006_carry[5]), .CO(sub_1006_carry[6]), .S(wsub[5]) );
  ADDF_X1M_A12TR sub_1006_u2_6 ( .A(rtgt[6]), .B(sub_1006_n9), .CI(
        sub_1006_carry[6]), .CO(sub_1006_carry[7]), .S(wsub[6]) );
  ADDF_X1M_A12TR sub_1006_u2_7 ( .A(rtgt[7]), .B(sub_1006_n4), .CI(
        sub_1006_carry[7]), .CO(sub_1006_carry[8]), .S(wsub[7]) );
  AND2_X1M_A12TR add_1004_u2 ( .A(wneg[0]), .B(rsrc[0]), .Y(add_1004_n1) );
  XOR2_X1M_A12TR add_1004_u1 ( .A(wneg[0]), .B(rsrc[0]), .Y(wadd[0]) );
  ADDF_X1M_A12TR add_1004_u1_1 ( .A(rsrc[1]), .B(rtgt[1]), .CI(add_1004_n1), 
        .CO(add_1004_carry[2]), .S(wadd[1]) );
  ADDF_X1M_A12TR add_1004_u1_2 ( .A(rsrc[2]), .B(rtgt[2]), .CI(
        add_1004_carry[2]), .CO(add_1004_carry[3]), .S(wadd[2]) );
  ADDF_X1M_A12TR add_1004_u1_3 ( .A(rsrc[3]), .B(rtgt[3]), .CI(
        add_1004_carry[3]), .CO(add_1004_carry[4]), .S(wadd[3]) );
  ADDF_X1M_A12TR add_1004_u1_4 ( .A(rsrc[4]), .B(rtgt[4]), .CI(
        add_1004_carry[4]), .CO(add_1004_carry[5]), .S(wadd[4]) );
  ADDF_X1M_A12TR add_1004_u1_5 ( .A(rsrc[5]), .B(rtgt[5]), .CI(
        add_1004_carry[5]), .CO(add_1004_carry[6]), .S(wadd[5]) );
  ADDF_X1M_A12TR add_1004_u1_6 ( .A(rsrc[6]), .B(rtgt[6]), .CI(
        add_1004_carry[6]), .CO(add_1004_carry[7]), .S(wadd[6]) );
  ADDF_X1M_A12TR add_1004_u1_7 ( .A(rsrc[7]), .B(rtgt[7]), .CI(
        add_1004_carry[7]), .CO(wadd[8]), .S(wadd[7]) );
  AND2_X1M_A12TR add_436_u2 ( .A(rireg[0]), .B(iwb_adr_o[1]), .Y(add_436_n1)
         );
  XOR2_X1M_A12TR add_436_u1 ( .A(rireg[0]), .B(iwb_adr_o[1]), .Y(n386) );
  ADDF_X1M_A12TR add_436_u1_1 ( .A(iwb_adr_o[2]), .B(rireg[1]), .CI(add_436_n1), .CO(add_436_carry[2]), .S(n387) );
  ADDF_X1M_A12TR add_436_u1_2 ( .A(iwb_adr_o[3]), .B(rireg[2]), .CI(
        add_436_carry[2]), .CO(add_436_carry[3]), .S(n388) );
  ADDF_X1M_A12TR add_436_u1_3 ( .A(iwb_adr_o[4]), .B(rireg[3]), .CI(
        add_436_carry[3]), .CO(add_436_carry[4]), .S(n389) );
  ADDF_X1M_A12TR add_436_u1_4 ( .A(iwb_adr_o[5]), .B(rireg[4]), .CI(
        add_436_carry[4]), .CO(add_436_carry[5]), .S(n390) );
  ADDF_X1M_A12TR add_436_u1_5 ( .A(iwb_adr_o[6]), .B(rireg[5]), .CI(
        add_436_carry[5]), .CO(add_436_carry[6]), .S(n391) );
  ADDF_X1M_A12TR add_436_u1_6 ( .A(iwb_adr_o[7]), .B(rireg[6]), .CI(
        add_436_carry[6]), .CO(add_436_carry[7]), .S(n392) );
  ADDF_X1M_A12TR add_436_u1_7 ( .A(iwb_adr_o[8]), .B(rireg[7]), .CI(
        add_436_carry[7]), .CO(add_436_carry[8]), .S(n393) );
  ADDF_X1M_A12TR add_436_u1_8 ( .A(iwb_adr_o[9]), .B(rireg[8]), .CI(
        add_436_carry[8]), .CO(add_436_carry[9]), .S(n394) );
  ADDF_X1M_A12TR add_436_u1_9 ( .A(iwb_adr_o[10]), .B(rireg[9]), .CI(
        add_436_carry[9]), .CO(add_436_carry[10]), .S(n395) );
  ADDF_X1M_A12TR add_436_u1_10 ( .A(iwb_adr_o[11]), .B(rireg[10]), .CI(
        add_436_carry[10]), .CO(add_436_carry[11]), .S(n396) );
  ADDF_X1M_A12TR add_436_u1_11 ( .A(iwb_adr_o[12]), .B(rireg[10]), .CI(
        add_436_carry[11]), .CO(add_436_carry[12]), .S(n397) );
  ADDF_X1M_A12TR add_436_u1_12 ( .A(iwb_adr_o[13]), .B(rireg[10]), .CI(
        add_436_carry[12]), .CO(add_436_carry[13]), .S(n398) );
  ADDF_X1M_A12TR add_436_u1_13 ( .A(iwb_adr_o[14]), .B(rireg[10]), .CI(
        add_436_carry[13]), .CO(add_436_carry[14]), .S(n399) );
  ADDF_X1M_A12TR add_436_u1_14 ( .A(iwb_adr_o[15]), .B(rireg[10]), .CI(
        add_436_carry[14]), .CO(add_436_carry[15]), .S(n400) );
  ADDF_X1M_A12TR add_436_u1_15 ( .A(iwb_adr_o[16]), .B(rireg[10]), .CI(
        add_436_carry[15]), .CO(add_436_carry[16]), .S(n401) );
  ADDF_X1M_A12TR add_436_u1_16 ( .A(iwb_adr_o[17]), .B(rireg[10]), .CI(
        add_436_carry[16]), .CO(add_436_carry[17]), .S(n402) );
  ADDF_X1M_A12TR add_436_u1_17 ( .A(iwb_adr_o[18]), .B(rireg[10]), .CI(
        add_436_carry[17]), .CO(add_436_carry[18]), .S(n403) );
  ADDF_X1M_A12TR add_436_u1_18 ( .A(iwb_adr_o[19]), .B(rireg[10]), .CI(
        add_436_carry[18]), .CO(), .S(n404) );
  XOR2_X0P5M_A12TR add_433_u2 ( .A(add_433_carry[18]), .B(iwb_adr_o[19]), .Y(
        wpcinc[18]) );
  INV_X1M_A12TR add_433_u1 ( .A(iwb_adr_o[1]), .Y(wpcinc[0]) );
  ADDH_X1M_A12TR add_433_u1_1_1 ( .A(iwb_adr_o[2]), .B(iwb_adr_o[1]), .CO(
        add_433_carry[2]), .S(wpcinc[1]) );
  ADDH_X1M_A12TR add_433_u1_1_2 ( .A(iwb_adr_o[3]), .B(add_433_carry[2]), .CO(
        add_433_carry[3]), .S(wpcinc[2]) );
  ADDH_X1M_A12TR add_433_u1_1_3 ( .A(iwb_adr_o[4]), .B(add_433_carry[3]), .CO(
        add_433_carry[4]), .S(wpcinc[3]) );
  ADDH_X1M_A12TR add_433_u1_1_5 ( .A(iwb_adr_o[6]), .B(add_433_carry[5]), .CO(
        add_433_carry[6]), .S(wpcinc[5]) );
  ADDH_X1M_A12TR add_433_u1_1_6 ( .A(iwb_adr_o[7]), .B(add_433_carry[6]), .CO(
        add_433_carry[7]), .S(wpcinc[6]) );
  ADDH_X1M_A12TR add_433_u1_1_7 ( .A(iwb_adr_o[8]), .B(add_433_carry[7]), .CO(
        add_433_carry[8]), .S(wpcinc[7]) );
  ADDH_X1M_A12TR add_433_u1_1_8 ( .A(iwb_adr_o[9]), .B(add_433_carry[8]), .CO(
        add_433_carry[9]), .S(wpcinc[8]) );
  ADDH_X1M_A12TR add_433_u1_1_9 ( .A(iwb_adr_o[10]), .B(add_433_carry[9]), 
        .CO(add_433_carry[10]), .S(wpcinc[9]) );
  ADDH_X1M_A12TR add_433_u1_1_10 ( .A(iwb_adr_o[11]), .B(add_433_carry[10]), 
        .CO(add_433_carry[11]), .S(wpcinc[10]) );
  ADDH_X1M_A12TR add_433_u1_1_11 ( .A(iwb_adr_o[12]), .B(add_433_carry[11]), 
        .CO(add_433_carry[12]), .S(wpcinc[11]) );
  ADDH_X1M_A12TR add_433_u1_1_12 ( .A(iwb_adr_o[13]), .B(add_433_carry[12]), 
        .CO(add_433_carry[13]), .S(wpcinc[12]) );
  ADDH_X1M_A12TR add_433_u1_1_13 ( .A(iwb_adr_o[14]), .B(add_433_carry[13]), 
        .CO(add_433_carry[14]), .S(wpcinc[13]) );
  ADDH_X1M_A12TR add_433_u1_1_14 ( .A(iwb_adr_o[15]), .B(add_433_carry[14]), 
        .CO(add_433_carry[15]), .S(wpcinc[14]) );
  ADDH_X1M_A12TR add_433_u1_1_15 ( .A(iwb_adr_o[16]), .B(add_433_carry[15]), 
        .CO(add_433_carry[16]), .S(wpcinc[15]) );
  ADDH_X1M_A12TR add_433_u1_1_16 ( .A(iwb_adr_o[17]), .B(add_433_carry[16]), 
        .CO(add_433_carry[17]), .S(wpcinc[16]) );
  ADDH_X1M_A12TR add_433_u1_1_4 ( .A(iwb_adr_o[5]), .B(add_433_carry[4]), .CO(
        add_433_carry[5]), .S(wpcinc[4]) );
  ADDH_X1M_A12TR add_433_u1_1_17 ( .A(iwb_adr_o[18]), .B(add_433_carry[17]), 
        .CO(add_433_carry[18]), .S(wpcinc[17]) );
  XOR2_X0P5M_A12TR add_276_u2 ( .A(add_276_carry[16]), .B(rwdt[16]), .Y(n240)
         );
  INV_X1M_A12TR add_276_u1 ( .A(rwdt[0]), .Y(n224) );
  ADDH_X1M_A12TR add_276_u1_1_1 ( .A(rwdt[1]), .B(rwdt[0]), .CO(
        add_276_carry[2]), .S(n225) );
  ADDH_X1M_A12TR add_276_u1_1_2 ( .A(rwdt[2]), .B(add_276_carry[2]), .CO(
        add_276_carry[3]), .S(n226) );
  ADDH_X1M_A12TR add_276_u1_1_3 ( .A(rwdt[3]), .B(add_276_carry[3]), .CO(
        add_276_carry[4]), .S(n227) );
  ADDH_X1M_A12TR add_276_u1_1_4 ( .A(rwdt[4]), .B(add_276_carry[4]), .CO(
        add_276_carry[5]), .S(n228) );
  ADDH_X1M_A12TR add_276_u1_1_5 ( .A(rwdt[5]), .B(add_276_carry[5]), .CO(
        add_276_carry[6]), .S(n229) );
  ADDH_X1M_A12TR add_276_u1_1_6 ( .A(rwdt[6]), .B(add_276_carry[6]), .CO(
        add_276_carry[7]), .S(n230) );
  ADDH_X1M_A12TR add_276_u1_1_7 ( .A(rwdt[7]), .B(add_276_carry[7]), .CO(
        add_276_carry[8]), .S(n231) );
  ADDH_X1M_A12TR add_276_u1_1_8 ( .A(rwdt[8]), .B(add_276_carry[8]), .CO(
        add_276_carry[9]), .S(n232) );
  ADDH_X1M_A12TR add_276_u1_1_9 ( .A(rwdt[9]), .B(add_276_carry[9]), .CO(
        add_276_carry[10]), .S(n233) );
  ADDH_X1M_A12TR add_276_u1_1_10 ( .A(rwdt[10]), .B(add_276_carry[10]), .CO(
        add_276_carry[11]), .S(n234) );
  ADDH_X1M_A12TR add_276_u1_1_11 ( .A(rwdt[11]), .B(add_276_carry[11]), .CO(
        add_276_carry[12]), .S(n235) );
  ADDH_X1M_A12TR add_276_u1_1_12 ( .A(rwdt[12]), .B(add_276_carry[12]), .CO(
        add_276_carry[13]), .S(n236) );
  ADDH_X1M_A12TR add_276_u1_1_13 ( .A(rwdt[13]), .B(add_276_carry[13]), .CO(
        add_276_carry[14]), .S(n237) );
  ADDH_X1M_A12TR add_276_u1_1_14 ( .A(rwdt[14]), .B(add_276_carry[14]), .CO(
        add_276_carry[15]), .S(n238) );
  ADDH_X1M_A12TR add_276_u1_1_15 ( .A(rwdt[15]), .B(add_276_carry[15]), .CO(
        add_276_carry[16]), .S(n239) );
  OR2_X1M_A12TR sub_1477_u22 ( .A(sub_1477_n1), .B(rfsr0h[2]), .Y(sub_1477_n10) );
  OR2_X1M_A12TR sub_1477_u21 ( .A(sub_1477_n6), .B(rfsr0l[4]), .Y(sub_1477_n9)
         );
  OR2_X1M_A12TR sub_1477_u20 ( .A(rfsr0l[0]), .B(rfsr0l[1]), .Y(sub_1477_n8)
         );
  OR2_X1M_A12TR sub_1477_u19 ( .A(sub_1477_n8), .B(rfsr0l[2]), .Y(sub_1477_n7)
         );
  OR2_X1M_A12TR sub_1477_u18 ( .A(sub_1477_n7), .B(rfsr0l[3]), .Y(sub_1477_n6)
         );
  OR2_X1M_A12TR sub_1477_u17 ( .A(sub_1477_n9), .B(rfsr0l[5]), .Y(sub_1477_n5)
         );
  OR2_X1M_A12TR sub_1477_u16 ( .A(sub_1477_n5), .B(rfsr0l[6]), .Y(sub_1477_n4)
         );
  OR2_X1M_A12TR sub_1477_u15 ( .A(sub_1477_n4), .B(rfsr0l[7]), .Y(sub_1477_n3)
         );
  OR2_X1M_A12TR sub_1477_u14 ( .A(sub_1477_n3), .B(rfsr0h[0]), .Y(sub_1477_n2)
         );
  OR2_X1M_A12TR sub_1477_u13 ( .A(sub_1477_n2), .B(rfsr0h[1]), .Y(sub_1477_n1)
         );
  XNOR2_X1M_A12TR sub_1477_u12 ( .A(rfsr0l[5]), .B(sub_1477_n9), .Y(
        wfsrdec0[5]) );
  INV_X1M_A12TR sub_1477_u11 ( .A(rfsr0l[0]), .Y(wfsrdec0[0]) );
  XNOR2_X1M_A12TR sub_1477_u10 ( .A(rfsr0l[1]), .B(rfsr0l[0]), .Y(wfsrdec0[1])
         );
  XNOR2_X1M_A12TR sub_1477_u9 ( .A(rfsr0l[2]), .B(sub_1477_n8), .Y(wfsrdec0[2]) );
  XNOR2_X1M_A12TR sub_1477_u8 ( .A(rfsr0l[3]), .B(sub_1477_n7), .Y(wfsrdec0[3]) );
  XNOR2_X1M_A12TR sub_1477_u7 ( .A(rfsr0l[4]), .B(sub_1477_n6), .Y(wfsrdec0[4]) );
  XNOR2_X1M_A12TR sub_1477_u6 ( .A(rfsr0l[6]), .B(sub_1477_n5), .Y(wfsrdec0[6]) );
  XNOR2_X1M_A12TR sub_1477_u5 ( .A(rfsr0l[7]), .B(sub_1477_n4), .Y(wfsrdec0[7]) );
  XNOR2_X1M_A12TR sub_1477_u4 ( .A(rfsr0h[0]), .B(sub_1477_n3), .Y(wfsrdec0[8]) );
  XNOR2_X1M_A12TR sub_1477_u3 ( .A(rfsr0h[3]), .B(sub_1477_n10), .Y(
        wfsrdec0[11]) );
  XNOR2_X1M_A12TR sub_1477_u2 ( .A(rfsr0h[1]), .B(sub_1477_n2), .Y(wfsrdec0[9]) );
  XNOR2_X1M_A12TR sub_1477_u1 ( .A(rfsr0h[2]), .B(sub_1477_n1), .Y(
        wfsrdec0[10]) );
  AND2_X1M_A12TR add_1152_u9 ( .A(rfsr2h[1]), .B(add_1152_n2), .Y(add_1152_n3)
         );
  AND2_X1M_A12TR add_1152_u8 ( .A(rfsr2h[0]), .B(add_1152_carry_8_), .Y(
        add_1152_n2) );
  AND2_X1M_A12TR add_1152_u7 ( .A(rwreg[0]), .B(rfsr2l[0]), .Y(add_1152_n1) );
  XOR2_X1M_A12TR add_1152_u6 ( .A(rfsr2h[1]), .B(add_1152_n2), .Y(
        wfsrplusw2[9]) );
  XOR2_X1M_A12TR add_1152_u5 ( .A(rfsr2h[2]), .B(add_1152_n3), .Y(
        wfsrplusw2[10]) );
  NAND2_X1M_A12TR add_1152_u4 ( .A(rfsr2h[2]), .B(add_1152_n3), .Y(add_1152_n4) );
  XNOR2_X1M_A12TR add_1152_u3 ( .A(rfsr2h[3]), .B(add_1152_n4), .Y(
        wfsrplusw2[11]) );
  XOR2_X1M_A12TR add_1152_u2 ( .A(rwreg[0]), .B(rfsr2l[0]), .Y(wfsrplusw2[0])
         );
  XOR2_X1M_A12TR add_1152_u1 ( .A(rfsr2h[0]), .B(add_1152_carry_8_), .Y(
        wfsrplusw2[8]) );
  ADDF_X1M_A12TR add_1152_u1_1 ( .A(rfsr2l[1]), .B(rwreg[1]), .CI(add_1152_n1), 
        .CO(add_1152_carry_2_), .S(wfsrplusw2[1]) );
  ADDF_X1M_A12TR add_1152_u1_2 ( .A(rfsr2l[2]), .B(rwreg[2]), .CI(
        add_1152_carry_2_), .CO(add_1152_carry_3_), .S(wfsrplusw2[2]) );
  ADDF_X1M_A12TR add_1152_u1_3 ( .A(rfsr2l[3]), .B(rwreg[3]), .CI(
        add_1152_carry_3_), .CO(add_1152_carry_4_), .S(wfsrplusw2[3]) );
  ADDF_X1M_A12TR add_1152_u1_4 ( .A(rfsr2l[4]), .B(rwreg[4]), .CI(
        add_1152_carry_4_), .CO(add_1152_carry_5_), .S(wfsrplusw2[4]) );
  ADDF_X1M_A12TR add_1152_u1_5 ( .A(rfsr2l[5]), .B(rwreg[5]), .CI(
        add_1152_carry_5_), .CO(add_1152_carry_6_), .S(wfsrplusw2[5]) );
  ADDF_X1M_A12TR add_1152_u1_6 ( .A(rfsr2l[6]), .B(rwreg[6]), .CI(
        add_1152_carry_6_), .CO(add_1152_carry_7_), .S(wfsrplusw2[6]) );
  ADDF_X1M_A12TR add_1152_u1_7 ( .A(rfsr2l[7]), .B(rwreg[7]), .CI(
        add_1152_carry_7_), .CO(add_1152_carry_8_), .S(wfsrplusw2[7]) );
  INV_X1M_A12TR mult_1536_u155 ( .A(rsrc[6]), .Y(mult_1536_n171) );
  INV_X1M_A12TR mult_1536_u154 ( .A(rsrc[5]), .Y(mult_1536_n172) );
  INV_X1M_A12TR mult_1536_u153 ( .A(rsrc[4]), .Y(mult_1536_n173) );
  INV_X1M_A12TR mult_1536_u152 ( .A(rsrc[3]), .Y(mult_1536_n174) );
  INV_X1M_A12TR mult_1536_u151 ( .A(rsrc[2]), .Y(mult_1536_n175) );
  INV_X1M_A12TR mult_1536_u150 ( .A(rsrc[1]), .Y(mult_1536_n176) );
  INV_X1M_A12TR mult_1536_u149 ( .A(rsrc[0]), .Y(mult_1536_n177) );
  INV_X1M_A12TR mult_1536_u148 ( .A(rsrc[7]), .Y(mult_1536_n170) );
  INV_X1M_A12TR mult_1536_u147 ( .A(rtgt[6]), .Y(mult_1536_n163) );
  INV_X1M_A12TR mult_1536_u146 ( .A(rtgt[5]), .Y(mult_1536_n164) );
  INV_X1M_A12TR mult_1536_u145 ( .A(rtgt[3]), .Y(mult_1536_n166) );
  INV_X1M_A12TR mult_1536_u144 ( .A(rtgt[2]), .Y(mult_1536_n167) );
  INV_X1M_A12TR mult_1536_u143 ( .A(rtgt[1]), .Y(mult_1536_n168) );
  INV_X1M_A12TR mult_1536_u142 ( .A(rtgt[4]), .Y(mult_1536_n165) );
  INV_X1M_A12TR mult_1536_u141 ( .A(rtgt[7]), .Y(mult_1536_n162) );
  INV_X1M_A12TR mult_1536_u140 ( .A(wneg[0]), .Y(mult_1536_n169) );
  NOR2_X1M_A12TR mult_1536_u121 ( .A(mult_1536_n169), .B(mult_1536_n177), .Y(
        n17820) );
  NOR2_X1M_A12TR mult_1536_u120 ( .A(mult_1536_n168), .B(mult_1536_n177), .Y(
        mult_1536_n161) );
  NOR2_X1M_A12TR mult_1536_u119 ( .A(mult_1536_n167), .B(mult_1536_n177), .Y(
        mult_1536_n160) );
  NOR2_X1M_A12TR mult_1536_u118 ( .A(mult_1536_n166), .B(mult_1536_n177), .Y(
        mult_1536_n159) );
  NOR2_X1M_A12TR mult_1536_u117 ( .A(mult_1536_n165), .B(mult_1536_n177), .Y(
        mult_1536_n158) );
  NOR2_X1M_A12TR mult_1536_u116 ( .A(mult_1536_n164), .B(mult_1536_n177), .Y(
        mult_1536_n157) );
  NOR2_X1M_A12TR mult_1536_u115 ( .A(mult_1536_n163), .B(mult_1536_n177), .Y(
        mult_1536_n156) );
  NOR2_X1M_A12TR mult_1536_u114 ( .A(mult_1536_n162), .B(mult_1536_n177), .Y(
        mult_1536_n155) );
  NOR2_X1M_A12TR mult_1536_u113 ( .A(mult_1536_n169), .B(mult_1536_n176), .Y(
        mult_1536_n154) );
  NOR2_X1M_A12TR mult_1536_u112 ( .A(mult_1536_n168), .B(mult_1536_n176), .Y(
        mult_1536_n153) );
  NOR2_X1M_A12TR mult_1536_u111 ( .A(mult_1536_n167), .B(mult_1536_n176), .Y(
        mult_1536_n152) );
  NOR2_X1M_A12TR mult_1536_u110 ( .A(mult_1536_n166), .B(mult_1536_n176), .Y(
        mult_1536_n151) );
  NOR2_X1M_A12TR mult_1536_u109 ( .A(mult_1536_n165), .B(mult_1536_n176), .Y(
        mult_1536_n150) );
  NOR2_X1M_A12TR mult_1536_u108 ( .A(mult_1536_n164), .B(mult_1536_n176), .Y(
        mult_1536_n149) );
  NOR2_X1M_A12TR mult_1536_u107 ( .A(mult_1536_n163), .B(mult_1536_n176), .Y(
        mult_1536_n148) );
  NOR2_X1M_A12TR mult_1536_u106 ( .A(mult_1536_n162), .B(mult_1536_n176), .Y(
        mult_1536_n147) );
  NOR2_X1M_A12TR mult_1536_u105 ( .A(mult_1536_n169), .B(mult_1536_n175), .Y(
        mult_1536_n146) );
  NOR2_X1M_A12TR mult_1536_u104 ( .A(mult_1536_n168), .B(mult_1536_n175), .Y(
        mult_1536_n145) );
  NOR2_X1M_A12TR mult_1536_u103 ( .A(mult_1536_n167), .B(mult_1536_n175), .Y(
        mult_1536_n144) );
  NOR2_X1M_A12TR mult_1536_u102 ( .A(mult_1536_n166), .B(mult_1536_n175), .Y(
        mult_1536_n143) );
  NOR2_X1M_A12TR mult_1536_u101 ( .A(mult_1536_n165), .B(mult_1536_n175), .Y(
        mult_1536_n142) );
  NOR2_X1M_A12TR mult_1536_u100 ( .A(mult_1536_n164), .B(mult_1536_n175), .Y(
        mult_1536_n141) );
  NOR2_X1M_A12TR mult_1536_u99 ( .A(mult_1536_n163), .B(mult_1536_n175), .Y(
        mult_1536_n140) );
  NOR2_X1M_A12TR mult_1536_u98 ( .A(mult_1536_n162), .B(mult_1536_n175), .Y(
        mult_1536_n139) );
  NOR2_X1M_A12TR mult_1536_u97 ( .A(mult_1536_n169), .B(mult_1536_n174), .Y(
        mult_1536_n138) );
  NOR2_X1M_A12TR mult_1536_u96 ( .A(mult_1536_n168), .B(mult_1536_n174), .Y(
        mult_1536_n137) );
  NOR2_X1M_A12TR mult_1536_u95 ( .A(mult_1536_n167), .B(mult_1536_n174), .Y(
        mult_1536_n136) );
  NOR2_X1M_A12TR mult_1536_u94 ( .A(mult_1536_n166), .B(mult_1536_n174), .Y(
        mult_1536_n135) );
  NOR2_X1M_A12TR mult_1536_u93 ( .A(mult_1536_n165), .B(mult_1536_n174), .Y(
        mult_1536_n134) );
  NOR2_X1M_A12TR mult_1536_u92 ( .A(mult_1536_n164), .B(mult_1536_n174), .Y(
        mult_1536_n133) );
  NOR2_X1M_A12TR mult_1536_u91 ( .A(mult_1536_n163), .B(mult_1536_n174), .Y(
        mult_1536_n132) );
  NOR2_X1M_A12TR mult_1536_u90 ( .A(mult_1536_n162), .B(mult_1536_n174), .Y(
        mult_1536_n131) );
  NOR2_X1M_A12TR mult_1536_u89 ( .A(mult_1536_n169), .B(mult_1536_n173), .Y(
        mult_1536_n130) );
  NOR2_X1M_A12TR mult_1536_u88 ( .A(mult_1536_n168), .B(mult_1536_n173), .Y(
        mult_1536_n129) );
  NOR2_X1M_A12TR mult_1536_u87 ( .A(mult_1536_n167), .B(mult_1536_n173), .Y(
        mult_1536_n128) );
  NOR2_X1M_A12TR mult_1536_u86 ( .A(mult_1536_n166), .B(mult_1536_n173), .Y(
        mult_1536_n127) );
  NOR2_X1M_A12TR mult_1536_u85 ( .A(mult_1536_n165), .B(mult_1536_n173), .Y(
        mult_1536_n126) );
  NOR2_X1M_A12TR mult_1536_u84 ( .A(mult_1536_n164), .B(mult_1536_n173), .Y(
        mult_1536_n125) );
  NOR2_X1M_A12TR mult_1536_u83 ( .A(mult_1536_n163), .B(mult_1536_n173), .Y(
        mult_1536_n124) );
  NOR2_X1M_A12TR mult_1536_u82 ( .A(mult_1536_n162), .B(mult_1536_n173), .Y(
        mult_1536_n123) );
  NOR2_X1M_A12TR mult_1536_u81 ( .A(mult_1536_n169), .B(mult_1536_n172), .Y(
        mult_1536_n122) );
  NOR2_X1M_A12TR mult_1536_u80 ( .A(mult_1536_n168), .B(mult_1536_n172), .Y(
        mult_1536_n121) );
  NOR2_X1M_A12TR mult_1536_u79 ( .A(mult_1536_n167), .B(mult_1536_n172), .Y(
        mult_1536_n120) );
  NOR2_X1M_A12TR mult_1536_u78 ( .A(mult_1536_n166), .B(mult_1536_n172), .Y(
        mult_1536_n119) );
  NOR2_X1M_A12TR mult_1536_u77 ( .A(mult_1536_n165), .B(mult_1536_n172), .Y(
        mult_1536_n118) );
  NOR2_X1M_A12TR mult_1536_u76 ( .A(mult_1536_n164), .B(mult_1536_n172), .Y(
        mult_1536_n117) );
  NOR2_X1M_A12TR mult_1536_u75 ( .A(mult_1536_n163), .B(mult_1536_n172), .Y(
        mult_1536_n116) );
  NOR2_X1M_A12TR mult_1536_u74 ( .A(mult_1536_n162), .B(mult_1536_n172), .Y(
        mult_1536_n115) );
  NOR2_X1M_A12TR mult_1536_u73 ( .A(mult_1536_n169), .B(mult_1536_n171), .Y(
        mult_1536_n114) );
  NOR2_X1M_A12TR mult_1536_u72 ( .A(mult_1536_n168), .B(mult_1536_n171), .Y(
        mult_1536_n113) );
  NOR2_X1M_A12TR mult_1536_u71 ( .A(mult_1536_n167), .B(mult_1536_n171), .Y(
        mult_1536_n112) );
  NOR2_X1M_A12TR mult_1536_u70 ( .A(mult_1536_n166), .B(mult_1536_n171), .Y(
        mult_1536_n111) );
  NOR2_X1M_A12TR mult_1536_u69 ( .A(mult_1536_n165), .B(mult_1536_n171), .Y(
        mult_1536_n110) );
  NOR2_X1M_A12TR mult_1536_u68 ( .A(mult_1536_n164), .B(mult_1536_n171), .Y(
        mult_1536_n109) );
  NOR2_X1M_A12TR mult_1536_u67 ( .A(mult_1536_n163), .B(mult_1536_n171), .Y(
        mult_1536_n108) );
  NOR2_X1M_A12TR mult_1536_u66 ( .A(mult_1536_n162), .B(mult_1536_n171), .Y(
        mult_1536_n107) );
  NOR2_X1M_A12TR mult_1536_u65 ( .A(mult_1536_n169), .B(mult_1536_n170), .Y(
        mult_1536_n106) );
  NOR2_X1M_A12TR mult_1536_u64 ( .A(mult_1536_n168), .B(mult_1536_n170), .Y(
        mult_1536_n105) );
  NOR2_X1M_A12TR mult_1536_u63 ( .A(mult_1536_n167), .B(mult_1536_n170), .Y(
        mult_1536_n104) );
  NOR2_X1M_A12TR mult_1536_u62 ( .A(mult_1536_n166), .B(mult_1536_n170), .Y(
        mult_1536_n103) );
  NOR2_X1M_A12TR mult_1536_u61 ( .A(mult_1536_n165), .B(mult_1536_n170), .Y(
        mult_1536_n102) );
  NOR2_X1M_A12TR mult_1536_u60 ( .A(mult_1536_n164), .B(mult_1536_n170), .Y(
        mult_1536_n101) );
  NOR2_X1M_A12TR mult_1536_u59 ( .A(mult_1536_n163), .B(mult_1536_n170), .Y(
        mult_1536_n100) );
  NOR2_X1M_A12TR mult_1536_u58 ( .A(mult_1536_n162), .B(mult_1536_n170), .Y(
        mult_1536_n99) );
  ADDH_X1M_A12TR mult_1536_u57 ( .A(mult_1536_n160), .B(mult_1536_n153), .CO(
        mult_1536_n97), .S(mult_1536_n98) );
  ADDH_X1M_A12TR mult_1536_u56 ( .A(mult_1536_n145), .B(mult_1536_n138), .CO(
        mult_1536_n95), .S(mult_1536_n96) );
  ADDF_X1M_A12TR mult_1536_u55 ( .A(mult_1536_n159), .B(mult_1536_n152), .CI(
        mult_1536_n97), .CO(mult_1536_n93), .S(mult_1536_n94) );
  ADDH_X1M_A12TR mult_1536_u54 ( .A(mult_1536_n137), .B(mult_1536_n130), .CO(
        mult_1536_n91), .S(mult_1536_n92) );
  ADDF_X1M_A12TR mult_1536_u53 ( .A(mult_1536_n158), .B(mult_1536_n144), .CI(
        mult_1536_n151), .CO(mult_1536_n89), .S(mult_1536_n90) );
  ADDF_X1M_A12TR mult_1536_u52 ( .A(mult_1536_n95), .B(mult_1536_n92), .CI(
        mult_1536_n90), .CO(mult_1536_n87), .S(mult_1536_n88) );
  ADDH_X1M_A12TR mult_1536_u51 ( .A(mult_1536_n129), .B(mult_1536_n122), .CO(
        mult_1536_n85), .S(mult_1536_n86) );
  ADDF_X1M_A12TR mult_1536_u50 ( .A(mult_1536_n157), .B(mult_1536_n136), .CI(
        mult_1536_n143), .CO(mult_1536_n83), .S(mult_1536_n84) );
  ADDF_X1M_A12TR mult_1536_u49 ( .A(mult_1536_n150), .B(mult_1536_n91), .CI(
        mult_1536_n89), .CO(mult_1536_n81), .S(mult_1536_n82) );
  ADDF_X1M_A12TR mult_1536_u48 ( .A(mult_1536_n86), .B(mult_1536_n84), .CI(
        mult_1536_n87), .CO(mult_1536_n79), .S(mult_1536_n80) );
  ADDH_X1M_A12TR mult_1536_u47 ( .A(mult_1536_n121), .B(mult_1536_n114), .CO(
        mult_1536_n77), .S(mult_1536_n78) );
  ADDF_X1M_A12TR mult_1536_u46 ( .A(mult_1536_n156), .B(mult_1536_n128), .CI(
        mult_1536_n135), .CO(mult_1536_n75), .S(mult_1536_n76) );
  ADDF_X1M_A12TR mult_1536_u45 ( .A(mult_1536_n149), .B(mult_1536_n142), .CI(
        mult_1536_n85), .CO(mult_1536_n73), .S(mult_1536_n74) );
  ADDF_X1M_A12TR mult_1536_u44 ( .A(mult_1536_n83), .B(mult_1536_n78), .CI(
        mult_1536_n76), .CO(mult_1536_n71), .S(mult_1536_n72) );
  ADDF_X1M_A12TR mult_1536_u43 ( .A(mult_1536_n81), .B(mult_1536_n74), .CI(
        mult_1536_n72), .CO(mult_1536_n69), .S(mult_1536_n70) );
  ADDH_X1M_A12TR mult_1536_u42 ( .A(mult_1536_n113), .B(mult_1536_n106), .CO(
        mult_1536_n67), .S(mult_1536_n68) );
  ADDF_X1M_A12TR mult_1536_u41 ( .A(mult_1536_n155), .B(mult_1536_n120), .CI(
        mult_1536_n127), .CO(mult_1536_n65), .S(mult_1536_n66) );
  ADDF_X1M_A12TR mult_1536_u40 ( .A(mult_1536_n148), .B(mult_1536_n134), .CI(
        mult_1536_n141), .CO(mult_1536_n63), .S(mult_1536_n64) );
  ADDF_X1M_A12TR mult_1536_u39 ( .A(mult_1536_n77), .B(mult_1536_n75), .CI(
        mult_1536_n68), .CO(mult_1536_n61), .S(mult_1536_n62) );
  ADDF_X1M_A12TR mult_1536_u38 ( .A(mult_1536_n64), .B(mult_1536_n66), .CI(
        mult_1536_n73), .CO(mult_1536_n59), .S(mult_1536_n60) );
  ADDF_X1M_A12TR mult_1536_u37 ( .A(mult_1536_n71), .B(mult_1536_n62), .CI(
        mult_1536_n60), .CO(mult_1536_n57), .S(mult_1536_n58) );
  ADDH_X1M_A12TR mult_1536_u36 ( .A(mult_1536_n112), .B(mult_1536_n105), .CO(
        mult_1536_n55), .S(mult_1536_n56) );
  ADDF_X1M_A12TR mult_1536_u35 ( .A(mult_1536_n147), .B(mult_1536_n119), .CI(
        mult_1536_n126), .CO(mult_1536_n53), .S(mult_1536_n54) );
  ADDF_X1M_A12TR mult_1536_u34 ( .A(mult_1536_n140), .B(mult_1536_n133), .CI(
        mult_1536_n67), .CO(mult_1536_n51), .S(mult_1536_n52) );
  ADDF_X1M_A12TR mult_1536_u33 ( .A(mult_1536_n65), .B(mult_1536_n63), .CI(
        mult_1536_n56), .CO(mult_1536_n49), .S(mult_1536_n50) );
  ADDF_X1M_A12TR mult_1536_u32 ( .A(mult_1536_n54), .B(mult_1536_n61), .CI(
        mult_1536_n52), .CO(mult_1536_n47), .S(mult_1536_n48) );
  ADDF_X1M_A12TR mult_1536_u31 ( .A(mult_1536_n59), .B(mult_1536_n50), .CI(
        mult_1536_n48), .CO(mult_1536_n45), .S(mult_1536_n46) );
  ADDF_X1M_A12TR mult_1536_u30 ( .A(mult_1536_n139), .B(mult_1536_n104), .CI(
        mult_1536_n111), .CO(mult_1536_n43), .S(mult_1536_n44) );
  ADDF_X1M_A12TR mult_1536_u29 ( .A(mult_1536_n118), .B(mult_1536_n125), .CI(
        mult_1536_n132), .CO(mult_1536_n41), .S(mult_1536_n42) );
  ADDF_X1M_A12TR mult_1536_u28 ( .A(mult_1536_n55), .B(mult_1536_n53), .CI(
        mult_1536_n42), .CO(mult_1536_n39), .S(mult_1536_n40) );
  ADDF_X1M_A12TR mult_1536_u27 ( .A(mult_1536_n44), .B(mult_1536_n51), .CI(
        mult_1536_n49), .CO(mult_1536_n37), .S(mult_1536_n38) );
  ADDF_X1M_A12TR mult_1536_u26 ( .A(mult_1536_n40), .B(mult_1536_n47), .CI(
        mult_1536_n38), .CO(mult_1536_n35), .S(mult_1536_n36) );
  ADDF_X1M_A12TR mult_1536_u25 ( .A(mult_1536_n131), .B(mult_1536_n103), .CI(
        mult_1536_n110), .CO(mult_1536_n33), .S(mult_1536_n34) );
  ADDF_X1M_A12TR mult_1536_u24 ( .A(mult_1536_n124), .B(mult_1536_n117), .CI(
        mult_1536_n43), .CO(mult_1536_n31), .S(mult_1536_n32) );
  ADDF_X1M_A12TR mult_1536_u23 ( .A(mult_1536_n41), .B(mult_1536_n34), .CI(
        mult_1536_n39), .CO(mult_1536_n29), .S(mult_1536_n30) );
  ADDF_X1M_A12TR mult_1536_u22 ( .A(mult_1536_n32), .B(mult_1536_n37), .CI(
        mult_1536_n30), .CO(mult_1536_n27), .S(mult_1536_n28) );
  ADDF_X1M_A12TR mult_1536_u21 ( .A(mult_1536_n123), .B(mult_1536_n102), .CI(
        mult_1536_n109), .CO(mult_1536_n25), .S(mult_1536_n26) );
  ADDF_X1M_A12TR mult_1536_u20 ( .A(mult_1536_n116), .B(mult_1536_n33), .CI(
        mult_1536_n26), .CO(mult_1536_n23), .S(mult_1536_n24) );
  ADDF_X1M_A12TR mult_1536_u19 ( .A(mult_1536_n31), .B(mult_1536_n24), .CI(
        mult_1536_n29), .CO(mult_1536_n21), .S(mult_1536_n22) );
  ADDF_X1M_A12TR mult_1536_u18 ( .A(mult_1536_n115), .B(mult_1536_n101), .CI(
        mult_1536_n108), .CO(mult_1536_n19), .S(mult_1536_n20) );
  ADDF_X1M_A12TR mult_1536_u17 ( .A(mult_1536_n25), .B(mult_1536_n20), .CI(
        mult_1536_n23), .CO(mult_1536_n17), .S(mult_1536_n18) );
  ADDF_X1M_A12TR mult_1536_u16 ( .A(mult_1536_n107), .B(mult_1536_n100), .CI(
        mult_1536_n19), .CO(mult_1536_n15), .S(mult_1536_n16) );
  ADDH_X1M_A12TR mult_1536_u15 ( .A(mult_1536_n154), .B(mult_1536_n161), .CO(
        mult_1536_n14), .S(n1783) );
  ADDF_X1M_A12TR mult_1536_u14 ( .A(mult_1536_n146), .B(mult_1536_n14), .CI(
        mult_1536_n98), .CO(mult_1536_n13), .S(n17840) );
  ADDF_X1M_A12TR mult_1536_u13 ( .A(mult_1536_n96), .B(mult_1536_n13), .CI(
        mult_1536_n94), .CO(mult_1536_n12), .S(n1785) );
  ADDF_X1M_A12TR mult_1536_u12 ( .A(mult_1536_n93), .B(mult_1536_n88), .CI(
        mult_1536_n12), .CO(mult_1536_n11), .S(n1786) );
  ADDF_X1M_A12TR mult_1536_u11 ( .A(mult_1536_n82), .B(mult_1536_n80), .CI(
        mult_1536_n11), .CO(mult_1536_n10), .S(n17870) );
  ADDF_X1M_A12TR mult_1536_u10 ( .A(mult_1536_n79), .B(mult_1536_n70), .CI(
        mult_1536_n10), .CO(mult_1536_n9), .S(n1788) );
  ADDF_X1M_A12TR mult_1536_u9 ( .A(mult_1536_n69), .B(mult_1536_n58), .CI(
        mult_1536_n9), .CO(mult_1536_n8), .S(n1789) );
  ADDF_X1M_A12TR mult_1536_u8 ( .A(mult_1536_n57), .B(mult_1536_n46), .CI(
        mult_1536_n8), .CO(mult_1536_n7), .S(n17900) );
  ADDF_X1M_A12TR mult_1536_u7 ( .A(mult_1536_n45), .B(mult_1536_n36), .CI(
        mult_1536_n7), .CO(mult_1536_n6), .S(n1791) );
  ADDF_X1M_A12TR mult_1536_u6 ( .A(mult_1536_n35), .B(mult_1536_n28), .CI(
        mult_1536_n6), .CO(mult_1536_n5), .S(n1792) );
  ADDF_X1M_A12TR mult_1536_u5 ( .A(mult_1536_n27), .B(mult_1536_n22), .CI(
        mult_1536_n5), .CO(mult_1536_n4), .S(n1793) );
  ADDF_X1M_A12TR mult_1536_u4 ( .A(mult_1536_n18), .B(mult_1536_n21), .CI(
        mult_1536_n4), .CO(mult_1536_n3), .S(n1794) );
  ADDF_X1M_A12TR mult_1536_u3 ( .A(mult_1536_n16), .B(mult_1536_n17), .CI(
        mult_1536_n3), .CO(mult_1536_n2), .S(n1795) );
  ADDF_X1M_A12TR mult_1536_u2 ( .A(mult_1536_n99), .B(mult_1536_n15), .CI(
        mult_1536_n2), .CO(n17970), .S(n1796) );
endmodule

