
module oc8051_top ( wb_rst_i, wb_clk_i, wbi_adr_o, wbi_dat_i, wbi_stb_o, 
        wbi_ack_i, wbi_cyc_o, wbi_err_i, wbd_dat_i, wbd_dat_o, wbd_adr_o, 
        wbd_we_o, wbd_ack_i, wbd_stb_o, wbd_cyc_o, wbd_err_i, int0_i, int1_i, 
        p0_i, p0_o, p1_i, p1_o, p2_i, p2_o, p3_i, p3_o, rxd_i, txd_o, t0_i, 
        t1_i, t2_i, t2ex_i, ea_in );
  output [15:0] wbi_adr_o;
  input [31:0] wbi_dat_i;
  input [7:0] wbd_dat_i;
  output [7:0] wbd_dat_o;
  output [15:0] wbd_adr_o;
  input [7:0] p0_i;
  output [7:0] p0_o;
  input [7:0] p1_i;
  output [7:0] p1_o;
  input [7:0] p2_i;
  output [7:0] p2_o;
  input [7:0] p3_i;
  output [7:0] p3_o;
  input wb_rst_i, wb_clk_i, wbi_ack_i, wbi_err_i, wbd_ack_i, wbd_err_i, int0_i,
         int1_i, rxd_i, t0_i, t1_i, t2_i, t2ex_i, ea_in;
  output wbi_stb_o, wbi_cyc_o, wbd_we_o, wbd_stb_o, wbd_cyc_o, txd_o;
  wire   wbi_stb_o, n_logic0_, wbd_cyc_o, src_sel3, pc_wr, eq, rd, rmw, istb,
         mem_wait, wait_data, alu_cy, srcac, descy, desac, desov, bit_out,
         bit_addr_o, n_0_net_, bit_data, wr_o, wr_ind, cy, sfr_bit, intr,
         int_ack, reti, n_3_net_, comp_wait, n_5_net_, n2,
         oc8051_decoder1_n444, oc8051_decoder1_n441, oc8051_decoder1_n440,
         oc8051_decoder1_n439, oc8051_decoder1_n438, oc8051_decoder1_n437,
         oc8051_decoder1_n436, oc8051_decoder1_n435, oc8051_decoder1_n434,
         oc8051_decoder1_n433, oc8051_decoder1_n432, oc8051_decoder1_n431,
         oc8051_decoder1_n430, oc8051_decoder1_n429, oc8051_decoder1_n428,
         oc8051_decoder1_n427, oc8051_decoder1_n426, oc8051_decoder1_n425,
         oc8051_decoder1_n411, oc8051_decoder1_n410, oc8051_decoder1_n409,
         oc8051_decoder1_n404, oc8051_decoder1_n387, oc8051_decoder1_n386,
         oc8051_decoder1_n385, oc8051_decoder1_n384, oc8051_decoder1_n383,
         oc8051_decoder1_n382, oc8051_decoder1_n381, oc8051_decoder1_n380,
         oc8051_decoder1_n379, oc8051_decoder1_n378, oc8051_decoder1_n377,
         oc8051_decoder1_n376, oc8051_decoder1_n375, oc8051_decoder1_n374,
         oc8051_decoder1_n373, oc8051_decoder1_n372, oc8051_decoder1_n371,
         oc8051_decoder1_n370, oc8051_decoder1_n369, oc8051_decoder1_n368,
         oc8051_decoder1_n367, oc8051_decoder1_n366, oc8051_decoder1_n365,
         oc8051_decoder1_n364, oc8051_decoder1_n363, oc8051_decoder1_n362,
         oc8051_decoder1_n361, oc8051_decoder1_n360, oc8051_decoder1_n359,
         oc8051_decoder1_n358, oc8051_decoder1_n357, oc8051_decoder1_n356,
         oc8051_decoder1_n355, oc8051_decoder1_n354, oc8051_decoder1_n353,
         oc8051_decoder1_n352, oc8051_decoder1_n351, oc8051_decoder1_n350,
         oc8051_decoder1_n349, oc8051_decoder1_n348, oc8051_decoder1_n347,
         oc8051_decoder1_n346, oc8051_decoder1_n345, oc8051_decoder1_n344,
         oc8051_decoder1_n343, oc8051_decoder1_n342, oc8051_decoder1_n341,
         oc8051_decoder1_n340, oc8051_decoder1_n339, oc8051_decoder1_n338,
         oc8051_decoder1_n337, oc8051_decoder1_n336, oc8051_decoder1_n335,
         oc8051_decoder1_n334, oc8051_decoder1_n333, oc8051_decoder1_n332,
         oc8051_decoder1_n331, oc8051_decoder1_n330, oc8051_decoder1_n329,
         oc8051_decoder1_n328, oc8051_decoder1_n327, oc8051_decoder1_n326,
         oc8051_decoder1_n325, oc8051_decoder1_n324, oc8051_decoder1_n323,
         oc8051_decoder1_n322, oc8051_decoder1_n321, oc8051_decoder1_n320,
         oc8051_decoder1_n319, oc8051_decoder1_n318, oc8051_decoder1_n317,
         oc8051_decoder1_n316, oc8051_decoder1_n315, oc8051_decoder1_n314,
         oc8051_decoder1_n313, oc8051_decoder1_n312, oc8051_decoder1_n311,
         oc8051_decoder1_n310, oc8051_decoder1_n309, oc8051_decoder1_n308,
         oc8051_decoder1_n307, oc8051_decoder1_n306, oc8051_decoder1_n305,
         oc8051_decoder1_n304, oc8051_decoder1_n303, oc8051_decoder1_n302,
         oc8051_decoder1_n301, oc8051_decoder1_n300, oc8051_decoder1_n299,
         oc8051_decoder1_n298, oc8051_decoder1_n297, oc8051_decoder1_n296,
         oc8051_decoder1_n295, oc8051_decoder1_n294, oc8051_decoder1_n293,
         oc8051_decoder1_n292, oc8051_decoder1_n291, oc8051_decoder1_n290,
         oc8051_decoder1_n289, oc8051_decoder1_n288, oc8051_decoder1_n287,
         oc8051_decoder1_n286, oc8051_decoder1_n285, oc8051_decoder1_n284,
         oc8051_decoder1_n283, oc8051_decoder1_n282, oc8051_decoder1_n281,
         oc8051_decoder1_n280, oc8051_decoder1_n279, oc8051_decoder1_n278,
         oc8051_decoder1_n277, oc8051_decoder1_n276, oc8051_decoder1_n275,
         oc8051_decoder1_n274, oc8051_decoder1_n273, oc8051_decoder1_n272,
         oc8051_decoder1_n271, oc8051_decoder1_n270, oc8051_decoder1_n269,
         oc8051_decoder1_n268, oc8051_decoder1_n267, oc8051_decoder1_n266,
         oc8051_decoder1_n265, oc8051_decoder1_n264, oc8051_decoder1_n263,
         oc8051_decoder1_n262, oc8051_decoder1_n261, oc8051_decoder1_n260,
         oc8051_decoder1_n259, oc8051_decoder1_n258, oc8051_decoder1_n257,
         oc8051_decoder1_n256, oc8051_decoder1_n255, oc8051_decoder1_n254,
         oc8051_decoder1_n253, oc8051_decoder1_n252, oc8051_decoder1_n251,
         oc8051_decoder1_n250, oc8051_decoder1_n249, oc8051_decoder1_n248,
         oc8051_decoder1_n247, oc8051_decoder1_n246, oc8051_decoder1_n245,
         oc8051_decoder1_n244, oc8051_decoder1_n243, oc8051_decoder1_n242,
         oc8051_decoder1_n241, oc8051_decoder1_n240, oc8051_decoder1_n239,
         oc8051_decoder1_n238, oc8051_decoder1_n237, oc8051_decoder1_n236,
         oc8051_decoder1_n235, oc8051_decoder1_n234, oc8051_decoder1_n233,
         oc8051_decoder1_n232, oc8051_decoder1_n231, oc8051_decoder1_n230,
         oc8051_decoder1_n229, oc8051_decoder1_n228, oc8051_decoder1_n227,
         oc8051_decoder1_n226, oc8051_decoder1_n225, oc8051_decoder1_n224,
         oc8051_decoder1_n223, oc8051_decoder1_n222, oc8051_decoder1_n221,
         oc8051_decoder1_n220, oc8051_decoder1_n219, oc8051_decoder1_n218,
         oc8051_decoder1_n217, oc8051_decoder1_n216, oc8051_decoder1_n215,
         oc8051_decoder1_n214, oc8051_decoder1_n213, oc8051_decoder1_n212,
         oc8051_decoder1_n211, oc8051_decoder1_n210, oc8051_decoder1_n209,
         oc8051_decoder1_n208, oc8051_decoder1_n207, oc8051_decoder1_n206,
         oc8051_decoder1_n205, oc8051_decoder1_n204, oc8051_decoder1_n203,
         oc8051_decoder1_n202, oc8051_decoder1_n201, oc8051_decoder1_n200,
         oc8051_decoder1_n199, oc8051_decoder1_n198, oc8051_decoder1_n197,
         oc8051_decoder1_n196, oc8051_decoder1_n195, oc8051_decoder1_n194,
         oc8051_decoder1_n193, oc8051_decoder1_n192, oc8051_decoder1_n191,
         oc8051_decoder1_n190, oc8051_decoder1_n189, oc8051_decoder1_n188,
         oc8051_decoder1_n187, oc8051_decoder1_n186, oc8051_decoder1_n185,
         oc8051_decoder1_n184, oc8051_decoder1_n183, oc8051_decoder1_n182,
         oc8051_decoder1_n181, oc8051_decoder1_n180, oc8051_decoder1_n179,
         oc8051_decoder1_n178, oc8051_decoder1_n177, oc8051_decoder1_n176,
         oc8051_decoder1_n175, oc8051_decoder1_n174, oc8051_decoder1_n173,
         oc8051_decoder1_n172, oc8051_decoder1_n171, oc8051_decoder1_n170,
         oc8051_decoder1_n169, oc8051_decoder1_n168, oc8051_decoder1_n167,
         oc8051_decoder1_n166, oc8051_decoder1_n165, oc8051_decoder1_n164,
         oc8051_decoder1_n163, oc8051_decoder1_n162, oc8051_decoder1_n161,
         oc8051_decoder1_n160, oc8051_decoder1_n159, oc8051_decoder1_n158,
         oc8051_decoder1_n157, oc8051_decoder1_n156, oc8051_decoder1_n155,
         oc8051_decoder1_n154, oc8051_decoder1_n153, oc8051_decoder1_n152,
         oc8051_decoder1_n151, oc8051_decoder1_n150, oc8051_decoder1_n149,
         oc8051_decoder1_n148, oc8051_decoder1_n147, oc8051_decoder1_n146,
         oc8051_decoder1_n145, oc8051_decoder1_n144, oc8051_decoder1_n143,
         oc8051_decoder1_n142, oc8051_decoder1_n141, oc8051_decoder1_n140,
         oc8051_decoder1_n139, oc8051_decoder1_n138, oc8051_decoder1_n137,
         oc8051_decoder1_n136, oc8051_decoder1_n135, oc8051_decoder1_n134,
         oc8051_decoder1_n133, oc8051_decoder1_n132, oc8051_decoder1_n131,
         oc8051_decoder1_n130, oc8051_decoder1_n129, oc8051_decoder1_n128,
         oc8051_decoder1_n127, oc8051_decoder1_n126, oc8051_decoder1_n125,
         oc8051_decoder1_n124, oc8051_decoder1_n123, oc8051_decoder1_n122,
         oc8051_decoder1_n121, oc8051_decoder1_n120, oc8051_decoder1_n119,
         oc8051_decoder1_n118, oc8051_decoder1_n117, oc8051_decoder1_n116,
         oc8051_decoder1_n115, oc8051_decoder1_n114, oc8051_decoder1_n113,
         oc8051_decoder1_n112, oc8051_decoder1_n111, oc8051_decoder1_n110,
         oc8051_decoder1_n109, oc8051_decoder1_n108, oc8051_decoder1_n107,
         oc8051_decoder1_n106, oc8051_decoder1_n105, oc8051_decoder1_n104,
         oc8051_decoder1_n103, oc8051_decoder1_n102, oc8051_decoder1_n101,
         oc8051_decoder1_n100, oc8051_decoder1_n99, oc8051_decoder1_n98,
         oc8051_decoder1_n97, oc8051_decoder1_n96, oc8051_decoder1_n95,
         oc8051_decoder1_n94, oc8051_decoder1_n93, oc8051_decoder1_n92,
         oc8051_decoder1_n91, oc8051_decoder1_n90, oc8051_decoder1_n89,
         oc8051_decoder1_n88, oc8051_decoder1_n87, oc8051_decoder1_n86,
         oc8051_decoder1_n85, oc8051_decoder1_n84, oc8051_decoder1_n83,
         oc8051_decoder1_n82, oc8051_decoder1_n81, oc8051_decoder1_n80,
         oc8051_decoder1_n79, oc8051_decoder1_n78, oc8051_decoder1_n77,
         oc8051_decoder1_n76, oc8051_decoder1_n75, oc8051_decoder1_n74,
         oc8051_decoder1_n73, oc8051_decoder1_n72, oc8051_decoder1_n71,
         oc8051_decoder1_n70, oc8051_decoder1_n69, oc8051_decoder1_n68,
         oc8051_decoder1_n67, oc8051_decoder1_n66, oc8051_decoder1_n65,
         oc8051_decoder1_n64, oc8051_decoder1_n63, oc8051_decoder1_n62,
         oc8051_decoder1_n61, oc8051_decoder1_n60, oc8051_decoder1_n59,
         oc8051_decoder1_n58, oc8051_decoder1_n57, oc8051_decoder1_n56,
         oc8051_decoder1_n55, oc8051_decoder1_n54, oc8051_decoder1_n53,
         oc8051_decoder1_n52, oc8051_decoder1_n51, oc8051_decoder1_n50,
         oc8051_decoder1_n49, oc8051_decoder1_n48, oc8051_decoder1_n47,
         oc8051_decoder1_n46, oc8051_decoder1_n45, oc8051_decoder1_n44,
         oc8051_decoder1_n43, oc8051_decoder1_n42, oc8051_decoder1_n41,
         oc8051_decoder1_n40, oc8051_decoder1_n39, oc8051_decoder1_n38,
         oc8051_decoder1_n37, oc8051_decoder1_n36, oc8051_decoder1_n35,
         oc8051_decoder1_n34, oc8051_decoder1_n33, oc8051_decoder1_n32,
         oc8051_decoder1_n31, oc8051_decoder1_n30, oc8051_decoder1_n29,
         oc8051_decoder1_n28, oc8051_decoder1_n27, oc8051_decoder1_n26,
         oc8051_decoder1_n25, oc8051_decoder1_n24, oc8051_decoder1_n23,
         oc8051_decoder1_n22, oc8051_decoder1_n21, oc8051_decoder1_n20,
         oc8051_decoder1_n19, oc8051_decoder1_n18, oc8051_decoder1_n17,
         oc8051_decoder1_n16, oc8051_decoder1_n15, oc8051_decoder1_n14,
         oc8051_decoder1_n13, oc8051_decoder1_n12, oc8051_decoder1_n11,
         oc8051_decoder1_n10, oc8051_decoder1_n9, oc8051_decoder1_n8,
         oc8051_decoder1_n7, oc8051_decoder1_n6, oc8051_decoder1_n5,
         oc8051_decoder1_n4, oc8051_decoder1_n3, oc8051_decoder1_n2,
         oc8051_decoder1_n1, oc8051_decoder1_n424, oc8051_decoder1_n423,
         oc8051_decoder1_n422, oc8051_decoder1_n421, oc8051_decoder1_n420,
         oc8051_decoder1_n419, oc8051_decoder1_n418, oc8051_decoder1_n417,
         oc8051_decoder1_n416, oc8051_decoder1_n415, oc8051_decoder1_n414,
         oc8051_decoder1_n413, oc8051_decoder1_n412, oc8051_decoder1_n408,
         oc8051_decoder1_n407, oc8051_decoder1_n406, oc8051_decoder1_n405,
         oc8051_decoder1_n403, oc8051_decoder1_n402, oc8051_decoder1_n401,
         oc8051_decoder1_n400, oc8051_decoder1_n399, oc8051_decoder1_n398,
         oc8051_decoder1_n397, oc8051_decoder1_n396, oc8051_decoder1_n395,
         oc8051_decoder1_n394, oc8051_decoder1_n393, oc8051_decoder1_n392,
         oc8051_decoder1_n391, oc8051_decoder1_n390, oc8051_decoder1_n389,
         oc8051_decoder1_n388, oc8051_decoder1_n1806, oc8051_decoder1_n1805,
         oc8051_decoder1_n1804, oc8051_decoder1_wr,
         oc8051_decoder1_ram_wr_sel_0_, oc8051_decoder1_ram_wr_sel_1_,
         oc8051_decoder1_ram_rd_sel_0_, oc8051_decoder1_ram_rd_sel_1_,
         oc8051_decoder1_alu_op_0_, oc8051_decoder1_alu_op_1_,
         oc8051_decoder1_alu_op_2_, oc8051_decoder1_alu_op_3_,
         oc8051_decoder1_state_0_, oc8051_decoder1_state_1_, oc8051_alu1_n225,
         oc8051_alu1_n224, oc8051_alu1_n223, oc8051_alu1_n222,
         oc8051_alu1_n221, oc8051_alu1_n220, oc8051_alu1_n219,
         oc8051_alu1_n216, oc8051_alu1_n215, oc8051_alu1_n214,
         oc8051_alu1_n213, oc8051_alu1_n212, oc8051_alu1_n211,
         oc8051_alu1_n210, oc8051_alu1_n209, oc8051_alu1_n208,
         oc8051_alu1_n207, oc8051_alu1_n206, oc8051_alu1_n205,
         oc8051_alu1_n204, oc8051_alu1_n201, oc8051_alu1_n200,
         oc8051_alu1_n199, oc8051_alu1_n198, oc8051_alu1_n197,
         oc8051_alu1_n196, oc8051_alu1_n195, oc8051_alu1_n194,
         oc8051_alu1_n193, oc8051_alu1_n192, oc8051_alu1_n191,
         oc8051_alu1_n190, oc8051_alu1_n189, oc8051_alu1_n188,
         oc8051_alu1_n187, oc8051_alu1_n186, oc8051_alu1_n185,
         oc8051_alu1_n184, oc8051_alu1_n183, oc8051_alu1_n182,
         oc8051_alu1_n181, oc8051_alu1_n180, oc8051_alu1_n179,
         oc8051_alu1_n178, oc8051_alu1_n177, oc8051_alu1_n173,
         oc8051_alu1_n172, oc8051_alu1_n171, oc8051_alu1_n170,
         oc8051_alu1_n169, oc8051_alu1_n168, oc8051_alu1_n167,
         oc8051_alu1_n166, oc8051_alu1_n165, oc8051_alu1_n164,
         oc8051_alu1_n163, oc8051_alu1_n162, oc8051_alu1_n161,
         oc8051_alu1_n160, oc8051_alu1_n159, oc8051_alu1_n158,
         oc8051_alu1_n157, oc8051_alu1_n156, oc8051_alu1_n155,
         oc8051_alu1_n154, oc8051_alu1_n153, oc8051_alu1_n152,
         oc8051_alu1_n151, oc8051_alu1_n150, oc8051_alu1_n149,
         oc8051_alu1_n148, oc8051_alu1_n147, oc8051_alu1_n146,
         oc8051_alu1_n145, oc8051_alu1_n144, oc8051_alu1_n143,
         oc8051_alu1_n142, oc8051_alu1_n141, oc8051_alu1_n140,
         oc8051_alu1_n139, oc8051_alu1_n136, oc8051_alu1_n135,
         oc8051_alu1_n134, oc8051_alu1_n133, oc8051_alu1_n132,
         oc8051_alu1_n131, oc8051_alu1_n130, oc8051_alu1_n129,
         oc8051_alu1_n128, oc8051_alu1_n127, oc8051_alu1_n126,
         oc8051_alu1_n125, oc8051_alu1_n123, oc8051_alu1_n121,
         oc8051_alu1_n120, oc8051_alu1_n119, oc8051_alu1_n118,
         oc8051_alu1_n117, oc8051_alu1_n116, oc8051_alu1_n115,
         oc8051_alu1_n114, oc8051_alu1_n113, oc8051_alu1_n112,
         oc8051_alu1_n111, oc8051_alu1_n110, oc8051_alu1_n109,
         oc8051_alu1_n108, oc8051_alu1_n107, oc8051_alu1_n106,
         oc8051_alu1_n105, oc8051_alu1_n104, oc8051_alu1_n103,
         oc8051_alu1_n102, oc8051_alu1_n101, oc8051_alu1_n100, oc8051_alu1_n99,
         oc8051_alu1_n98, oc8051_alu1_n97, oc8051_alu1_n96, oc8051_alu1_n95,
         oc8051_alu1_n94, oc8051_alu1_n93, oc8051_alu1_n92, oc8051_alu1_n90,
         oc8051_alu1_n89, oc8051_alu1_n88, oc8051_alu1_n86, oc8051_alu1_n85,
         oc8051_alu1_n84, oc8051_alu1_n83, oc8051_alu1_n82, oc8051_alu1_n81,
         oc8051_alu1_n80, oc8051_alu1_n79, oc8051_alu1_n78, oc8051_alu1_n77,
         oc8051_alu1_n76, oc8051_alu1_n75, oc8051_alu1_n74, oc8051_alu1_n73,
         oc8051_alu1_n72, oc8051_alu1_n71, oc8051_alu1_n70, oc8051_alu1_n69,
         oc8051_alu1_n68, oc8051_alu1_n67, oc8051_alu1_n66, oc8051_alu1_n65,
         oc8051_alu1_n64, oc8051_alu1_n63, oc8051_alu1_n62, oc8051_alu1_n61,
         oc8051_alu1_n60, oc8051_alu1_n59, oc8051_alu1_n58, oc8051_alu1_n57,
         oc8051_alu1_n56, oc8051_alu1_n55, oc8051_alu1_n54, oc8051_alu1_n53,
         oc8051_alu1_n52, oc8051_alu1_n51, oc8051_alu1_n50, oc8051_alu1_n49,
         oc8051_alu1_n48, oc8051_alu1_n47, oc8051_alu1_n46, oc8051_alu1_n45,
         oc8051_alu1_n44, oc8051_alu1_n43, oc8051_alu1_n42, oc8051_alu1_n41,
         oc8051_alu1_n40, oc8051_alu1_n39, oc8051_alu1_n38, oc8051_alu1_n37,
         oc8051_alu1_n36, oc8051_alu1_n35, oc8051_alu1_n34, oc8051_alu1_n33,
         oc8051_alu1_n32, oc8051_alu1_n31, oc8051_alu1_n30, oc8051_alu1_n29,
         oc8051_alu1_n28, oc8051_alu1_n27, oc8051_alu1_n26, oc8051_alu1_n25,
         oc8051_alu1_n24, oc8051_alu1_n23, oc8051_alu1_n22, oc8051_alu1_n21,
         oc8051_alu1_n20, oc8051_alu1_n19, oc8051_alu1_n18, oc8051_alu1_n17,
         oc8051_alu1_n16, oc8051_alu1_n15, oc8051_alu1_n13, oc8051_alu1_n12,
         oc8051_alu1_n11, oc8051_alu1_n10, oc8051_alu1_n9, oc8051_alu1_n8,
         oc8051_alu1_n7, oc8051_alu1_n6, oc8051_alu1_n5, oc8051_alu1_n4,
         oc8051_alu1_n3, oc8051_alu1_n2, oc8051_alu1_n1,
         oc8051_alu1_sub_1_root_sub_189_2_carry_3_,
         oc8051_alu1_sub_1_root_sub_189_2_carry_2_,
         oc8051_alu1_sub_1_root_sub_189_2_carry_1_,
         oc8051_alu1_sub_1_root_sub_189_2_carry_0_, oc8051_alu1_r450_carry_3_,
         oc8051_alu1_r450_carry_2_, oc8051_alu1_n247, oc8051_alu1_n246,
         oc8051_alu1_n245, oc8051_alu1_n244, oc8051_alu1_n243,
         oc8051_alu1_n237, oc8051_alu1_n236, oc8051_alu1_n228,
         oc8051_alu1_n227, oc8051_alu1_n218, oc8051_alu1_n217,
         oc8051_alu1_n203, oc8051_alu1_n202, oc8051_alu1_n176,
         oc8051_alu1_n175, oc8051_alu1_n174, oc8051_alu1_n138,
         oc8051_alu1_n137, oc8051_alu1_n124, oc8051_alu1_n122, oc8051_alu1_n91,
         oc8051_alu1_n87, oc8051_alu1_u3_u2_z_0, oc8051_alu1_u3_u1_z_2,
         oc8051_alu1_n14, oc8051_alu1_n240, oc8051_alu1_n2200,
         oc8051_alu1_n2190, oc8051_alu1_n2180, oc8051_alu1_n2170,
         oc8051_alu1_n2160, oc8051_alu1_n2150, oc8051_alu1_n2140,
         oc8051_alu1_n2130, oc8051_alu1_n1810, oc8051_alu1_n1800,
         oc8051_alu1_n1790, oc8051_alu1_n1780, oc8051_alu1_n1770,
         oc8051_alu1_n1520, oc8051_alu1_n1510, oc8051_alu1_n1410,
         oc8051_alu1_n1400, oc8051_alu1_n1390, oc8051_alu1_n1380,
         oc8051_alu1_n1370, oc8051_alu1_n1360, oc8051_alu1_n1350,
         oc8051_alu1_n1340, oc8051_alu1_sub4_4_, oc8051_alu1_addc_1_,
         oc8051_alu1_add4_0_, oc8051_alu1_add4_1_, oc8051_alu1_add4_2_,
         oc8051_alu1_add4_3_, oc8051_alu1_add4_4_, oc8051_alu1_divov,
         oc8051_alu1_mulov, oc8051_alu1_malicious1,
         oc8051_alu1_alu_malicious_n7, oc8051_alu1_alu_malicious_n6,
         oc8051_alu1_alu_malicious_n5, oc8051_alu1_alu_malicious_n4,
         oc8051_alu1_alu_malicious_n3, oc8051_alu1_alu_malicious_n2,
         oc8051_alu1_alu_malicious_n1, oc8051_alu1_alu_malicious_n9,
         oc8051_alu1_alu_malicious_n8, oc8051_alu1_alu_malicious_n70,
         oc8051_alu1_alu_malicious_state_0_,
         oc8051_alu1_alu_malicious_state_1_, oc8051_alu1_oc8051_mul1_n22,
         oc8051_alu1_oc8051_mul1_n21, oc8051_alu1_oc8051_mul1_n20,
         oc8051_alu1_oc8051_mul1_n19, oc8051_alu1_oc8051_mul1_n18,
         oc8051_alu1_oc8051_mul1_n16, oc8051_alu1_oc8051_mul1_n15,
         oc8051_alu1_oc8051_mul1_n14, oc8051_alu1_oc8051_mul1_n13,
         oc8051_alu1_oc8051_mul1_n12, oc8051_alu1_oc8051_mul1_n11,
         oc8051_alu1_oc8051_mul1_n10, oc8051_alu1_oc8051_mul1_n9,
         oc8051_alu1_oc8051_mul1_n8, oc8051_alu1_oc8051_mul1_n7,
         oc8051_alu1_oc8051_mul1_n6, oc8051_alu1_oc8051_mul1_n5,
         oc8051_alu1_oc8051_mul1_n4, oc8051_alu1_oc8051_mul1_n3,
         oc8051_alu1_oc8051_mul1_n2, oc8051_alu1_oc8051_mul1_n1,
         oc8051_alu1_oc8051_mul1_add_96_carry_10_,
         oc8051_alu1_oc8051_mul1_add_96_carry_9_,
         oc8051_alu1_oc8051_mul1_add_96_carry_8_,
         oc8051_alu1_oc8051_mul1_add_96_carry_7_,
         oc8051_alu1_oc8051_mul1_add_96_carry_6_,
         oc8051_alu1_oc8051_mul1_add_96_carry_5_,
         oc8051_alu1_oc8051_mul1_add_96_carry_4_,
         oc8051_alu1_oc8051_mul1_add_96_carry_3_, oc8051_alu1_oc8051_mul1_n17,
         oc8051_alu1_oc8051_mul1_shifted_2_,
         oc8051_alu1_oc8051_mul1_shifted_3_,
         oc8051_alu1_oc8051_mul1_shifted_4_,
         oc8051_alu1_oc8051_mul1_shifted_5_,
         oc8051_alu1_oc8051_mul1_shifted_6_,
         oc8051_alu1_oc8051_mul1_shifted_7_,
         oc8051_alu1_oc8051_mul1_shifted_8_,
         oc8051_alu1_oc8051_mul1_shifted_9_,
         oc8051_alu1_oc8051_mul1_shifted_10_,
         oc8051_alu1_oc8051_mul1_shifted_11_,
         oc8051_alu1_oc8051_mul1_shifted_12_,
         oc8051_alu1_oc8051_mul1_shifted_13_,
         oc8051_alu1_oc8051_mul1_shifted_14_,
         oc8051_alu1_oc8051_mul1_shifted_15_, oc8051_alu1_oc8051_mul1_n80,
         oc8051_alu1_oc8051_mul1_n70, oc8051_alu1_oc8051_mul1_cycle_0_,
         oc8051_alu1_oc8051_mul1_cycle_1_, oc8051_alu1_oc8051_mul1_mult_90_n33,
         oc8051_alu1_oc8051_mul1_mult_90_n32,
         oc8051_alu1_oc8051_mul1_mult_90_n31,
         oc8051_alu1_oc8051_mul1_mult_90_n30,
         oc8051_alu1_oc8051_mul1_mult_90_n29,
         oc8051_alu1_oc8051_mul1_mult_90_n28,
         oc8051_alu1_oc8051_mul1_mult_90_n27,
         oc8051_alu1_oc8051_mul1_mult_90_n26,
         oc8051_alu1_oc8051_mul1_mult_90_n25,
         oc8051_alu1_oc8051_mul1_mult_90_n24,
         oc8051_alu1_oc8051_mul1_mult_90_n23,
         oc8051_alu1_oc8051_mul1_mult_90_n22,
         oc8051_alu1_oc8051_mul1_mult_90_n21,
         oc8051_alu1_oc8051_mul1_mult_90_n20,
         oc8051_alu1_oc8051_mul1_mult_90_n19,
         oc8051_alu1_oc8051_mul1_mult_90_n18,
         oc8051_alu1_oc8051_mul1_mult_90_n17,
         oc8051_alu1_oc8051_mul1_mult_90_n16,
         oc8051_alu1_oc8051_mul1_mult_90_n15,
         oc8051_alu1_oc8051_mul1_mult_90_n14,
         oc8051_alu1_oc8051_mul1_mult_90_n13,
         oc8051_alu1_oc8051_mul1_mult_90_n12,
         oc8051_alu1_oc8051_mul1_mult_90_n11,
         oc8051_alu1_oc8051_mul1_mult_90_n10,
         oc8051_alu1_oc8051_mul1_mult_90_n9,
         oc8051_alu1_oc8051_mul1_mult_90_n8,
         oc8051_alu1_oc8051_mul1_mult_90_n7,
         oc8051_alu1_oc8051_mul1_mult_90_n6,
         oc8051_alu1_oc8051_mul1_mult_90_n5,
         oc8051_alu1_oc8051_mul1_mult_90_n4,
         oc8051_alu1_oc8051_mul1_mult_90_n3,
         oc8051_alu1_oc8051_mul1_mult_90_n2, oc8051_alu1_oc8051_div1_n30,
         oc8051_alu1_oc8051_div1_n29, oc8051_alu1_oc8051_div1_n28,
         oc8051_alu1_oc8051_div1_n27, oc8051_alu1_oc8051_div1_n24,
         oc8051_alu1_oc8051_div1_n23, oc8051_alu1_oc8051_div1_n22,
         oc8051_alu1_oc8051_div1_n21, oc8051_alu1_oc8051_div1_n20,
         oc8051_alu1_oc8051_div1_n19, oc8051_alu1_oc8051_div1_n18,
         oc8051_alu1_oc8051_div1_n17, oc8051_alu1_oc8051_div1_n16,
         oc8051_alu1_oc8051_div1_n15, oc8051_alu1_oc8051_div1_n14,
         oc8051_alu1_oc8051_div1_n13, oc8051_alu1_oc8051_div1_n12,
         oc8051_alu1_oc8051_div1_n11, oc8051_alu1_oc8051_div1_n10,
         oc8051_alu1_oc8051_div1_n9, oc8051_alu1_oc8051_div1_n8,
         oc8051_alu1_oc8051_div1_n7, oc8051_alu1_oc8051_div1_n6,
         oc8051_alu1_oc8051_div1_n5, oc8051_alu1_oc8051_div1_n4,
         oc8051_alu1_oc8051_div1_n3, oc8051_alu1_oc8051_div1_n2,
         oc8051_alu1_oc8051_div1_n26, oc8051_alu1_oc8051_div1_n25,
         oc8051_alu1_oc8051_div1_cmp1_0_, oc8051_alu1_oc8051_div1_rem1_0_,
         oc8051_alu1_oc8051_div1_rem1_1_, oc8051_alu1_oc8051_div1_rem1_2_,
         oc8051_alu1_oc8051_div1_rem1_3_, oc8051_alu1_oc8051_div1_rem1_4_,
         oc8051_alu1_oc8051_div1_rem1_5_, oc8051_alu1_oc8051_div1_rem1_6_,
         oc8051_alu1_oc8051_div1_rem1_7_, oc8051_alu1_oc8051_div1_rem2_1_,
         oc8051_alu1_oc8051_div1_rem2_2_, oc8051_alu1_oc8051_div1_rem2_3_,
         oc8051_alu1_oc8051_div1_rem2_4_, oc8051_alu1_oc8051_div1_rem2_5_,
         oc8051_alu1_oc8051_div1_rem2_6_, oc8051_alu1_oc8051_div1_rem2_7_,
         oc8051_alu1_oc8051_div1_cmp0_7_, oc8051_alu1_oc8051_div1_cmp1_1_,
         oc8051_alu1_oc8051_div1_cmp1_2_, oc8051_alu1_oc8051_div1_cmp1_3_,
         oc8051_alu1_oc8051_div1_cmp1_4_, oc8051_alu1_oc8051_div1_cmp1_5_,
         oc8051_alu1_oc8051_div1_cmp1_6_, oc8051_alu1_oc8051_div1_cmp1_7_,
         oc8051_alu1_oc8051_div1_cycle_0_, oc8051_alu1_oc8051_div1_cycle_1_,
         oc8051_alu1_oc8051_div1_sub_98_n1,
         oc8051_alu1_oc8051_div1_sub_98_b_not_0_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_1_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_2_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_3_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_4_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_5_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_6_,
         oc8051_alu1_oc8051_div1_sub_98_b_not_7_,
         oc8051_alu1_oc8051_div1_sub_94_n1, oc8051_alu1_sub_205_n14,
         oc8051_alu1_sub_205_n13, oc8051_alu1_sub_205_n12,
         oc8051_alu1_sub_205_n11, oc8051_alu1_sub_205_n10,
         oc8051_alu1_sub_205_n9, oc8051_alu1_sub_205_n8,
         oc8051_alu1_sub_205_n7, oc8051_alu1_sub_205_n6,
         oc8051_alu1_sub_205_n5, oc8051_alu1_sub_205_n4,
         oc8051_alu1_sub_205_n3, oc8051_alu1_sub_205_n2,
         oc8051_alu1_sub_205_n1, oc8051_ram_top1_n75, oc8051_ram_top1_n74,
         oc8051_ram_top1_n73, oc8051_ram_top1_n72, oc8051_ram_top1_n71,
         oc8051_ram_top1_n70, oc8051_ram_top1_n69, oc8051_ram_top1_n68,
         oc8051_ram_top1_n67, oc8051_ram_top1_n66, oc8051_ram_top1_n65,
         oc8051_ram_top1_n64, oc8051_ram_top1_n63, oc8051_ram_top1_n62,
         oc8051_ram_top1_n61, oc8051_ram_top1_n60, oc8051_ram_top1_n59,
         oc8051_ram_top1_n58, oc8051_ram_top1_n57, oc8051_ram_top1_n56,
         oc8051_ram_top1_n55, oc8051_ram_top1_n54, oc8051_ram_top1_n52,
         oc8051_ram_top1_n51, oc8051_ram_top1_n50, oc8051_ram_top1_n49,
         oc8051_ram_top1_n48, oc8051_ram_top1_n47, oc8051_ram_top1_n46,
         oc8051_ram_top1_n45, oc8051_ram_top1_n44, oc8051_ram_top1_n43,
         oc8051_ram_top1_n42, oc8051_ram_top1_n41, oc8051_ram_top1_n40,
         oc8051_ram_top1_n39, oc8051_ram_top1_n38, oc8051_ram_top1_n37,
         oc8051_ram_top1_n36, oc8051_ram_top1_n35, oc8051_ram_top1_n34,
         oc8051_ram_top1_n33, oc8051_ram_top1_n32, oc8051_ram_top1_n31,
         oc8051_ram_top1_n30, oc8051_ram_top1_n29, oc8051_ram_top1_n28,
         oc8051_ram_top1_n27, oc8051_ram_top1_n26, oc8051_ram_top1_n25,
         oc8051_ram_top1_n24, oc8051_ram_top1_n23, oc8051_ram_top1_n22,
         oc8051_ram_top1_n21, oc8051_ram_top1_n20, oc8051_ram_top1_n19,
         oc8051_ram_top1_n18, oc8051_ram_top1_n17, oc8051_ram_top1_n16,
         oc8051_ram_top1_n15, oc8051_ram_top1_n14, oc8051_ram_top1_n13,
         oc8051_ram_top1_n12, oc8051_ram_top1_n11, oc8051_ram_top1_n10,
         oc8051_ram_top1_n9, oc8051_ram_top1_n7, oc8051_ram_top1_n6,
         oc8051_ram_top1_n5, oc8051_ram_top1_n4, oc8051_ram_top1_n3,
         oc8051_ram_top1_n2, oc8051_ram_top1_n1, oc8051_ram_top1_n53,
         oc8051_ram_top1_n8, oc8051_ram_top1_bit_addr_r,
         oc8051_ram_top1_wr_addr_m_2_, oc8051_ram_top1_wr_addr_m_3_,
         oc8051_ram_top1_wr_addr_m_4_, oc8051_ram_top1_wr_addr_m_5_,
         oc8051_ram_top1_wr_addr_m_6_, oc8051_ram_top1_rd_addr_m_0_,
         oc8051_ram_top1_rd_addr_m_1_, oc8051_ram_top1_rd_addr_m_2_,
         oc8051_ram_top1_rd_addr_m_4_, oc8051_ram_top1_rd_addr_m_5_,
         oc8051_ram_top1_rd_addr_m_6_, oc8051_ram_top1_rd_en_r,
         oc8051_ram_top1__logic1_, oc8051_ram_top1_n280, oc8051_ram_top1_n270,
         oc8051_ram_top1_n260, oc8051_ram_top1_oc8051_idata__logic1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3432,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3431,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3430,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3428,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3424,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3419,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3417,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3416,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3415,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3413,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3411,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3409,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3408,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3342,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3324,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3255,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3237,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3219,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3218,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3183,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3182,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3164,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3163,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3123,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3122,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3121,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3120,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3119,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3118,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3117,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3116,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3115,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3114,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3113,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3112,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3111,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3110,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3109,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3108,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3107,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3106,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3105,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3104,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3103,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3102,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3101,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3100,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3099,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3098,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3097,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3096,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3095,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3094,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3093,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3092,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3091,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3090,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3089,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3088,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3087,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3086,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3085,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3084,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3083,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3082,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3081,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3080,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3079,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3078,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3077,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3076,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3075,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3074,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3073,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3072,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3071,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3070,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3069,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3068,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3067,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3066,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3065,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3064,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3063,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3062,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3061,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3060,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3059,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3058,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3057,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3056,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3055,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3054,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3053,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3052,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3051,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3050,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3049,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3048,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3047,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3046,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3045,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3044,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3043,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3042,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3041,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3040,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3039,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3038,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3037,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3036,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3035,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3034,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3033,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3032,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3031,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3030,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3029,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3028,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3027,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3026,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3025,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3024,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3023,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3022,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3021,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3020,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3019,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3018,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3017,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3016,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3015,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3014,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3013,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3012,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3011,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3010,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3009,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3008,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3007,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3006,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3005,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3004,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3003,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3002,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3001,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3000,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2999,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2998,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2997,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2996,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2995,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2994,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2993,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2992,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2991,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2990,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2989,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2988,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2987,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2986,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2985,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2984,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2983,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2982,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2981,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2980,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2979,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2978,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2977,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2976,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2975,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2974,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2973,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2972,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2971,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2970,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2969,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2968,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2967,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2966,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2965,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2964,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2963,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2962,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2961,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2960,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2959,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2958,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2957,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2956,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2955,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2954,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2953,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2952,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2951,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2950,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2949,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2948,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2947,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2946,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2945,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2944,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2943,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2942,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2941,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2940,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2939,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2938,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2937,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2936,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2935,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2934,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2933,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2932,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2931,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2930,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2929,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2928,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2927,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2926,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2925,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2924,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2923,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2922,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2921,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2920,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2919,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2918,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2917,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2916,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2915,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2914,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2913,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2912,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2911,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2910,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2909,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2908,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2907,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2906,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2905,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2904,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2903,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2902,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2901,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2900,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2899,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2898,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2897,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2896,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2895,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2894,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2893,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2892,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2891,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2890,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2889,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2888,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2887,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2886,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2885,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2884,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2883,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2882,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2881,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2880,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2879,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2878,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2877,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2876,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2875,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2874,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2873,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2872,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2871,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2870,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2869,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2868,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2867,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2866,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2865,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2864,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2863,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2862,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2861,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2860,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2859,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2858,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2857,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2856,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2855,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2854,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2853,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2852,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2851,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2850,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2849,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2848,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2847,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2846,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2845,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2844,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2843,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2842,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2841,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2840,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2839,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2838,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2837,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2836,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2835,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2834,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2833,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2832,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2831,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2830,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2829,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2828,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2827,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2826,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2825,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2824,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2823,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2822,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2821,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2820,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2819,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2818,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2817,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2816,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2815,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2814,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2813,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2812,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2811,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2810,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2809,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2808,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2807,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2806,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2805,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2804,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2803,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2802,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2801,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2800,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2799,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2798,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2797,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2796,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2795,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2794,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2793,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2792,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2791,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2790,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2789,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2788,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2787,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2786,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2785,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2784,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2783,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2782,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2781,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2780,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2779,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2778,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2777,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2776,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2775,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2774,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2773,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2772,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2771,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2770,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2769,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2768,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2767,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2766,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2765,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2764,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2763,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2762,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2761,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2760,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2759,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2758,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2757,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2756,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2755,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2754,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2753,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2752,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2751,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2750,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2749,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2748,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2747,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2746,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2745,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2744,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2743,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2742,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2741,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2740,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2739,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2738,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2737,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2736,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2735,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2734,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2733,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2732,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2731,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2730,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2729,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2728,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2727,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2726,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2725,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2724,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2723,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2722,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2721,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2720,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2719,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2718,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2717,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2716,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2715,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2714,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2713,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2712,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2711,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2710,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2709,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2708,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2707,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2706,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2705,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2704,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2703,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2702,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2701,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2700,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2699,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2698,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2697,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2696,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2695,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2694,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2693,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2692,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2691,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2690,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2689,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2688,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2687,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2686,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2685,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2684,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2683,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2682,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2681,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2680,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2679,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2678,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2677,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2676,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2675,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2674,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2673,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2672,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2671,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2670,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2669,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2668,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2667,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2666,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2665,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2664,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2663,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2662,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2661,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2660,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2659,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2658,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2657,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2656,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2655,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2654,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2653,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2652,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2651,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2650,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2649,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2648,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2647,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2646,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2645,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2644,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2643,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2642,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2641,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2640,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2639,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2638,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2637,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2636,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2635,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2634,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2633,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2632,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2631,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2630,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2629,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2628,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2627,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2626,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n568,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n567,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n566,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n565,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n564,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n563,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n562,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n561,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n560,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n559,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n558,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n557,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n556,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n555,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n554,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n553,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n552,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n551,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n550,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n549,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n548,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n547,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n546,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n545,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n544,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n543,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n542,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n541,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n540,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n539,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n538,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n537,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n536,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n535,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n534,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n533,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n532,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n531,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n530,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n529,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n528,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n527,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n526,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n525,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n524,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n523,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n522,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n521,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n520,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n519,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n518,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n517,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n516,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n515,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n514,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n513,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n512,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n511,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n510,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n509,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n508,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n507,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n506,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n505,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n504,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n503,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n502,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n501,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n500,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n499,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n498,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n497,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n496,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n495,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n494,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n493,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n492,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n491,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n490,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n489,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n488,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n487,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n486,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n485,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n484,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n483,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n482,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n481,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n480,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n479,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n478,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n477,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n476,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n475,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n474,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n473,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n472,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n471,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n470,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n469,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n468,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n467,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n466,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n465,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n464,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n463,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n462,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n461,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n460,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n459,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n458,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n457,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n456,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n455,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n454,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n453,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n452,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n451,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n450,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n449,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n448,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n447,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n446,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n445,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n444,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n443,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n442,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n441,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n440,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n439,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n438,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n437,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n436,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n435,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n434,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n433,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n432,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n431,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n430,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n429,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n428,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n427,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n426,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n425,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n424,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n423,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n422,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n421,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n420,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n419,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n418,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n417,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n416,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n415,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n414,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n413,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n412,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n411,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n410,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n409,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n408,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n407,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n406,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n405,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n404,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n403,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n402,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n401,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n400,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n399,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n398,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n397,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n396,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n395,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n374,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n373,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n372,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n371,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n370,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n369,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n368,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n367,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n366,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n365,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n364,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n363,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n362,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n361,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n360,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n359,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n358,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n357,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n356,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n355,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n354,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n353,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n352,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n351,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n350,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n349,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n348,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n307,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n306,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n305,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n304,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n303,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n302,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n301,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n300,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n299,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n298,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n297,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n296,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n295,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n294,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n293,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n292,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n291,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n290,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n289,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n288,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n287,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n286,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n285,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n284,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n283,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n282,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n281,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n240,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n239,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n238,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n237,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n236,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n235,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n234,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n233,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n232,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n231,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n210,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n209,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n208,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n207,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n206,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n205,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n204,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n203,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n202,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n201,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n180,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n179,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n178,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n177,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n176,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n175,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n174,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n173,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n172,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n171,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n150,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n149,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n148,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n147,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n146,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n145,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n144,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n143,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n142,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n141,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n120,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n119,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n118,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n117,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n116,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n115,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n114,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n113,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n112,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n111,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n90,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n89,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n88,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n87,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n86,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n85,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n84,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n83,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n82,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n81,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n60,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n59,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n58,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n57,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n56,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n55,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n54,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n53,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n52,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n51,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n30,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n29,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n28,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n27,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n26,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n25,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n24,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n23,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n22,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n21,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2625,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2624,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2623,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2622,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2621,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2620,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2619,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2618,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2617,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2616,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2615,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2614,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2613,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2612,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2611,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2610,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2609,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2608,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2607,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2606,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2605,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2604,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2603,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2602,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2601,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2600,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2599,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2598,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2597,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2596,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2595,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2594,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2593,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2592,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2591,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2590,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2589,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2588,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2587,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2586,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2585,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2584,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2583,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2582,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2581,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2580,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2579,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2578,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2577,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2576,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2575,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2574,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2573,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2572,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2571,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2570,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2569,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2568,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2567,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2566,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2565,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2564,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2563,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2562,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2561,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2560,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2559,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2558,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2557,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2556,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2555,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2554,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2553,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2552,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2551,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2550,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2549,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2548,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2547,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2546,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2545,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2544,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2543,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2542,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2541,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2540,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2539,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2538,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2537,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2536,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2535,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2534,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2533,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2532,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2531,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2530,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2529,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2528,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2527,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2526,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2525,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2524,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2523,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2522,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2521,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2520,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2519,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2518,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2517,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2516,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2515,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2514,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2513,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2512,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2511,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2510,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2509,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2508,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2507,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2506,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2505,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2504,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2503,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2502,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2501,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2500,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2499,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2498,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2497,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2496,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2495,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2494,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2493,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2492,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2491,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2490,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2489,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2488,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2487,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2486,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2485,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2484,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2483,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2482,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2481,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2480,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2479,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2478,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2477,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2476,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2475,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2474,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2473,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2472,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2471,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2470,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2469,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2468,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2467,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2466,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2465,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2464,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2463,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2462,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2461,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2460,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2459,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2458,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2457,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2456,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2455,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2454,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2453,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2452,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2451,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2450,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2449,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2448,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2447,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2446,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2445,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2444,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2443,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2442,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2441,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2440,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2439,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2438,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2437,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2436,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2435,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2434,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2433,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2432,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2431,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2430,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2429,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2428,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2427,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2426,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2425,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2424,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2423,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2422,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2421,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2420,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2419,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2418,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2417,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2416,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2415,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2414,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2413,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2412,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2411,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2410,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2409,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2408,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2407,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2406,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2405,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2404,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2403,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2402,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2401,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2400,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2399,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2398,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2397,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2396,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2395,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2394,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2393,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2392,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2391,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2390,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2389,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2388,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2387,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2386,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2385,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2384,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2383,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2382,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2381,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2380,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2379,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2378,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2377,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2376,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2375,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2374,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2373,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2372,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2371,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2370,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2369,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2368,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2367,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2366,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2365,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2364,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2363,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2362,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2361,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2360,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2359,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2358,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2357,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2356,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2355,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2354,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2353,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2352,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2351,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2350,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2349,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2348,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2347,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2346,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2345,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2344,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2343,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2342,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2341,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2340,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2339,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2338,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2337,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2336,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2335,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2334,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2333,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2332,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2331,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2330,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2329,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2328,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2327,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2326,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2325,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2324,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2323,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2322,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2321,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2320,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2319,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2318,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2317,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2316,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2315,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2314,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2313,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2312,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2311,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2310,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2309,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2308,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2307,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2306,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2305,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2304,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2303,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2302,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2301,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2300,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2299,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2298,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2297,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2296,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2295,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2294,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2293,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2292,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2291,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2290,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2289,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2288,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2287,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2286,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2285,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2284,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2283,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2282,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2281,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2280,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2279,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2278,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2277,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2276,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2275,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2274,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2273,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2272,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2271,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2270,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2269,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2268,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2267,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2266,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2265,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2264,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2263,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2262,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2261,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2260,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2259,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2258,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2257,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2256,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2255,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2254,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2253,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2252,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2251,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2250,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2249,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2248,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2247,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2246,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2245,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2244,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2243,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2242,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2241,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2240,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2239,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2238,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2237,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2236,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2235,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2234,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2233,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2232,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2231,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2230,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2229,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2228,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2227,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2226,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2225,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2224,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2223,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2222,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2221,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2220,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2219,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2218,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2217,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2216,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2215,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2214,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2213,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2212,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2211,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2210,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2209,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2208,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2207,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2206,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2205,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2204,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2203,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2202,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2201,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2200,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2199,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2198,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2197,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2196,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2195,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2194,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2193,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2192,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2191,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2190,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2189,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2188,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2187,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2186,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2185,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2184,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2183,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2182,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2181,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2180,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2179,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2178,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2177,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2176,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2175,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2174,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2173,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2172,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2171,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2170,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2169,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2168,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2167,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2166,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2165,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2164,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2163,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2162,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2161,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2160,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2159,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2158,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2157,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2156,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2155,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2154,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2153,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2152,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2151,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2150,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2149,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2148,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2147,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2146,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2145,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2144,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2143,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2142,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2141,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2140,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2139,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2138,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2137,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2136,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2135,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2134,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2133,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2132,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2131,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2130,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2129,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2128,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2127,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2126,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2125,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2124,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2123,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2122,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2121,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2120,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2119,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2118,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2117,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2116,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2115,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2114,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2113,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2112,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2111,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2110,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2109,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2108,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2107,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2106,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2105,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2104,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2103,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2102,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2101,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2100,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2099,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2098,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2097,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2096,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2095,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2094,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2093,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2092,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2091,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2090,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2089,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2088,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2087,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2086,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2085,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2084,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2083,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2082,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2081,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2080,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2079,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2078,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2077,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2076,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2075,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2074,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2073,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2072,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2071,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2070,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2069,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2068,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2067,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2066,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2065,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2064,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2063,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2062,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2061,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2060,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2059,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2058,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2057,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2056,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2055,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2054,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2053,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2052,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2051,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2050,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2049,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2048,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2047,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2046,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2045,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2044,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2043,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2042,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2041,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2040,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2039,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2038,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2037,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2036,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2035,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2034,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2033,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2032,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2031,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2030,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2029,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2028,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2027,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2026,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2025,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2024,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2023,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2022,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2021,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2020,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2019,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2018,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2017,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2016,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2015,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2014,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2013,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2012,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2011,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2010,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2009,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2008,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2007,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2006,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2005,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2004,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2003,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2002,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2001,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2000,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1999,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1998,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1997,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1996,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1995,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1994,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1993,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1992,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1991,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1990,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1989,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1988,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1987,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1986,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1985,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1984,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1983,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1982,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1981,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1980,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1979,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1978,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1977,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1976,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1975,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1974,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1973,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1972,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1971,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1970,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1969,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1968,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1967,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1966,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1965,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1964,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1963,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1962,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1961,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1960,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1959,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1958,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1957,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1956,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1955,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1954,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1953,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1952,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1951,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1950,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1949,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1948,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1947,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1946,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1945,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1944,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1943,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1942,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1941,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1940,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1939,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1938,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1937,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1936,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1935,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1934,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1933,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1932,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1931,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1930,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1929,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1928,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1927,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1926,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1925,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1924,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1923,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1922,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1921,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1920,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1919,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1918,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1917,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1916,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1915,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1914,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1913,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1912,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1911,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1910,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1909,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1908,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1907,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1906,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1905,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1904,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1903,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1902,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1901,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1900,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1899,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1898,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1897,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1896,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1895,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1894,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1893,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1892,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1891,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1890,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1889,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1888,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1887,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1886,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1885,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1884,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1883,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1882,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1881,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1880,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1879,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1878,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1877,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1876,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1875,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1874,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1873,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1872,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1871,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1870,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1869,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1868,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1867,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1866,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1865,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1864,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1863,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1862,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1861,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1860,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1859,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1858,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1857,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1856,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1855,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1854,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1853,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1852,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1851,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1850,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1849,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1848,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1847,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1846,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1845,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1844,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1843,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1842,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1841,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1840,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1839,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1838,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1837,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1836,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1835,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1834,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1833,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1832,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1831,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1830,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1829,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1828,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1827,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1826,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1825,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1824,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1823,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1822,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1821,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1820,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1819,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1818,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1817,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1816,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1815,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1814,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1813,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1812,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1811,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1810,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1809,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1808,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1807,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1806,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1805,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1804,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1803,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1802,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1801,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1800,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1799,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1798,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1797,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1796,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1795,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1794,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1793,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1792,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1791,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1790,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1789,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1788,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1787,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1786,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1785,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1784,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1783,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1782,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1781,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1780,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1779,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1778,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1777,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1776,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1775,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1774,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1773,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1772,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1771,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1770,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1769,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1768,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1767,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1766,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1765,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1764,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1763,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1762,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1761,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1760,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1759,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1758,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1757,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1756,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1755,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1754,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1753,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1752,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1751,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1750,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1749,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1748,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1747,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1746,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1745,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1744,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1743,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1742,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1741,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1740,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1739,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1738,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1737,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1736,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1735,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1734,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1733,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1732,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1731,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1730,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1729,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1728,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1727,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1726,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1725,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1724,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1723,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1722,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1721,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1720,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1719,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1718,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1717,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1716,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1715,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1714,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1713,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1712,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1711,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1710,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1709,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1708,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1707,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1706,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1705,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1704,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1703,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1702,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1701,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1700,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1699,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1698,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1697,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1696,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1695,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1694,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1693,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1692,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1691,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1690,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1689,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1688,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1687,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1686,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1685,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1684,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1683,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1682,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1681,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1680,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1679,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1678,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1677,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1676,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1675,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1674,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1673,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1672,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1671,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1670,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1669,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1668,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1667,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1666,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1665,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1664,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1663,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1662,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1661,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1660,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1659,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1658,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1657,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1656,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1655,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1654,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1653,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1652,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1651,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1650,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1649,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1648,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1647,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1646,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1645,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1644,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1643,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1642,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1641,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1640,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1639,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1638,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1637,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1636,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1635,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1634,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1633,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1632,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1631,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1630,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1629,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1628,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1627,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1626,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1625,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1624,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1623,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1622,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1621,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1620,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1619,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1618,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1617,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1616,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1615,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1614,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1613,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1612,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1611,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1610,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1609,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1608,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1607,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1606,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1605,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1604,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1603,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1602,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1601,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1600,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1599,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1598,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1597,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1596,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1595,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1594,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1593,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1592,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1591,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1590,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1589,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1588,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1587,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1586,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1585,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1584,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1583,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1582,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1581,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1580,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1579,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1578,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1577,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1576,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1575,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1574,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1573,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1572,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1571,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1570,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1569,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1568,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1567,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1566,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1565,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1564,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1563,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1562,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1561,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1560,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1559,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1558,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1557,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1556,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1555,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1554,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1553,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1552,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1551,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1550,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1549,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1548,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1547,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1546,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1545,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1544,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1543,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1542,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1541,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1540,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1539,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1538,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1537,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1536,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1535,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1534,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1533,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1532,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1531,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1530,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1529,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1528,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1527,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1526,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1525,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1524,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1523,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1522,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1521,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1520,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1519,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1518,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1517,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1516,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1515,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1514,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1513,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1512,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1511,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1510,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1509,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1508,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1507,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1506,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1505,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1504,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1503,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1502,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1501,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1500,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1499,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1498,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1497,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1496,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1495,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1494,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1493,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1492,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1491,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1490,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1489,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1488,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1487,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1486,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1485,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1484,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1483,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1482,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1481,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1480,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1479,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1478,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1477,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1476,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1475,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1474,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1473,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1472,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1471,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1470,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1469,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1468,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1467,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1466,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1465,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1464,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1463,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1462,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1461,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1460,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1459,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1458,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1457,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1456,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1455,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1454,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1453,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1452,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1451,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1450,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1449,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1448,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1447,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1446,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1445,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1444,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1443,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1442,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1441,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1440,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1439,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1438,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1437,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1436,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1435,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1434,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1433,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1432,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1431,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1430,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1429,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1428,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1427,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1426,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1425,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1424,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1423,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1422,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1421,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1420,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1419,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1418,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1417,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1416,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1415,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1414,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1413,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1412,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1411,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1410,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1409,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1408,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1407,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1406,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1405,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1404,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1403,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1402,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1401,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1400,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1399,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1398,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1397,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1396,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1395,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1394,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1393,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1392,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1391,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1390,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1389,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1388,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1387,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1386,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1385,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1384,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1383,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1382,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1381,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1380,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1379,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1378,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1377,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1376,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1375,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1374,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1373,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1372,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1371,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1370,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1369,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1368,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1367,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1366,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1365,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1364,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1363,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1362,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1361,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1360,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1359,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1358,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1357,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1356,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1355,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1354,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1353,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1352,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1351,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1350,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1349,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1348,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1347,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1346,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1345,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1344,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1343,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1342,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1341,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1340,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1339,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1338,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1337,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1336,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1335,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1334,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1333,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1332,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1331,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1330,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1329,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1328,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1327,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1326,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1325,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1324,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1323,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1322,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1321,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1320,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1319,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1318,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1317,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1316,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1315,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1314,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1313,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1312,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1311,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1310,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1309,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1308,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1307,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1306,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1305,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1304,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1303,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1302,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1301,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1300,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1299,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1298,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1297,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1296,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1295,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1294,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1293,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1292,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1291,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1290,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1289,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1288,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1287,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1286,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1285,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1284,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1283,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1282,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1281,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1280,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1279,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1278,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1277,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1276,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1275,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1274,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1273,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1272,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1271,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1270,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1269,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1268,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1267,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1266,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1265,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1264,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1263,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1262,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1261,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1260,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1259,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1258,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1257,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1256,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1255,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1254,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1253,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1252,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1251,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1250,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1249,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1248,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1247,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1246,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1245,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1244,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1243,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1242,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1241,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1240,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1239,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1238,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1237,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1236,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1235,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1234,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1233,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1232,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1231,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1230,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1229,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1228,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1227,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1226,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1225,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1224,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1223,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1222,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1221,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1220,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1219,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1218,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1217,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1216,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1215,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1214,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1213,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1212,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1211,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1210,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1209,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1208,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1207,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1206,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1205,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1204,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1203,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1202,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1201,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1200,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1199,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1198,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1197,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1196,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1195,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1194,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1193,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1192,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1191,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1190,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1189,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1188,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1187,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1186,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1185,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1184,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1183,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1182,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1181,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1180,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1179,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1178,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1177,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1176,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1175,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1174,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1173,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1172,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1171,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1170,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1169,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1168,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1167,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1166,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1165,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1164,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1163,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1162,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1161,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1160,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1159,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1158,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1157,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1156,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1155,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1154,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1153,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1152,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1151,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1150,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1149,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1148,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1147,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1146,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1145,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1144,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1143,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1142,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1141,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1140,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1139,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1138,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1137,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1136,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1135,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1134,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1133,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1132,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1131,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1130,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1129,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1128,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1127,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1126,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1125,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1124,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1123,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1122,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1121,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1120,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1119,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1118,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1117,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1116,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1115,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1114,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1113,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1112,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1111,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1110,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1109,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1108,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1107,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1106,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1105,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1104,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1103,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1102,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1101,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1100,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1099,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1098,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1097,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1096,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1095,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1094,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1093,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1092,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1091,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1090,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1089,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1088,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1087,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1086,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1085,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1084,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1083,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1082,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1081,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1080,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1079,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1078,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1077,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1076,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1075,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1074,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1073,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1072,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1071,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1070,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1069,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1068,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1067,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1066,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1065,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1064,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1063,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1062,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1061,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1060,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1059,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1058,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1057,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1056,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1055,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1054,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1053,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1052,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1051,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1050,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1049,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1048,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1047,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1046,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1045,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1044,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1043,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1042,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1041,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1040,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1039,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1038,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1037,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1036,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1035,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1034,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1033,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1032,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1031,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1030,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1029,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1028,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1027,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1026,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1025,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1024,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1023,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1022,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1021,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1020,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1019,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1018,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1017,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1016,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1015,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1014,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1013,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1012,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1011,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1010,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1009,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1008,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1007,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1006,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1005,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1004,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1003,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1002,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1001,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1000,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n999,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n998,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n997,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n996,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n995,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n994,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n993,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n992,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n991,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n990,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n989,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n988,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n987,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n986,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n985,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n984,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n983,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n982,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n981,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n980,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n979,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n978,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n977,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n976,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n975,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n974,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n973,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n972,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n971,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n970,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n969,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n968,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n967,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n966,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n965,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n964,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n963,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n962,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n961,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n960,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n959,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n958,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n957,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n956,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n955,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n954,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n953,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n952,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n951,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n950,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n949,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n948,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n947,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n946,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n945,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n944,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n943,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n942,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n941,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n940,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n939,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n938,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n937,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n936,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n935,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n934,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n933,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n932,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n931,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n930,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n929,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n928,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n927,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n926,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n925,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n924,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n923,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n922,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n921,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n920,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n919,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n918,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n917,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n916,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n915,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n914,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n913,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n912,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n911,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n910,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n909,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n908,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n907,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n906,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n905,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n904,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n903,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n902,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n901,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n900,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n899,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n898,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n897,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n896,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n895,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n894,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n893,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n892,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n891,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n890,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n889,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n888,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n887,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n886,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n885,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n884,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n883,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n882,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n881,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n880,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n879,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n878,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n877,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n876,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n875,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n874,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n873,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n872,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n871,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n870,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n869,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n868,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n867,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n866,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n865,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n864,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n863,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n862,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n861,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n860,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n859,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n858,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n857,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n856,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n855,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n854,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n853,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n852,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n851,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n850,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n849,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n848,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n847,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n846,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n845,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n844,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n843,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n842,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n841,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n840,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n839,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n838,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n837,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n836,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n835,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n834,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n833,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n832,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n831,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n830,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n829,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n828,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n827,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n826,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n825,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n824,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n823,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n822,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n821,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n820,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n819,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n818,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n817,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n816,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n815,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n814,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n813,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n812,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n811,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n810,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n809,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n808,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n807,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n806,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n805,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n804,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n803,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n802,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n801,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n800,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n799,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n798,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n797,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n796,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n795,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n794,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n793,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n792,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n791,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n790,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n789,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n788,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n787,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n786,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n785,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n784,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n783,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n782,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n781,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n780,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n779,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n778,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n777,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n776,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n775,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n774,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n773,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n772,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n771,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n770,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n769,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n768,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n767,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n766,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n765,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n764,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n763,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n762,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n761,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n760,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n759,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n758,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n757,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n756,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n755,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n754,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n753,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n752,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n751,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n750,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n749,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n748,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n747,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n746,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n745,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n744,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n743,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n742,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n741,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n740,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n739,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n738,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n737,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n736,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n735,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n734,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n733,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n732,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n731,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n730,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n729,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n728,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n727,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n726,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n725,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n724,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n723,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n722,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n721,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n720,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n719,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n718,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n717,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n716,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n715,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n714,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n713,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n712,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n711,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n710,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n709,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n708,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n707,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n706,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n705,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n704,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n703,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n702,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n701,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n700,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n699,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n698,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n697,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n696,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n695,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n694,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n693,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n692,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n691,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n690,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n689,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n688,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n687,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n686,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n685,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n684,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n683,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n682,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n681,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n680,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n679,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n678,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n677,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n676,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n675,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n674,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n673,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n672,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n671,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n670,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n669,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n668,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n667,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n666,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n665,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n664,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n663,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n662,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n661,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n660,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n659,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n658,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n657,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n656,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n655,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n654,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n653,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n652,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n651,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n650,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n649,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n648,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n647,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n646,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n645,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n644,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n643,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n642,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n641,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n640,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n639,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n638,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n637,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n636,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n635,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n634,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n633,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n632,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n631,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n630,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n629,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n628,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n627,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n626,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n625,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n624,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n623,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n622,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n621,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n620,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n619,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n618,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n617,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n616,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n615,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n614,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n613,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n612,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n611,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n610,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n609,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n608,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n607,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n606,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n605,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n604,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n603,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n602,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n601,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n600,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n599,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n598,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n597,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n596,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n595,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n594,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n593,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n592,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n591,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n590,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n589,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n588,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n587,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n586,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n585,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n584,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n583,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n582,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n581,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n580,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n579,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n578,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n577,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n576,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n575,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n574,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n573,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n572,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n571,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n570,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4110,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4010,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3910,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3810,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3710,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3610,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3510,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3435,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__7_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_0_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_1_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_2_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_3_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_4_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_5_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_6_,
         oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_7_,
         oc8051_alu_src_sel1_n61, oc8051_alu_src_sel1_n60,
         oc8051_alu_src_sel1_n59, oc8051_alu_src_sel1_n58,
         oc8051_alu_src_sel1_n57, oc8051_alu_src_sel1_n56,
         oc8051_alu_src_sel1_n55, oc8051_alu_src_sel1_n54,
         oc8051_alu_src_sel1_n53, oc8051_alu_src_sel1_n52,
         oc8051_alu_src_sel1_n51, oc8051_alu_src_sel1_n50,
         oc8051_alu_src_sel1_n49, oc8051_alu_src_sel1_n48,
         oc8051_alu_src_sel1_n47, oc8051_alu_src_sel1_n46,
         oc8051_alu_src_sel1_n45, oc8051_alu_src_sel1_n44,
         oc8051_alu_src_sel1_n43, oc8051_alu_src_sel1_n42,
         oc8051_alu_src_sel1_n41, oc8051_alu_src_sel1_n40,
         oc8051_alu_src_sel1_n39, oc8051_alu_src_sel1_n38,
         oc8051_alu_src_sel1_n37, oc8051_alu_src_sel1_n36,
         oc8051_alu_src_sel1_n35, oc8051_alu_src_sel1_n34,
         oc8051_alu_src_sel1_n33, oc8051_alu_src_sel1_n32,
         oc8051_alu_src_sel1_n28, oc8051_alu_src_sel1_n27,
         oc8051_alu_src_sel1_n26, oc8051_alu_src_sel1_n24,
         oc8051_alu_src_sel1_n23, oc8051_alu_src_sel1_n22,
         oc8051_alu_src_sel1_n21, oc8051_alu_src_sel1_n20,
         oc8051_alu_src_sel1_n19, oc8051_alu_src_sel1_n18,
         oc8051_alu_src_sel1_n17, oc8051_alu_src_sel1_n16,
         oc8051_alu_src_sel1_n15, oc8051_alu_src_sel1_n14,
         oc8051_alu_src_sel1_n13, oc8051_alu_src_sel1_n12,
         oc8051_alu_src_sel1_n11, oc8051_alu_src_sel1_n10,
         oc8051_alu_src_sel1_n9, oc8051_alu_src_sel1_n8,
         oc8051_alu_src_sel1_n7, oc8051_alu_src_sel1_n6,
         oc8051_alu_src_sel1_n5, oc8051_alu_src_sel1_n4,
         oc8051_alu_src_sel1_n3, oc8051_alu_src_sel1_n2,
         oc8051_alu_src_sel1_n1, oc8051_alu_src_sel1_n31,
         oc8051_alu_src_sel1_n30, oc8051_alu_src_sel1_n29,
         oc8051_alu_src_sel1_n25, oc8051_alu_src_sel1_op2_r_0_,
         oc8051_alu_src_sel1_op2_r_1_, oc8051_alu_src_sel1_op2_r_2_,
         oc8051_alu_src_sel1_op2_r_3_, oc8051_alu_src_sel1_op2_r_4_,
         oc8051_alu_src_sel1_op2_r_5_, oc8051_alu_src_sel1_op2_r_6_,
         oc8051_alu_src_sel1_op2_r_7_, oc8051_comp1_n10, oc8051_comp1_n9,
         oc8051_comp1_n8, oc8051_comp1_n7, oc8051_comp1_n6, oc8051_comp1_n5,
         oc8051_comp1_n4, oc8051_comp1_n3, oc8051_comp1_n2, oc8051_comp1_n1,
         oc8051_cy_select1_n1, oc8051_indi_addr1_n98, oc8051_indi_addr1_n97,
         oc8051_indi_addr1_n96, oc8051_indi_addr1_n95, oc8051_indi_addr1_n94,
         oc8051_indi_addr1_n93, oc8051_indi_addr1_n92, oc8051_indi_addr1_n27,
         oc8051_indi_addr1_n26, oc8051_indi_addr1_n25, oc8051_indi_addr1_n24,
         oc8051_indi_addr1_n23, oc8051_indi_addr1_n22, oc8051_indi_addr1_n21,
         oc8051_indi_addr1_n20, oc8051_indi_addr1_n19, oc8051_indi_addr1_n18,
         oc8051_indi_addr1_n17, oc8051_indi_addr1_n16, oc8051_indi_addr1_n15,
         oc8051_indi_addr1_n14, oc8051_indi_addr1_n13, oc8051_indi_addr1_n12,
         oc8051_indi_addr1_n11, oc8051_indi_addr1_n10, oc8051_indi_addr1_n9,
         oc8051_indi_addr1_n8, oc8051_indi_addr1_n7, oc8051_indi_addr1_n6,
         oc8051_indi_addr1_n5, oc8051_indi_addr1_n4, oc8051_indi_addr1_n3,
         oc8051_indi_addr1_n2, oc8051_indi_addr1_n1, oc8051_indi_addr1_n91,
         oc8051_indi_addr1_n90, oc8051_indi_addr1_n89, oc8051_indi_addr1_n88,
         oc8051_indi_addr1_n87, oc8051_indi_addr1_n86, oc8051_indi_addr1_n85,
         oc8051_indi_addr1_n84, oc8051_indi_addr1_n83, oc8051_indi_addr1_n82,
         oc8051_indi_addr1_n81, oc8051_indi_addr1_n80, oc8051_indi_addr1_n79,
         oc8051_indi_addr1_n78, oc8051_indi_addr1_n77, oc8051_indi_addr1_n76,
         oc8051_indi_addr1_n75, oc8051_indi_addr1_n74, oc8051_indi_addr1_n73,
         oc8051_indi_addr1_n72, oc8051_indi_addr1_n71, oc8051_indi_addr1_n70,
         oc8051_indi_addr1_n69, oc8051_indi_addr1_n68, oc8051_indi_addr1_n67,
         oc8051_indi_addr1_n66, oc8051_indi_addr1_n65, oc8051_indi_addr1_n64,
         oc8051_indi_addr1_n63, oc8051_indi_addr1_n62, oc8051_indi_addr1_n61,
         oc8051_indi_addr1_n60, oc8051_indi_addr1_n59, oc8051_indi_addr1_n58,
         oc8051_indi_addr1_n57, oc8051_indi_addr1_n56, oc8051_indi_addr1_n55,
         oc8051_indi_addr1_n54, oc8051_indi_addr1_n53, oc8051_indi_addr1_n52,
         oc8051_indi_addr1_n51, oc8051_indi_addr1_n50, oc8051_indi_addr1_n49,
         oc8051_indi_addr1_n48, oc8051_indi_addr1_n47, oc8051_indi_addr1_n46,
         oc8051_indi_addr1_n45, oc8051_indi_addr1_n44, oc8051_indi_addr1_n43,
         oc8051_indi_addr1_n42, oc8051_indi_addr1_n41, oc8051_indi_addr1_n40,
         oc8051_indi_addr1_n39, oc8051_indi_addr1_n38, oc8051_indi_addr1_n37,
         oc8051_indi_addr1_n36, oc8051_indi_addr1_n35, oc8051_indi_addr1_n34,
         oc8051_indi_addr1_n33, oc8051_indi_addr1_n32, oc8051_indi_addr1_n31,
         oc8051_indi_addr1_n30, oc8051_indi_addr1_n29, oc8051_indi_addr1_n28,
         oc8051_indi_addr1_n106, oc8051_indi_addr1_n105,
         oc8051_indi_addr1_n104, oc8051_indi_addr1_n103,
         oc8051_indi_addr1_n102, oc8051_indi_addr1_n101,
         oc8051_indi_addr1_n100, oc8051_indi_addr1_n99,
         oc8051_indi_addr1_wr_bit_r, oc8051_indi_addr1_buff_7__0_,
         oc8051_indi_addr1_buff_7__1_, oc8051_indi_addr1_buff_7__2_,
         oc8051_indi_addr1_buff_7__3_, oc8051_indi_addr1_buff_7__4_,
         oc8051_indi_addr1_buff_7__5_, oc8051_indi_addr1_buff_7__6_,
         oc8051_indi_addr1_buff_7__7_, oc8051_indi_addr1_buff_6__0_,
         oc8051_indi_addr1_buff_6__1_, oc8051_indi_addr1_buff_6__2_,
         oc8051_indi_addr1_buff_6__3_, oc8051_indi_addr1_buff_6__4_,
         oc8051_indi_addr1_buff_6__5_, oc8051_indi_addr1_buff_6__6_,
         oc8051_indi_addr1_buff_6__7_, oc8051_indi_addr1_buff_5__0_,
         oc8051_indi_addr1_buff_5__1_, oc8051_indi_addr1_buff_5__2_,
         oc8051_indi_addr1_buff_5__3_, oc8051_indi_addr1_buff_5__4_,
         oc8051_indi_addr1_buff_5__5_, oc8051_indi_addr1_buff_5__6_,
         oc8051_indi_addr1_buff_5__7_, oc8051_indi_addr1_buff_4__0_,
         oc8051_indi_addr1_buff_4__1_, oc8051_indi_addr1_buff_4__2_,
         oc8051_indi_addr1_buff_4__3_, oc8051_indi_addr1_buff_4__4_,
         oc8051_indi_addr1_buff_4__5_, oc8051_indi_addr1_buff_4__6_,
         oc8051_indi_addr1_buff_4__7_, oc8051_indi_addr1_buff_3__0_,
         oc8051_indi_addr1_buff_3__1_, oc8051_indi_addr1_buff_3__2_,
         oc8051_indi_addr1_buff_3__3_, oc8051_indi_addr1_buff_3__4_,
         oc8051_indi_addr1_buff_3__5_, oc8051_indi_addr1_buff_3__6_,
         oc8051_indi_addr1_buff_3__7_, oc8051_indi_addr1_buff_2__0_,
         oc8051_indi_addr1_buff_2__1_, oc8051_indi_addr1_buff_2__2_,
         oc8051_indi_addr1_buff_2__3_, oc8051_indi_addr1_buff_2__4_,
         oc8051_indi_addr1_buff_2__5_, oc8051_indi_addr1_buff_2__6_,
         oc8051_indi_addr1_buff_2__7_, oc8051_indi_addr1_buff_1__0_,
         oc8051_indi_addr1_buff_1__1_, oc8051_indi_addr1_buff_1__2_,
         oc8051_indi_addr1_buff_1__3_, oc8051_indi_addr1_buff_1__4_,
         oc8051_indi_addr1_buff_1__5_, oc8051_indi_addr1_buff_1__6_,
         oc8051_indi_addr1_buff_1__7_, oc8051_indi_addr1_buff_0__0_,
         oc8051_indi_addr1_buff_0__1_, oc8051_indi_addr1_buff_0__2_,
         oc8051_indi_addr1_buff_0__3_, oc8051_indi_addr1_buff_0__4_,
         oc8051_indi_addr1_buff_0__5_, oc8051_indi_addr1_buff_0__6_,
         oc8051_indi_addr1_buff_0__7_, oc8051_memory_interface1_n691,
         oc8051_memory_interface1_n682, oc8051_memory_interface1_n681,
         oc8051_memory_interface1_n680, oc8051_memory_interface1_n679,
         oc8051_memory_interface1_n678, oc8051_memory_interface1_n677,
         oc8051_memory_interface1_n676, oc8051_memory_interface1_n675,
         oc8051_memory_interface1_n674, oc8051_memory_interface1_n673,
         oc8051_memory_interface1_n672, oc8051_memory_interface1_n671,
         oc8051_memory_interface1_n670, oc8051_memory_interface1_n669,
         oc8051_memory_interface1_n668, oc8051_memory_interface1_n667,
         oc8051_memory_interface1_n666, oc8051_memory_interface1_n649,
         oc8051_memory_interface1_n648, oc8051_memory_interface1_n647,
         oc8051_memory_interface1_n646, oc8051_memory_interface1_n645,
         oc8051_memory_interface1_n644, oc8051_memory_interface1_n643,
         oc8051_memory_interface1_n642, oc8051_memory_interface1_n641,
         oc8051_memory_interface1_n640, oc8051_memory_interface1_n639,
         oc8051_memory_interface1_n638, oc8051_memory_interface1_n637,
         oc8051_memory_interface1_n636, oc8051_memory_interface1_n635,
         oc8051_memory_interface1_n634, oc8051_memory_interface1_n633,
         oc8051_memory_interface1_n632, oc8051_memory_interface1_n631,
         oc8051_memory_interface1_n630, oc8051_memory_interface1_n629,
         oc8051_memory_interface1_n628, oc8051_memory_interface1_n627,
         oc8051_memory_interface1_n626, oc8051_memory_interface1_n625,
         oc8051_memory_interface1_n624, oc8051_memory_interface1_n623,
         oc8051_memory_interface1_n622, oc8051_memory_interface1_n621,
         oc8051_memory_interface1_n620, oc8051_memory_interface1_n619,
         oc8051_memory_interface1_n618, oc8051_memory_interface1_n617,
         oc8051_memory_interface1_n616, oc8051_memory_interface1_n615,
         oc8051_memory_interface1_n614, oc8051_memory_interface1_n613,
         oc8051_memory_interface1_n612, oc8051_memory_interface1_n611,
         oc8051_memory_interface1_n610, oc8051_memory_interface1_n609,
         oc8051_memory_interface1_n608, oc8051_memory_interface1_n607,
         oc8051_memory_interface1_n606, oc8051_memory_interface1_n605,
         oc8051_memory_interface1_n604, oc8051_memory_interface1_n603,
         oc8051_memory_interface1_n602, oc8051_memory_interface1_n601,
         oc8051_memory_interface1_n600, oc8051_memory_interface1_n599,
         oc8051_memory_interface1_n598, oc8051_memory_interface1_n597,
         oc8051_memory_interface1_n596, oc8051_memory_interface1_n595,
         oc8051_memory_interface1_n594, oc8051_memory_interface1_n593,
         oc8051_memory_interface1_n592, oc8051_memory_interface1_n591,
         oc8051_memory_interface1_n590, oc8051_memory_interface1_n589,
         oc8051_memory_interface1_n588, oc8051_memory_interface1_n587,
         oc8051_memory_interface1_n586, oc8051_memory_interface1_n585,
         oc8051_memory_interface1_n584, oc8051_memory_interface1_n583,
         oc8051_memory_interface1_n582, oc8051_memory_interface1_n581,
         oc8051_memory_interface1_n580, oc8051_memory_interface1_n579,
         oc8051_memory_interface1_n578, oc8051_memory_interface1_n577,
         oc8051_memory_interface1_n576, oc8051_memory_interface1_n575,
         oc8051_memory_interface1_n574, oc8051_memory_interface1_n573,
         oc8051_memory_interface1_n572, oc8051_memory_interface1_n571,
         oc8051_memory_interface1_n570, oc8051_memory_interface1_n541,
         oc8051_memory_interface1_n539, oc8051_memory_interface1_n537,
         oc8051_memory_interface1_n535, oc8051_memory_interface1_n533,
         oc8051_memory_interface1_n531, oc8051_memory_interface1_n529,
         oc8051_memory_interface1_n527, oc8051_memory_interface1_n443,
         oc8051_memory_interface1_n442, oc8051_memory_interface1_n441,
         oc8051_memory_interface1_n424, oc8051_memory_interface1_n423,
         oc8051_memory_interface1_n422, oc8051_memory_interface1_n421,
         oc8051_memory_interface1_n420, oc8051_memory_interface1_n419,
         oc8051_memory_interface1_n418, oc8051_memory_interface1_n417,
         oc8051_memory_interface1_n400, oc8051_memory_interface1_n399,
         oc8051_memory_interface1_n398, oc8051_memory_interface1_n397,
         oc8051_memory_interface1_n396, oc8051_memory_interface1_n395,
         oc8051_memory_interface1_n394, oc8051_memory_interface1_n393,
         oc8051_memory_interface1_n392, oc8051_memory_interface1_n391,
         oc8051_memory_interface1_n390, oc8051_memory_interface1_n389,
         oc8051_memory_interface1_n388, oc8051_memory_interface1_n387,
         oc8051_memory_interface1_n386, oc8051_memory_interface1_n385,
         oc8051_memory_interface1_n376, oc8051_memory_interface1_n375,
         oc8051_memory_interface1_n374, oc8051_memory_interface1_n373,
         oc8051_memory_interface1_n372, oc8051_memory_interface1_n371,
         oc8051_memory_interface1_n370, oc8051_memory_interface1_n369,
         oc8051_memory_interface1_n368, oc8051_memory_interface1_n367,
         oc8051_memory_interface1_n366, oc8051_memory_interface1_n365,
         oc8051_memory_interface1_n364, oc8051_memory_interface1_n363,
         oc8051_memory_interface1_n362, oc8051_memory_interface1_n361,
         oc8051_memory_interface1_n360, oc8051_memory_interface1_n359,
         oc8051_memory_interface1_n358, oc8051_memory_interface1_n357,
         oc8051_memory_interface1_n356, oc8051_memory_interface1_n355,
         oc8051_memory_interface1_n354, oc8051_memory_interface1_n353,
         oc8051_memory_interface1_n352, oc8051_memory_interface1_n351,
         oc8051_memory_interface1_n350, oc8051_memory_interface1_n349,
         oc8051_memory_interface1_n348, oc8051_memory_interface1_n347,
         oc8051_memory_interface1_n346, oc8051_memory_interface1_n345,
         oc8051_memory_interface1_n344, oc8051_memory_interface1_n343,
         oc8051_memory_interface1_n342, oc8051_memory_interface1_n341,
         oc8051_memory_interface1_n340, oc8051_memory_interface1_n339,
         oc8051_memory_interface1_n338, oc8051_memory_interface1_n337,
         oc8051_memory_interface1_n336, oc8051_memory_interface1_n335,
         oc8051_memory_interface1_n334, oc8051_memory_interface1_n333,
         oc8051_memory_interface1_n332, oc8051_memory_interface1_n331,
         oc8051_memory_interface1_n330, oc8051_memory_interface1_n329,
         oc8051_memory_interface1_n328, oc8051_memory_interface1_n327,
         oc8051_memory_interface1_n326, oc8051_memory_interface1_n325,
         oc8051_memory_interface1_n324, oc8051_memory_interface1_n323,
         oc8051_memory_interface1_n321, oc8051_memory_interface1_n320,
         oc8051_memory_interface1_n319, oc8051_memory_interface1_n318,
         oc8051_memory_interface1_n317, oc8051_memory_interface1_n316,
         oc8051_memory_interface1_n315, oc8051_memory_interface1_n314,
         oc8051_memory_interface1_n313, oc8051_memory_interface1_n312,
         oc8051_memory_interface1_n311, oc8051_memory_interface1_n310,
         oc8051_memory_interface1_n309, oc8051_memory_interface1_n308,
         oc8051_memory_interface1_n307, oc8051_memory_interface1_n306,
         oc8051_memory_interface1_n305, oc8051_memory_interface1_n304,
         oc8051_memory_interface1_n303, oc8051_memory_interface1_n302,
         oc8051_memory_interface1_n301, oc8051_memory_interface1_n300,
         oc8051_memory_interface1_n299, oc8051_memory_interface1_n298,
         oc8051_memory_interface1_n297, oc8051_memory_interface1_n296,
         oc8051_memory_interface1_n295, oc8051_memory_interface1_n294,
         oc8051_memory_interface1_n293, oc8051_memory_interface1_n292,
         oc8051_memory_interface1_n291, oc8051_memory_interface1_n290,
         oc8051_memory_interface1_n289, oc8051_memory_interface1_n288,
         oc8051_memory_interface1_n287, oc8051_memory_interface1_n286,
         oc8051_memory_interface1_n285, oc8051_memory_interface1_n284,
         oc8051_memory_interface1_n283, oc8051_memory_interface1_n282,
         oc8051_memory_interface1_n281, oc8051_memory_interface1_n280,
         oc8051_memory_interface1_n279, oc8051_memory_interface1_n278,
         oc8051_memory_interface1_n277, oc8051_memory_interface1_n276,
         oc8051_memory_interface1_n275, oc8051_memory_interface1_n274,
         oc8051_memory_interface1_n273, oc8051_memory_interface1_n272,
         oc8051_memory_interface1_n271, oc8051_memory_interface1_n270,
         oc8051_memory_interface1_n269, oc8051_memory_interface1_n268,
         oc8051_memory_interface1_n267, oc8051_memory_interface1_n266,
         oc8051_memory_interface1_n265, oc8051_memory_interface1_n264,
         oc8051_memory_interface1_n263, oc8051_memory_interface1_n262,
         oc8051_memory_interface1_n261, oc8051_memory_interface1_n260,
         oc8051_memory_interface1_n259, oc8051_memory_interface1_n258,
         oc8051_memory_interface1_n257, oc8051_memory_interface1_n256,
         oc8051_memory_interface1_n255, oc8051_memory_interface1_n254,
         oc8051_memory_interface1_n253, oc8051_memory_interface1_n252,
         oc8051_memory_interface1_n251, oc8051_memory_interface1_n250,
         oc8051_memory_interface1_n249, oc8051_memory_interface1_n248,
         oc8051_memory_interface1_n247, oc8051_memory_interface1_n246,
         oc8051_memory_interface1_n245, oc8051_memory_interface1_n244,
         oc8051_memory_interface1_n243, oc8051_memory_interface1_n242,
         oc8051_memory_interface1_n241, oc8051_memory_interface1_n240,
         oc8051_memory_interface1_n239, oc8051_memory_interface1_n238,
         oc8051_memory_interface1_n237, oc8051_memory_interface1_n236,
         oc8051_memory_interface1_n235, oc8051_memory_interface1_n234,
         oc8051_memory_interface1_n233, oc8051_memory_interface1_n232,
         oc8051_memory_interface1_n231, oc8051_memory_interface1_n230,
         oc8051_memory_interface1_n229, oc8051_memory_interface1_n228,
         oc8051_memory_interface1_n227, oc8051_memory_interface1_n226,
         oc8051_memory_interface1_n225, oc8051_memory_interface1_n224,
         oc8051_memory_interface1_n223, oc8051_memory_interface1_n222,
         oc8051_memory_interface1_n221, oc8051_memory_interface1_n220,
         oc8051_memory_interface1_n219, oc8051_memory_interface1_n218,
         oc8051_memory_interface1_n217, oc8051_memory_interface1_n216,
         oc8051_memory_interface1_n215, oc8051_memory_interface1_n214,
         oc8051_memory_interface1_n213, oc8051_memory_interface1_n212,
         oc8051_memory_interface1_n211, oc8051_memory_interface1_n210,
         oc8051_memory_interface1_n209, oc8051_memory_interface1_n208,
         oc8051_memory_interface1_n207, oc8051_memory_interface1_n206,
         oc8051_memory_interface1_n205, oc8051_memory_interface1_n204,
         oc8051_memory_interface1_n203, oc8051_memory_interface1_n202,
         oc8051_memory_interface1_n201, oc8051_memory_interface1_n200,
         oc8051_memory_interface1_n199, oc8051_memory_interface1_n198,
         oc8051_memory_interface1_n197, oc8051_memory_interface1_n196,
         oc8051_memory_interface1_n195, oc8051_memory_interface1_n194,
         oc8051_memory_interface1_n193, oc8051_memory_interface1_n192,
         oc8051_memory_interface1_n191, oc8051_memory_interface1_n190,
         oc8051_memory_interface1_n189, oc8051_memory_interface1_n188,
         oc8051_memory_interface1_n187, oc8051_memory_interface1_n186,
         oc8051_memory_interface1_n185, oc8051_memory_interface1_n184,
         oc8051_memory_interface1_n183, oc8051_memory_interface1_n182,
         oc8051_memory_interface1_n181, oc8051_memory_interface1_n180,
         oc8051_memory_interface1_n179, oc8051_memory_interface1_n178,
         oc8051_memory_interface1_n177, oc8051_memory_interface1_n176,
         oc8051_memory_interface1_n175, oc8051_memory_interface1_n174,
         oc8051_memory_interface1_n173, oc8051_memory_interface1_n172,
         oc8051_memory_interface1_n171, oc8051_memory_interface1_n170,
         oc8051_memory_interface1_n169, oc8051_memory_interface1_n168,
         oc8051_memory_interface1_n167, oc8051_memory_interface1_n166,
         oc8051_memory_interface1_n165, oc8051_memory_interface1_n164,
         oc8051_memory_interface1_n163, oc8051_memory_interface1_n162,
         oc8051_memory_interface1_n161, oc8051_memory_interface1_n160,
         oc8051_memory_interface1_n159, oc8051_memory_interface1_n158,
         oc8051_memory_interface1_n157, oc8051_memory_interface1_n156,
         oc8051_memory_interface1_n155, oc8051_memory_interface1_n154,
         oc8051_memory_interface1_n153, oc8051_memory_interface1_n152,
         oc8051_memory_interface1_n151, oc8051_memory_interface1_n150,
         oc8051_memory_interface1_n149, oc8051_memory_interface1_n148,
         oc8051_memory_interface1_n147, oc8051_memory_interface1_n146,
         oc8051_memory_interface1_n145, oc8051_memory_interface1_n144,
         oc8051_memory_interface1_n143, oc8051_memory_interface1_n142,
         oc8051_memory_interface1_n141, oc8051_memory_interface1_n140,
         oc8051_memory_interface1_n139, oc8051_memory_interface1_n138,
         oc8051_memory_interface1_n137, oc8051_memory_interface1_n136,
         oc8051_memory_interface1_n135, oc8051_memory_interface1_n134,
         oc8051_memory_interface1_n133, oc8051_memory_interface1_n132,
         oc8051_memory_interface1_n131, oc8051_memory_interface1_n130,
         oc8051_memory_interface1_n129, oc8051_memory_interface1_n128,
         oc8051_memory_interface1_n127, oc8051_memory_interface1_n126,
         oc8051_memory_interface1_n125, oc8051_memory_interface1_n124,
         oc8051_memory_interface1_n123, oc8051_memory_interface1_n122,
         oc8051_memory_interface1_n121, oc8051_memory_interface1_n120,
         oc8051_memory_interface1_n119, oc8051_memory_interface1_n118,
         oc8051_memory_interface1_n117, oc8051_memory_interface1_n116,
         oc8051_memory_interface1_n115, oc8051_memory_interface1_n114,
         oc8051_memory_interface1_n113, oc8051_memory_interface1_n112,
         oc8051_memory_interface1_n111, oc8051_memory_interface1_n110,
         oc8051_memory_interface1_n109, oc8051_memory_interface1_n108,
         oc8051_memory_interface1_n107, oc8051_memory_interface1_n106,
         oc8051_memory_interface1_n105, oc8051_memory_interface1_n104,
         oc8051_memory_interface1_n103, oc8051_memory_interface1_n102,
         oc8051_memory_interface1_n101, oc8051_memory_interface1_n100,
         oc8051_memory_interface1_n99, oc8051_memory_interface1_n98,
         oc8051_memory_interface1_n97, oc8051_memory_interface1_n96,
         oc8051_memory_interface1_n95, oc8051_memory_interface1_n94,
         oc8051_memory_interface1_n93, oc8051_memory_interface1_n92,
         oc8051_memory_interface1_n91, oc8051_memory_interface1_n90,
         oc8051_memory_interface1_n89, oc8051_memory_interface1_n88,
         oc8051_memory_interface1_n87, oc8051_memory_interface1_n86,
         oc8051_memory_interface1_n85, oc8051_memory_interface1_n84,
         oc8051_memory_interface1_n83, oc8051_memory_interface1_n82,
         oc8051_memory_interface1_n81, oc8051_memory_interface1_n80,
         oc8051_memory_interface1_n79, oc8051_memory_interface1_n78,
         oc8051_memory_interface1_n77, oc8051_memory_interface1_n76,
         oc8051_memory_interface1_n75, oc8051_memory_interface1_n74,
         oc8051_memory_interface1_n73, oc8051_memory_interface1_n72,
         oc8051_memory_interface1_n71, oc8051_memory_interface1_n70,
         oc8051_memory_interface1_n69, oc8051_memory_interface1_n68,
         oc8051_memory_interface1_n67, oc8051_memory_interface1_n66,
         oc8051_memory_interface1_n65, oc8051_memory_interface1_n64,
         oc8051_memory_interface1_n63, oc8051_memory_interface1_n62,
         oc8051_memory_interface1_n61, oc8051_memory_interface1_n60,
         oc8051_memory_interface1_n59, oc8051_memory_interface1_n58,
         oc8051_memory_interface1_n57, oc8051_memory_interface1_n56,
         oc8051_memory_interface1_n55, oc8051_memory_interface1_n54,
         oc8051_memory_interface1_n53, oc8051_memory_interface1_n52,
         oc8051_memory_interface1_n51, oc8051_memory_interface1_n50,
         oc8051_memory_interface1_n49, oc8051_memory_interface1_n48,
         oc8051_memory_interface1_n47, oc8051_memory_interface1_n46,
         oc8051_memory_interface1_n45, oc8051_memory_interface1_n44,
         oc8051_memory_interface1_n43, oc8051_memory_interface1_n42,
         oc8051_memory_interface1_n41, oc8051_memory_interface1_n40,
         oc8051_memory_interface1_n39, oc8051_memory_interface1_n38,
         oc8051_memory_interface1_n37, oc8051_memory_interface1_n36,
         oc8051_memory_interface1_n35, oc8051_memory_interface1_n34,
         oc8051_memory_interface1_n33, oc8051_memory_interface1_n32,
         oc8051_memory_interface1_n31, oc8051_memory_interface1_n30,
         oc8051_memory_interface1_n29, oc8051_memory_interface1_n28,
         oc8051_memory_interface1_n27, oc8051_memory_interface1_n26,
         oc8051_memory_interface1_n25, oc8051_memory_interface1_n24,
         oc8051_memory_interface1_n23, oc8051_memory_interface1_n22,
         oc8051_memory_interface1_n21, oc8051_memory_interface1_n20,
         oc8051_memory_interface1_n19, oc8051_memory_interface1_n18,
         oc8051_memory_interface1_n17, oc8051_memory_interface1_n16,
         oc8051_memory_interface1_n15, oc8051_memory_interface1_n14,
         oc8051_memory_interface1_n13, oc8051_memory_interface1_n12,
         oc8051_memory_interface1_n11, oc8051_memory_interface1_n10,
         oc8051_memory_interface1_n9, oc8051_memory_interface1_n8,
         oc8051_memory_interface1_n7, oc8051_memory_interface1_n6,
         oc8051_memory_interface1_n5, oc8051_memory_interface1_n4,
         oc8051_memory_interface1_n3, oc8051_memory_interface1_n2,
         oc8051_memory_interface1_n1, oc8051_memory_interface1_r390_carry_8_,
         oc8051_memory_interface1_r390_carry_7_,
         oc8051_memory_interface1_r390_carry_6_,
         oc8051_memory_interface1_r390_carry_5_,
         oc8051_memory_interface1_r390_carry_4_,
         oc8051_memory_interface1_r390_carry_3_,
         oc8051_memory_interface1_r390_carry_2_,
         oc8051_memory_interface1_add_2_root_add_937_2_carry_3_,
         oc8051_memory_interface1_add_2_root_add_937_2_carry_2_,
         oc8051_memory_interface1_add_0_root_add_937_2_carry_2_,
         oc8051_memory_interface1_n569, oc8051_memory_interface1_n568,
         oc8051_memory_interface1_n567, oc8051_memory_interface1_n566,
         oc8051_memory_interface1_n565, oc8051_memory_interface1_n564,
         oc8051_memory_interface1_n563, oc8051_memory_interface1_n562,
         oc8051_memory_interface1_n561, oc8051_memory_interface1_n560,
         oc8051_memory_interface1_n559, oc8051_memory_interface1_n558,
         oc8051_memory_interface1_n557, oc8051_memory_interface1_n556,
         oc8051_memory_interface1_n555, oc8051_memory_interface1_n554,
         oc8051_memory_interface1_n553, oc8051_memory_interface1_n552,
         oc8051_memory_interface1_n551, oc8051_memory_interface1_n550,
         oc8051_memory_interface1_n549, oc8051_memory_interface1_n548,
         oc8051_memory_interface1_n547, oc8051_memory_interface1_n546,
         oc8051_memory_interface1_n545, oc8051_memory_interface1_n544,
         oc8051_memory_interface1_n543, oc8051_memory_interface1_n542,
         oc8051_memory_interface1_n540, oc8051_memory_interface1_n538,
         oc8051_memory_interface1_n536, oc8051_memory_interface1_n534,
         oc8051_memory_interface1_n532, oc8051_memory_interface1_n530,
         oc8051_memory_interface1_n528, oc8051_memory_interface1_n526,
         oc8051_memory_interface1_n525, oc8051_memory_interface1_n524,
         oc8051_memory_interface1_n523, oc8051_memory_interface1_n522,
         oc8051_memory_interface1_n521, oc8051_memory_interface1_n520,
         oc8051_memory_interface1_n519, oc8051_memory_interface1_n518,
         oc8051_memory_interface1_n517, oc8051_memory_interface1_n516,
         oc8051_memory_interface1_n515, oc8051_memory_interface1_n514,
         oc8051_memory_interface1_n513, oc8051_memory_interface1_n512,
         oc8051_memory_interface1_n511, oc8051_memory_interface1_n510,
         oc8051_memory_interface1_n509, oc8051_memory_interface1_n508,
         oc8051_memory_interface1_n507, oc8051_memory_interface1_n506,
         oc8051_memory_interface1_n505, oc8051_memory_interface1_n504,
         oc8051_memory_interface1_n503, oc8051_memory_interface1_n502,
         oc8051_memory_interface1_n501, oc8051_memory_interface1_n500,
         oc8051_memory_interface1_n499, oc8051_memory_interface1_n498,
         oc8051_memory_interface1_n497, oc8051_memory_interface1_n496,
         oc8051_memory_interface1_n495, oc8051_memory_interface1_n494,
         oc8051_memory_interface1_n493, oc8051_memory_interface1_n492,
         oc8051_memory_interface1_n491, oc8051_memory_interface1_n490,
         oc8051_memory_interface1_n489, oc8051_memory_interface1_n488,
         oc8051_memory_interface1_n487, oc8051_memory_interface1_n486,
         oc8051_memory_interface1_n485, oc8051_memory_interface1_n484,
         oc8051_memory_interface1_n483, oc8051_memory_interface1_n482,
         oc8051_memory_interface1_n481, oc8051_memory_interface1_n480,
         oc8051_memory_interface1_n479, oc8051_memory_interface1_n478,
         oc8051_memory_interface1_n477, oc8051_memory_interface1_n476,
         oc8051_memory_interface1_n475, oc8051_memory_interface1_n474,
         oc8051_memory_interface1_n473, oc8051_memory_interface1_n472,
         oc8051_memory_interface1_n471, oc8051_memory_interface1_n470,
         oc8051_memory_interface1_n469, oc8051_memory_interface1_n468,
         oc8051_memory_interface1_n467, oc8051_memory_interface1_n466,
         oc8051_memory_interface1_n465, oc8051_memory_interface1_n464,
         oc8051_memory_interface1_n463, oc8051_memory_interface1_n462,
         oc8051_memory_interface1_n461, oc8051_memory_interface1_n460,
         oc8051_memory_interface1_n459, oc8051_memory_interface1_n458,
         oc8051_memory_interface1_n457, oc8051_memory_interface1_n456,
         oc8051_memory_interface1_n455, oc8051_memory_interface1_n454,
         oc8051_memory_interface1_n453, oc8051_memory_interface1_n452,
         oc8051_memory_interface1_n451, oc8051_memory_interface1_n450,
         oc8051_memory_interface1_n449, oc8051_memory_interface1_n448,
         oc8051_memory_interface1_n447, oc8051_memory_interface1_n446,
         oc8051_memory_interface1_n445, oc8051_memory_interface1_n444,
         oc8051_memory_interface1_n440, oc8051_memory_interface1_n439,
         oc8051_memory_interface1_n438, oc8051_memory_interface1_n437,
         oc8051_memory_interface1_n436, oc8051_memory_interface1_n435,
         oc8051_memory_interface1_n434, oc8051_memory_interface1_n433,
         oc8051_memory_interface1_n432, oc8051_memory_interface1_n431,
         oc8051_memory_interface1_n430, oc8051_memory_interface1_n429,
         oc8051_memory_interface1_n428, oc8051_memory_interface1_n427,
         oc8051_memory_interface1_n426, oc8051_memory_interface1_n425,
         oc8051_memory_interface1_n416, oc8051_memory_interface1_n415,
         oc8051_memory_interface1_n414, oc8051_memory_interface1_n413,
         oc8051_memory_interface1_n412, oc8051_memory_interface1_n411,
         oc8051_memory_interface1_n410, oc8051_memory_interface1_n409,
         oc8051_memory_interface1_n408, oc8051_memory_interface1_n407,
         oc8051_memory_interface1_n406, oc8051_memory_interface1_n405,
         oc8051_memory_interface1_n404, oc8051_memory_interface1_n403,
         oc8051_memory_interface1_n402, oc8051_memory_interface1_n401,
         oc8051_memory_interface1_n384, oc8051_memory_interface1_n383,
         oc8051_memory_interface1_n382, oc8051_memory_interface1_n381,
         oc8051_memory_interface1_n380, oc8051_memory_interface1_n379,
         oc8051_memory_interface1_n378, oc8051_memory_interface1_n377,
         oc8051_memory_interface1_n322, oc8051_memory_interface1_u3_u7_z_15,
         oc8051_memory_interface1_u3_u7_z_14,
         oc8051_memory_interface1_u3_u7_z_13,
         oc8051_memory_interface1_u3_u7_z_12,
         oc8051_memory_interface1_u3_u7_z_11,
         oc8051_memory_interface1_u3_u7_z_10,
         oc8051_memory_interface1_u3_u7_z_9,
         oc8051_memory_interface1_u3_u7_z_8, oc8051_memory_interface1_n5360,
         oc8051_memory_interface1_pc_wr_r, oc8051_memory_interface1_n4560,
         oc8051_memory_interface1_n4550, oc8051_memory_interface1_n4540,
         oc8051_memory_interface1_n4530, oc8051_memory_interface1_n4520,
         oc8051_memory_interface1_n4510, oc8051_memory_interface1_n4500,
         oc8051_memory_interface1_n4490, oc8051_memory_interface1_n4480,
         oc8051_memory_interface1_n4470, oc8051_memory_interface1_n4460,
         oc8051_memory_interface1_n4450, oc8051_memory_interface1_n4440,
         oc8051_memory_interface1_n4430, oc8051_memory_interface1_n4420,
         oc8051_memory_interface1_n4410, oc8051_memory_interface1_n4260,
         oc8051_memory_interface1_n4250, oc8051_memory_interface1_n4240,
         oc8051_memory_interface1_n4230, oc8051_memory_interface1_n4220,
         oc8051_memory_interface1_n4210, oc8051_memory_interface1_n4200,
         oc8051_memory_interface1_n4190, oc8051_memory_interface1_n4180,
         oc8051_memory_interface1_n4170, oc8051_memory_interface1_n4160,
         oc8051_memory_interface1_n4150, oc8051_memory_interface1_n4140,
         oc8051_memory_interface1_n4130, oc8051_memory_interface1_n4120,
         oc8051_memory_interface1_n4110, oc8051_memory_interface1_n4100,
         oc8051_memory_interface1_n4090, oc8051_memory_interface1_pc_buf_0_,
         oc8051_memory_interface1_pc_buf_1_,
         oc8051_memory_interface1_pc_buf_2_,
         oc8051_memory_interface1_pc_buf_3_,
         oc8051_memory_interface1_pc_buf_4_,
         oc8051_memory_interface1_pc_buf_5_,
         oc8051_memory_interface1_pc_buf_6_,
         oc8051_memory_interface1_pc_buf_7_,
         oc8051_memory_interface1_pc_buf_8_,
         oc8051_memory_interface1_pc_buf_9_,
         oc8051_memory_interface1_pc_buf_10_,
         oc8051_memory_interface1_pc_buf_11_,
         oc8051_memory_interface1_pc_buf_12_,
         oc8051_memory_interface1_pc_buf_13_,
         oc8051_memory_interface1_pc_buf_14_,
         oc8051_memory_interface1_pc_buf_15_, oc8051_memory_interface1_n4060,
         oc8051_memory_interface1_n4050, oc8051_memory_interface1_n4040,
         oc8051_memory_interface1_n4030, oc8051_memory_interface1_n4020,
         oc8051_memory_interface1_n4010, oc8051_memory_interface1_n4000,
         oc8051_memory_interface1_n3990, oc8051_memory_interface1_n3900,
         oc8051_memory_interface1_n3890, oc8051_memory_interface1_n3880,
         oc8051_memory_interface1_n3870, oc8051_memory_interface1_n3860,
         oc8051_memory_interface1_n3850, oc8051_memory_interface1_n3840,
         oc8051_memory_interface1_n3830,
         oc8051_memory_interface1_pcs_source_0_,
         oc8051_memory_interface1_pcs_source_1_,
         oc8051_memory_interface1_pcs_source_2_,
         oc8051_memory_interface1_pcs_source_3_,
         oc8051_memory_interface1_pcs_source_4_,
         oc8051_memory_interface1_pcs_source_5_,
         oc8051_memory_interface1_pcs_source_6_,
         oc8051_memory_interface1_pcs_source_7_,
         oc8051_memory_interface1_n3700, oc8051_memory_interface1_int_ack_buff,
         oc8051_memory_interface1_n1980,
         oc8051_memory_interface1_int_vec_buff_0_,
         oc8051_memory_interface1_int_vec_buff_1_,
         oc8051_memory_interface1_int_vec_buff_2_,
         oc8051_memory_interface1_int_vec_buff_3_,
         oc8051_memory_interface1_int_vec_buff_4_,
         oc8051_memory_interface1_int_vec_buff_5_,
         oc8051_memory_interface1_int_vec_buff_6_,
         oc8051_memory_interface1_int_vec_buff_7_,
         oc8051_memory_interface1_int_ack_t,
         oc8051_memory_interface1_ddat_ir_0_,
         oc8051_memory_interface1_ddat_ir_1_,
         oc8051_memory_interface1_ddat_ir_2_,
         oc8051_memory_interface1_ddat_ir_3_,
         oc8051_memory_interface1_ddat_ir_4_,
         oc8051_memory_interface1_ddat_ir_5_,
         oc8051_memory_interface1_ddat_ir_6_,
         oc8051_memory_interface1_ddat_ir_7_, oc8051_memory_interface1_dack_ir,
         oc8051_memory_interface1_op1_0_, oc8051_memory_interface1_op1_1_,
         oc8051_memory_interface1_op1_2_, oc8051_memory_interface1_op1_3_,
         oc8051_memory_interface1_op1_4_, oc8051_memory_interface1_op1_5_,
         oc8051_memory_interface1_op1_6_, oc8051_memory_interface1_op1_7_,
         oc8051_memory_interface1_op_pos_0_,
         oc8051_memory_interface1_op_pos_1_,
         oc8051_memory_interface1_op_pos_2_, oc8051_memory_interface1_cdone,
         oc8051_memory_interface1_cdata_0_, oc8051_memory_interface1_cdata_1_,
         oc8051_memory_interface1_cdata_2_, oc8051_memory_interface1_cdata_3_,
         oc8051_memory_interface1_cdata_4_, oc8051_memory_interface1_cdata_5_,
         oc8051_memory_interface1_cdata_6_, oc8051_memory_interface1_cdata_7_,
         oc8051_memory_interface1_inc_pc, oc8051_memory_interface1_idat_cur_0_,
         oc8051_memory_interface1_idat_cur_1_,
         oc8051_memory_interface1_idat_cur_2_,
         oc8051_memory_interface1_idat_cur_3_,
         oc8051_memory_interface1_idat_cur_4_,
         oc8051_memory_interface1_idat_cur_5_,
         oc8051_memory_interface1_idat_cur_6_,
         oc8051_memory_interface1_idat_cur_7_,
         oc8051_memory_interface1_idat_cur_8_,
         oc8051_memory_interface1_idat_cur_9_,
         oc8051_memory_interface1_idat_cur_10_,
         oc8051_memory_interface1_idat_cur_11_,
         oc8051_memory_interface1_idat_cur_12_,
         oc8051_memory_interface1_idat_cur_13_,
         oc8051_memory_interface1_idat_cur_14_,
         oc8051_memory_interface1_idat_cur_15_,
         oc8051_memory_interface1_idat_cur_16_,
         oc8051_memory_interface1_idat_cur_17_,
         oc8051_memory_interface1_idat_cur_18_,
         oc8051_memory_interface1_idat_cur_19_,
         oc8051_memory_interface1_idat_cur_20_,
         oc8051_memory_interface1_idat_cur_21_,
         oc8051_memory_interface1_idat_cur_22_,
         oc8051_memory_interface1_idat_cur_23_,
         oc8051_memory_interface1_idat_cur_24_,
         oc8051_memory_interface1_idat_cur_25_,
         oc8051_memory_interface1_idat_cur_26_,
         oc8051_memory_interface1_idat_cur_27_,
         oc8051_memory_interface1_idat_cur_28_,
         oc8051_memory_interface1_idat_cur_29_,
         oc8051_memory_interface1_idat_cur_30_,
         oc8051_memory_interface1_idat_cur_31_,
         oc8051_memory_interface1_idat_old_0_,
         oc8051_memory_interface1_idat_old_1_,
         oc8051_memory_interface1_idat_old_2_,
         oc8051_memory_interface1_idat_old_3_,
         oc8051_memory_interface1_idat_old_4_,
         oc8051_memory_interface1_idat_old_5_,
         oc8051_memory_interface1_idat_old_6_,
         oc8051_memory_interface1_idat_old_7_,
         oc8051_memory_interface1_idat_old_8_,
         oc8051_memory_interface1_idat_old_9_,
         oc8051_memory_interface1_idat_old_10_,
         oc8051_memory_interface1_idat_old_11_,
         oc8051_memory_interface1_idat_old_12_,
         oc8051_memory_interface1_idat_old_13_,
         oc8051_memory_interface1_idat_old_14_,
         oc8051_memory_interface1_idat_old_15_,
         oc8051_memory_interface1_idat_old_16_,
         oc8051_memory_interface1_idat_old_17_,
         oc8051_memory_interface1_idat_old_18_,
         oc8051_memory_interface1_idat_old_19_,
         oc8051_memory_interface1_idat_old_20_,
         oc8051_memory_interface1_idat_old_21_,
         oc8051_memory_interface1_idat_old_22_,
         oc8051_memory_interface1_idat_old_23_,
         oc8051_memory_interface1_idat_old_24_,
         oc8051_memory_interface1_idat_old_25_,
         oc8051_memory_interface1_idat_old_26_,
         oc8051_memory_interface1_idat_old_27_,
         oc8051_memory_interface1_idat_old_28_,
         oc8051_memory_interface1_idat_old_29_,
         oc8051_memory_interface1_idat_old_30_,
         oc8051_memory_interface1_idat_old_31_, oc8051_memory_interface1_n1290,
         oc8051_memory_interface1_pc_out_7_,
         oc8051_memory_interface1_pc_out_15_,
         oc8051_memory_interface1_iadr_t_0_,
         oc8051_memory_interface1_iadr_t_1_,
         oc8051_memory_interface1_iadr_t_2_,
         oc8051_memory_interface1_iadr_t_3_,
         oc8051_memory_interface1_iadr_t_4_,
         oc8051_memory_interface1_iadr_t_5_,
         oc8051_memory_interface1_iadr_t_6_,
         oc8051_memory_interface1_iadr_t_7_,
         oc8051_memory_interface1_iadr_t_8_,
         oc8051_memory_interface1_iadr_t_9_,
         oc8051_memory_interface1_iadr_t_10_,
         oc8051_memory_interface1_iadr_t_11_,
         oc8051_memory_interface1_iadr_t_12_,
         oc8051_memory_interface1_iadr_t_13_,
         oc8051_memory_interface1_iadr_t_14_,
         oc8051_memory_interface1_iadr_t_15_, oc8051_memory_interface1_n810,
         oc8051_memory_interface1_rd_addr_r, oc8051_memory_interface1_istb_t,
         oc8051_memory_interface1_pc_wr_r2, oc8051_memory_interface1_imem_wait,
         oc8051_memory_interface1_dmem_wait, oc8051_memory_interface1_istb_o,
         oc8051_memory_interface1_rd_ind, oc8051_sfr1_n259, oc8051_sfr1_n258,
         oc8051_sfr1_n257, oc8051_sfr1_n256, oc8051_sfr1_n255,
         oc8051_sfr1_n254, oc8051_sfr1_n253, oc8051_sfr1_n252,
         oc8051_sfr1_n251, oc8051_sfr1_n250, oc8051_sfr1_n249,
         oc8051_sfr1_n248, oc8051_sfr1_n247, oc8051_sfr1_n246,
         oc8051_sfr1_n245, oc8051_sfr1_n236, oc8051_sfr1_n235,
         oc8051_sfr1_n234, oc8051_sfr1_n233, oc8051_sfr1_n232,
         oc8051_sfr1_n231, oc8051_sfr1_n230, oc8051_sfr1_n229,
         oc8051_sfr1_n228, oc8051_sfr1_n227, oc8051_sfr1_n226,
         oc8051_sfr1_n225, oc8051_sfr1_n224, oc8051_sfr1_n223,
         oc8051_sfr1_n222, oc8051_sfr1_n221, oc8051_sfr1_n220,
         oc8051_sfr1_n219, oc8051_sfr1_n218, oc8051_sfr1_n217,
         oc8051_sfr1_n216, oc8051_sfr1_n215, oc8051_sfr1_n214,
         oc8051_sfr1_n213, oc8051_sfr1_n212, oc8051_sfr1_n211,
         oc8051_sfr1_n210, oc8051_sfr1_n209, oc8051_sfr1_n208,
         oc8051_sfr1_n207, oc8051_sfr1_n206, oc8051_sfr1_n205,
         oc8051_sfr1_n204, oc8051_sfr1_n203, oc8051_sfr1_n202,
         oc8051_sfr1_n201, oc8051_sfr1_n200, oc8051_sfr1_n199,
         oc8051_sfr1_n198, oc8051_sfr1_n197, oc8051_sfr1_n196,
         oc8051_sfr1_n195, oc8051_sfr1_n194, oc8051_sfr1_n193,
         oc8051_sfr1_n192, oc8051_sfr1_n191, oc8051_sfr1_n190,
         oc8051_sfr1_n189, oc8051_sfr1_n188, oc8051_sfr1_n187,
         oc8051_sfr1_n186, oc8051_sfr1_n185, oc8051_sfr1_n184,
         oc8051_sfr1_n183, oc8051_sfr1_n182, oc8051_sfr1_n181,
         oc8051_sfr1_n180, oc8051_sfr1_n179, oc8051_sfr1_n178,
         oc8051_sfr1_n177, oc8051_sfr1_n176, oc8051_sfr1_n175,
         oc8051_sfr1_n174, oc8051_sfr1_n173, oc8051_sfr1_n172,
         oc8051_sfr1_n171, oc8051_sfr1_n170, oc8051_sfr1_n169,
         oc8051_sfr1_n168, oc8051_sfr1_n167, oc8051_sfr1_n166,
         oc8051_sfr1_n165, oc8051_sfr1_n164, oc8051_sfr1_n163,
         oc8051_sfr1_n162, oc8051_sfr1_n161, oc8051_sfr1_n160,
         oc8051_sfr1_n159, oc8051_sfr1_n158, oc8051_sfr1_n157,
         oc8051_sfr1_n156, oc8051_sfr1_n155, oc8051_sfr1_n154,
         oc8051_sfr1_n153, oc8051_sfr1_n152, oc8051_sfr1_n151,
         oc8051_sfr1_n150, oc8051_sfr1_n149, oc8051_sfr1_n148,
         oc8051_sfr1_n147, oc8051_sfr1_n146, oc8051_sfr1_n145,
         oc8051_sfr1_n144, oc8051_sfr1_n143, oc8051_sfr1_n142,
         oc8051_sfr1_n141, oc8051_sfr1_n140, oc8051_sfr1_n139,
         oc8051_sfr1_n138, oc8051_sfr1_n137, oc8051_sfr1_n136,
         oc8051_sfr1_n135, oc8051_sfr1_n134, oc8051_sfr1_n133,
         oc8051_sfr1_n132, oc8051_sfr1_n131, oc8051_sfr1_n130,
         oc8051_sfr1_n129, oc8051_sfr1_n128, oc8051_sfr1_n127,
         oc8051_sfr1_n126, oc8051_sfr1_n125, oc8051_sfr1_n124,
         oc8051_sfr1_n123, oc8051_sfr1_n122, oc8051_sfr1_n121,
         oc8051_sfr1_n120, oc8051_sfr1_n119, oc8051_sfr1_n118,
         oc8051_sfr1_n117, oc8051_sfr1_n116, oc8051_sfr1_n115,
         oc8051_sfr1_n114, oc8051_sfr1_n113, oc8051_sfr1_n112,
         oc8051_sfr1_n111, oc8051_sfr1_n110, oc8051_sfr1_n109,
         oc8051_sfr1_n108, oc8051_sfr1_n107, oc8051_sfr1_n106,
         oc8051_sfr1_n105, oc8051_sfr1_n104, oc8051_sfr1_n103,
         oc8051_sfr1_n102, oc8051_sfr1_n101, oc8051_sfr1_n100, oc8051_sfr1_n99,
         oc8051_sfr1_n98, oc8051_sfr1_n97, oc8051_sfr1_n96, oc8051_sfr1_n95,
         oc8051_sfr1_n94, oc8051_sfr1_n93, oc8051_sfr1_n92, oc8051_sfr1_n91,
         oc8051_sfr1_n90, oc8051_sfr1_n89, oc8051_sfr1_n88, oc8051_sfr1_n87,
         oc8051_sfr1_n86, oc8051_sfr1_n85, oc8051_sfr1_n84, oc8051_sfr1_n83,
         oc8051_sfr1_n82, oc8051_sfr1_n81, oc8051_sfr1_n80, oc8051_sfr1_n79,
         oc8051_sfr1_n78, oc8051_sfr1_n77, oc8051_sfr1_n76, oc8051_sfr1_n75,
         oc8051_sfr1_n74, oc8051_sfr1_n73, oc8051_sfr1_n72, oc8051_sfr1_n71,
         oc8051_sfr1_n70, oc8051_sfr1_n69, oc8051_sfr1_n68, oc8051_sfr1_n67,
         oc8051_sfr1_n66, oc8051_sfr1_n65, oc8051_sfr1_n64, oc8051_sfr1_n63,
         oc8051_sfr1_n62, oc8051_sfr1_n61, oc8051_sfr1_n60, oc8051_sfr1_n59,
         oc8051_sfr1_n58, oc8051_sfr1_n57, oc8051_sfr1_n56, oc8051_sfr1_n55,
         oc8051_sfr1_n54, oc8051_sfr1_n53, oc8051_sfr1_n52, oc8051_sfr1_n51,
         oc8051_sfr1_n50, oc8051_sfr1_n49, oc8051_sfr1_n48, oc8051_sfr1_n47,
         oc8051_sfr1_n46, oc8051_sfr1_n45, oc8051_sfr1_n44, oc8051_sfr1_n43,
         oc8051_sfr1_n42, oc8051_sfr1_n41, oc8051_sfr1_n40, oc8051_sfr1_n39,
         oc8051_sfr1_n38, oc8051_sfr1_n37, oc8051_sfr1_n36, oc8051_sfr1_n35,
         oc8051_sfr1_n34, oc8051_sfr1_n33, oc8051_sfr1_n32, oc8051_sfr1_n31,
         oc8051_sfr1_n30, oc8051_sfr1_n29, oc8051_sfr1_n28, oc8051_sfr1_n27,
         oc8051_sfr1_n26, oc8051_sfr1_n25, oc8051_sfr1_n24, oc8051_sfr1_n23,
         oc8051_sfr1_n22, oc8051_sfr1_n21, oc8051_sfr1_n20, oc8051_sfr1_n19,
         oc8051_sfr1_n18, oc8051_sfr1_n17, oc8051_sfr1_n16, oc8051_sfr1_n15,
         oc8051_sfr1_n14, oc8051_sfr1_n13, oc8051_sfr1_n12, oc8051_sfr1_n11,
         oc8051_sfr1_n10, oc8051_sfr1_n9, oc8051_sfr1_n8, oc8051_sfr1_n7,
         oc8051_sfr1_n6, oc8051_sfr1_n5, oc8051_sfr1_n4, oc8051_sfr1_n3,
         oc8051_sfr1_n2, oc8051_sfr1_int_src_2_, oc8051_sfr1_n244,
         oc8051_sfr1_n243, oc8051_sfr1_n242, oc8051_sfr1_n241,
         oc8051_sfr1_n240, oc8051_sfr1_n239, oc8051_sfr1_n238,
         oc8051_sfr1_n237, oc8051_sfr1_n1520, oc8051_sfr1_n1510,
         oc8051_sfr1_n1500, oc8051_sfr1_prescaler_0_, oc8051_sfr1_prescaler_1_,
         oc8051_sfr1_prescaler_2_, oc8051_sfr1_prescaler_3_, oc8051_sfr1_n1400,
         oc8051_sfr1_n1380, oc8051_sfr1_n1370, oc8051_sfr1_n1360,
         oc8051_sfr1_n1350, oc8051_sfr1_n1340, oc8051_sfr1_n1330,
         oc8051_sfr1_n1320, oc8051_sfr1_n1310, oc8051_sfr1_n1300,
         oc8051_sfr1_n1290, oc8051_sfr1_n1280, oc8051_sfr1_n1270,
         oc8051_sfr1_n1020, oc8051_sfr1_t2con_0_, oc8051_sfr1_t2con_1_,
         oc8051_sfr1_t2con_2_, oc8051_sfr1_t2con_3_, oc8051_sfr1_t2con_6_,
         oc8051_sfr1_t2con_7_, oc8051_sfr1_ip_0_, oc8051_sfr1_ip_1_,
         oc8051_sfr1_ip_2_, oc8051_sfr1_ip_3_, oc8051_sfr1_ip_4_,
         oc8051_sfr1_ip_5_, oc8051_sfr1_ip_6_, oc8051_sfr1_ip_7_,
         oc8051_sfr1_tcon_0_, oc8051_sfr1_tcon_1_, oc8051_sfr1_tcon_2_,
         oc8051_sfr1_tcon_3_, oc8051_sfr1_tcon_5_, oc8051_sfr1_tcon_7_,
         oc8051_sfr1_ie_0_, oc8051_sfr1_ie_1_, oc8051_sfr1_ie_2_,
         oc8051_sfr1_ie_3_, oc8051_sfr1_ie_4_, oc8051_sfr1_ie_5_,
         oc8051_sfr1_ie_6_, oc8051_sfr1_ie_7_, oc8051_sfr1_tr1,
         oc8051_sfr1_tr0, oc8051_sfr1_tc2_int, oc8051_sfr1_tf0,
         oc8051_sfr1_scon_0_, oc8051_sfr1_scon_1_, oc8051_sfr1_scon_2_,
         oc8051_sfr1_scon_3_, oc8051_sfr1_scon_4_, oc8051_sfr1_scon_5_,
         oc8051_sfr1_scon_6_, oc8051_sfr1_scon_7_, oc8051_sfr1_tclk,
         oc8051_sfr1_rclk, oc8051_sfr1_pres_ow, oc8051_sfr1_tf1,
         oc8051_sfr1_brate2, oc8051_sfr1_uart_int, oc8051_sfr1_p3_data_0_,
         oc8051_sfr1_p3_data_1_, oc8051_sfr1_p3_data_2_,
         oc8051_sfr1_p3_data_3_, oc8051_sfr1_p3_data_4_,
         oc8051_sfr1_p3_data_5_, oc8051_sfr1_p3_data_6_,
         oc8051_sfr1_p3_data_7_, oc8051_sfr1_p2_data_0_,
         oc8051_sfr1_p2_data_1_, oc8051_sfr1_p2_data_2_,
         oc8051_sfr1_p2_data_3_, oc8051_sfr1_p2_data_4_,
         oc8051_sfr1_p2_data_5_, oc8051_sfr1_p2_data_6_,
         oc8051_sfr1_p2_data_7_, oc8051_sfr1_p1_data_0_,
         oc8051_sfr1_p1_data_1_, oc8051_sfr1_p1_data_2_,
         oc8051_sfr1_p1_data_3_, oc8051_sfr1_p1_data_4_,
         oc8051_sfr1_p1_data_5_, oc8051_sfr1_p1_data_6_,
         oc8051_sfr1_p1_data_7_, oc8051_sfr1_p0_data_0_,
         oc8051_sfr1_p0_data_1_, oc8051_sfr1_p0_data_2_,
         oc8051_sfr1_p0_data_3_, oc8051_sfr1_p0_data_4_,
         oc8051_sfr1_p0_data_5_, oc8051_sfr1_p0_data_6_,
         oc8051_sfr1_p0_data_7_, oc8051_sfr1_b_reg_0_, oc8051_sfr1_b_reg_1_,
         oc8051_sfr1_b_reg_2_, oc8051_sfr1_b_reg_3_, oc8051_sfr1_b_reg_4_,
         oc8051_sfr1_b_reg_5_, oc8051_sfr1_b_reg_6_, oc8051_sfr1_b_reg_7_,
         oc8051_sfr1_wr_bit_r, oc8051_sfr1_psw_0_, oc8051_sfr1_psw_1_,
         oc8051_sfr1_psw_2_, oc8051_sfr1_psw_3_, oc8051_sfr1_psw_4_,
         oc8051_sfr1_psw_5_, oc8051_sfr1_oc8051_acc1_n66,
         oc8051_sfr1_oc8051_acc1_n65, oc8051_sfr1_oc8051_acc1_n64,
         oc8051_sfr1_oc8051_acc1_n63, oc8051_sfr1_oc8051_acc1_n62,
         oc8051_sfr1_oc8051_acc1_n61, oc8051_sfr1_oc8051_acc1_n60,
         oc8051_sfr1_oc8051_acc1_n59, oc8051_sfr1_oc8051_acc1_n58,
         oc8051_sfr1_oc8051_acc1_n57, oc8051_sfr1_oc8051_acc1_n56,
         oc8051_sfr1_oc8051_acc1_n55, oc8051_sfr1_oc8051_acc1_n54,
         oc8051_sfr1_oc8051_acc1_n53, oc8051_sfr1_oc8051_acc1_n52,
         oc8051_sfr1_oc8051_acc1_n51, oc8051_sfr1_oc8051_acc1_n50,
         oc8051_sfr1_oc8051_acc1_n49, oc8051_sfr1_oc8051_acc1_n48,
         oc8051_sfr1_oc8051_acc1_n47, oc8051_sfr1_oc8051_acc1_n46,
         oc8051_sfr1_oc8051_acc1_n45, oc8051_sfr1_oc8051_acc1_n44,
         oc8051_sfr1_oc8051_acc1_n43, oc8051_sfr1_oc8051_acc1_n42,
         oc8051_sfr1_oc8051_acc1_n41, oc8051_sfr1_oc8051_acc1_n40,
         oc8051_sfr1_oc8051_acc1_n39, oc8051_sfr1_oc8051_acc1_n38,
         oc8051_sfr1_oc8051_acc1_n37, oc8051_sfr1_oc8051_acc1_n36,
         oc8051_sfr1_oc8051_acc1_n35, oc8051_sfr1_oc8051_acc1_n34,
         oc8051_sfr1_oc8051_acc1_n33, oc8051_sfr1_oc8051_acc1_n32,
         oc8051_sfr1_oc8051_acc1_n31, oc8051_sfr1_oc8051_acc1_n30,
         oc8051_sfr1_oc8051_acc1_n29, oc8051_sfr1_oc8051_acc1_n28,
         oc8051_sfr1_oc8051_acc1_n27, oc8051_sfr1_oc8051_acc1_n26,
         oc8051_sfr1_oc8051_acc1_n25, oc8051_sfr1_oc8051_acc1_n24,
         oc8051_sfr1_oc8051_acc1_n23, oc8051_sfr1_oc8051_acc1_n22,
         oc8051_sfr1_oc8051_acc1_n21, oc8051_sfr1_oc8051_acc1_n20,
         oc8051_sfr1_oc8051_acc1_n19, oc8051_sfr1_oc8051_acc1_n18,
         oc8051_sfr1_oc8051_acc1_n17, oc8051_sfr1_oc8051_acc1_n16,
         oc8051_sfr1_oc8051_acc1_n15, oc8051_sfr1_oc8051_acc1_n14,
         oc8051_sfr1_oc8051_acc1_n13, oc8051_sfr1_oc8051_acc1_n12,
         oc8051_sfr1_oc8051_acc1_n11, oc8051_sfr1_oc8051_acc1_n10,
         oc8051_sfr1_oc8051_acc1_n9, oc8051_sfr1_oc8051_acc1_n8,
         oc8051_sfr1_oc8051_acc1_n7, oc8051_sfr1_oc8051_acc1_n6,
         oc8051_sfr1_oc8051_acc1_n5, oc8051_sfr1_oc8051_acc1_n4,
         oc8051_sfr1_oc8051_acc1_n3, oc8051_sfr1_oc8051_acc1_n2,
         oc8051_sfr1_oc8051_acc1_n1, oc8051_sfr1_oc8051_acc1_acc_0_,
         oc8051_sfr1_oc8051_acc1_acc_1_, oc8051_sfr1_oc8051_acc1_acc_2_,
         oc8051_sfr1_oc8051_acc1_acc_3_, oc8051_sfr1_oc8051_acc1_acc_4_,
         oc8051_sfr1_oc8051_acc1_acc_5_, oc8051_sfr1_oc8051_acc1_acc_6_,
         oc8051_sfr1_oc8051_acc1_acc_7_, oc8051_sfr1_oc8051_b_register_n28,
         oc8051_sfr1_oc8051_b_register_n27, oc8051_sfr1_oc8051_b_register_n26,
         oc8051_sfr1_oc8051_b_register_n25, oc8051_sfr1_oc8051_b_register_n24,
         oc8051_sfr1_oc8051_b_register_n23, oc8051_sfr1_oc8051_b_register_n22,
         oc8051_sfr1_oc8051_b_register_n21, oc8051_sfr1_oc8051_b_register_n20,
         oc8051_sfr1_oc8051_b_register_n19, oc8051_sfr1_oc8051_b_register_n18,
         oc8051_sfr1_oc8051_b_register_n17, oc8051_sfr1_oc8051_b_register_n16,
         oc8051_sfr1_oc8051_b_register_n15, oc8051_sfr1_oc8051_b_register_n14,
         oc8051_sfr1_oc8051_b_register_n13, oc8051_sfr1_oc8051_b_register_n12,
         oc8051_sfr1_oc8051_b_register_n11, oc8051_sfr1_oc8051_b_register_n10,
         oc8051_sfr1_oc8051_b_register_n9, oc8051_sfr1_oc8051_b_register_n8,
         oc8051_sfr1_oc8051_b_register_n7, oc8051_sfr1_oc8051_b_register_n6,
         oc8051_sfr1_oc8051_b_register_n5, oc8051_sfr1_oc8051_b_register_n4,
         oc8051_sfr1_oc8051_b_register_n3, oc8051_sfr1_oc8051_b_register_n2,
         oc8051_sfr1_oc8051_b_register_n1, oc8051_sfr1_oc8051_b_register_n39,
         oc8051_sfr1_oc8051_b_register_n38, oc8051_sfr1_oc8051_b_register_n37,
         oc8051_sfr1_oc8051_b_register_n36, oc8051_sfr1_oc8051_b_register_n35,
         oc8051_sfr1_oc8051_b_register_n34, oc8051_sfr1_oc8051_b_register_n33,
         oc8051_sfr1_oc8051_b_register_n32, oc8051_sfr1_oc8051_sp1_n5,
         oc8051_sfr1_oc8051_sp1_n4, oc8051_sfr1_oc8051_sp1_n3,
         oc8051_sfr1_oc8051_sp1_n2, oc8051_sfr1_oc8051_sp1_n1,
         oc8051_sfr1_oc8051_sp1_r313_carry_7_,
         oc8051_sfr1_oc8051_sp1_r313_carry_6_,
         oc8051_sfr1_oc8051_sp1_r313_carry_5_,
         oc8051_sfr1_oc8051_sp1_r313_carry_4_,
         oc8051_sfr1_oc8051_sp1_r313_carry_3_,
         oc8051_sfr1_oc8051_sp1_r313_carry_2_,
         oc8051_sfr1_oc8051_sp1_r313_carry_1_,
         oc8051_sfr1_oc8051_sp1_r313_b_as_0_, oc8051_sfr1_oc8051_sp1_n22,
         oc8051_sfr1_oc8051_sp1_u3_u2_z_0, oc8051_sfr1_oc8051_sp1_pop,
         oc8051_sfr1_oc8051_sp1_n31, oc8051_sfr1_oc8051_sp1_n30,
         oc8051_sfr1_oc8051_sp1_n29, oc8051_sfr1_oc8051_sp1_n28,
         oc8051_sfr1_oc8051_sp1_n27, oc8051_sfr1_oc8051_sp1_n26,
         oc8051_sfr1_oc8051_sp1_n25, oc8051_sfr1_oc8051_sp1_n24,
         oc8051_sfr1_oc8051_sp1_n20, oc8051_sfr1_oc8051_sp1_n19,
         oc8051_sfr1_oc8051_sp1_n18, oc8051_sfr1_oc8051_sp1_n17,
         oc8051_sfr1_oc8051_sp1_n16, oc8051_sfr1_oc8051_sp1_n15,
         oc8051_sfr1_oc8051_sp1_n14, oc8051_sfr1_oc8051_sp1_n13,
         oc8051_sfr1_oc8051_sp1_sp_0_, oc8051_sfr1_oc8051_sp1_sp_1_,
         oc8051_sfr1_oc8051_sp1_sp_2_, oc8051_sfr1_oc8051_sp1_sp_3_,
         oc8051_sfr1_oc8051_sp1_sp_4_, oc8051_sfr1_oc8051_sp1_sp_5_,
         oc8051_sfr1_oc8051_sp1_sp_6_, oc8051_sfr1_oc8051_sp1_sp_7_,
         oc8051_sfr1_oc8051_dptr1_n15, oc8051_sfr1_oc8051_dptr1_n14,
         oc8051_sfr1_oc8051_dptr1_n13, oc8051_sfr1_oc8051_dptr1_n12,
         oc8051_sfr1_oc8051_dptr1_n11, oc8051_sfr1_oc8051_dptr1_n10,
         oc8051_sfr1_oc8051_dptr1_n9, oc8051_sfr1_oc8051_dptr1_n8,
         oc8051_sfr1_oc8051_dptr1_n7, oc8051_sfr1_oc8051_dptr1_n6,
         oc8051_sfr1_oc8051_dptr1_n5, oc8051_sfr1_oc8051_dptr1_n4,
         oc8051_sfr1_oc8051_dptr1_n3, oc8051_sfr1_oc8051_dptr1_n2,
         oc8051_sfr1_oc8051_dptr1_n1, oc8051_sfr1_oc8051_dptr1_n33,
         oc8051_sfr1_oc8051_dptr1_n32, oc8051_sfr1_oc8051_dptr1_n31,
         oc8051_sfr1_oc8051_dptr1_n30, oc8051_sfr1_oc8051_dptr1_n29,
         oc8051_sfr1_oc8051_dptr1_n28, oc8051_sfr1_oc8051_dptr1_n27,
         oc8051_sfr1_oc8051_dptr1_n26, oc8051_sfr1_oc8051_dptr1_n25,
         oc8051_sfr1_oc8051_dptr1_n24, oc8051_sfr1_oc8051_dptr1_n23,
         oc8051_sfr1_oc8051_dptr1_n22, oc8051_sfr1_oc8051_dptr1_n21,
         oc8051_sfr1_oc8051_dptr1_n20, oc8051_sfr1_oc8051_dptr1_n19,
         oc8051_sfr1_oc8051_dptr1_n18, oc8051_sfr1_oc8051_psw1_n40,
         oc8051_sfr1_oc8051_psw1_n39, oc8051_sfr1_oc8051_psw1_n38,
         oc8051_sfr1_oc8051_psw1_n37, oc8051_sfr1_oc8051_psw1_n36,
         oc8051_sfr1_oc8051_psw1_n35, oc8051_sfr1_oc8051_psw1_n34,
         oc8051_sfr1_oc8051_psw1_n33, oc8051_sfr1_oc8051_psw1_n32,
         oc8051_sfr1_oc8051_psw1_n31, oc8051_sfr1_oc8051_psw1_n30,
         oc8051_sfr1_oc8051_psw1_n29, oc8051_sfr1_oc8051_psw1_n28,
         oc8051_sfr1_oc8051_psw1_n27, oc8051_sfr1_oc8051_psw1_n26,
         oc8051_sfr1_oc8051_psw1_n25, oc8051_sfr1_oc8051_psw1_n24,
         oc8051_sfr1_oc8051_psw1_n23, oc8051_sfr1_oc8051_psw1_n22,
         oc8051_sfr1_oc8051_psw1_n21, oc8051_sfr1_oc8051_psw1_n20,
         oc8051_sfr1_oc8051_psw1_n19, oc8051_sfr1_oc8051_psw1_n18,
         oc8051_sfr1_oc8051_psw1_n17, oc8051_sfr1_oc8051_psw1_n16,
         oc8051_sfr1_oc8051_psw1_n15, oc8051_sfr1_oc8051_psw1_n14,
         oc8051_sfr1_oc8051_psw1_n13, oc8051_sfr1_oc8051_psw1_n12,
         oc8051_sfr1_oc8051_psw1_n11, oc8051_sfr1_oc8051_psw1_n10,
         oc8051_sfr1_oc8051_psw1_n9, oc8051_sfr1_oc8051_psw1_n8,
         oc8051_sfr1_oc8051_psw1_n7, oc8051_sfr1_oc8051_psw1_n6,
         oc8051_sfr1_oc8051_psw1_n5, oc8051_sfr1_oc8051_psw1_n4,
         oc8051_sfr1_oc8051_psw1_n3, oc8051_sfr1_oc8051_psw1_n2,
         oc8051_sfr1_oc8051_psw1_n49, oc8051_sfr1_oc8051_psw1_n48,
         oc8051_sfr1_oc8051_psw1_n47, oc8051_sfr1_oc8051_psw1_n46,
         oc8051_sfr1_oc8051_psw1_n45, oc8051_sfr1_oc8051_psw1_n44,
         oc8051_sfr1_oc8051_psw1_n43, oc8051_sfr1_oc8051_psw1_n1,
         oc8051_sfr1_oc8051_ports1_n106, oc8051_sfr1_oc8051_ports1_n105,
         oc8051_sfr1_oc8051_ports1_n104, oc8051_sfr1_oc8051_ports1_n103,
         oc8051_sfr1_oc8051_ports1_n102, oc8051_sfr1_oc8051_ports1_n101,
         oc8051_sfr1_oc8051_ports1_n100, oc8051_sfr1_oc8051_ports1_n99,
         oc8051_sfr1_oc8051_ports1_n98, oc8051_sfr1_oc8051_ports1_n97,
         oc8051_sfr1_oc8051_ports1_n96, oc8051_sfr1_oc8051_ports1_n95,
         oc8051_sfr1_oc8051_ports1_n94, oc8051_sfr1_oc8051_ports1_n93,
         oc8051_sfr1_oc8051_ports1_n92, oc8051_sfr1_oc8051_ports1_n91,
         oc8051_sfr1_oc8051_ports1_n90, oc8051_sfr1_oc8051_ports1_n89,
         oc8051_sfr1_oc8051_ports1_n88, oc8051_sfr1_oc8051_ports1_n87,
         oc8051_sfr1_oc8051_ports1_n86, oc8051_sfr1_oc8051_ports1_n85,
         oc8051_sfr1_oc8051_ports1_n84, oc8051_sfr1_oc8051_ports1_n83,
         oc8051_sfr1_oc8051_ports1_n82, oc8051_sfr1_oc8051_ports1_n81,
         oc8051_sfr1_oc8051_ports1_n80, oc8051_sfr1_oc8051_ports1_n79,
         oc8051_sfr1_oc8051_ports1_n78, oc8051_sfr1_oc8051_ports1_n77,
         oc8051_sfr1_oc8051_ports1_n76, oc8051_sfr1_oc8051_ports1_n75,
         oc8051_sfr1_oc8051_ports1_n74, oc8051_sfr1_oc8051_ports1_n73,
         oc8051_sfr1_oc8051_ports1_n72, oc8051_sfr1_oc8051_ports1_n71,
         oc8051_sfr1_oc8051_ports1_n70, oc8051_sfr1_oc8051_ports1_n69,
         oc8051_sfr1_oc8051_ports1_n68, oc8051_sfr1_oc8051_ports1_n67,
         oc8051_sfr1_oc8051_ports1_n66, oc8051_sfr1_oc8051_ports1_n65,
         oc8051_sfr1_oc8051_ports1_n64, oc8051_sfr1_oc8051_ports1_n63,
         oc8051_sfr1_oc8051_ports1_n62, oc8051_sfr1_oc8051_ports1_n61,
         oc8051_sfr1_oc8051_ports1_n60, oc8051_sfr1_oc8051_ports1_n59,
         oc8051_sfr1_oc8051_ports1_n58, oc8051_sfr1_oc8051_ports1_n57,
         oc8051_sfr1_oc8051_ports1_n56, oc8051_sfr1_oc8051_ports1_n55,
         oc8051_sfr1_oc8051_ports1_n54, oc8051_sfr1_oc8051_ports1_n53,
         oc8051_sfr1_oc8051_ports1_n52, oc8051_sfr1_oc8051_ports1_n51,
         oc8051_sfr1_oc8051_ports1_n50, oc8051_sfr1_oc8051_ports1_n49,
         oc8051_sfr1_oc8051_ports1_n48, oc8051_sfr1_oc8051_ports1_n47,
         oc8051_sfr1_oc8051_ports1_n46, oc8051_sfr1_oc8051_ports1_n45,
         oc8051_sfr1_oc8051_ports1_n44, oc8051_sfr1_oc8051_ports1_n43,
         oc8051_sfr1_oc8051_ports1_n42, oc8051_sfr1_oc8051_ports1_n41,
         oc8051_sfr1_oc8051_ports1_n40, oc8051_sfr1_oc8051_ports1_n39,
         oc8051_sfr1_oc8051_ports1_n38, oc8051_sfr1_oc8051_ports1_n37,
         oc8051_sfr1_oc8051_ports1_n36, oc8051_sfr1_oc8051_ports1_n35,
         oc8051_sfr1_oc8051_ports1_n34, oc8051_sfr1_oc8051_ports1_n33,
         oc8051_sfr1_oc8051_ports1_n32, oc8051_sfr1_oc8051_ports1_n31,
         oc8051_sfr1_oc8051_ports1_n30, oc8051_sfr1_oc8051_ports1_n29,
         oc8051_sfr1_oc8051_ports1_n28, oc8051_sfr1_oc8051_ports1_n27,
         oc8051_sfr1_oc8051_ports1_n26, oc8051_sfr1_oc8051_ports1_n25,
         oc8051_sfr1_oc8051_ports1_n24, oc8051_sfr1_oc8051_ports1_n23,
         oc8051_sfr1_oc8051_ports1_n22, oc8051_sfr1_oc8051_ports1_n21,
         oc8051_sfr1_oc8051_ports1_n20, oc8051_sfr1_oc8051_ports1_n19,
         oc8051_sfr1_oc8051_ports1_n18, oc8051_sfr1_oc8051_ports1_n17,
         oc8051_sfr1_oc8051_ports1_n16, oc8051_sfr1_oc8051_ports1_n15,
         oc8051_sfr1_oc8051_ports1_n14, oc8051_sfr1_oc8051_ports1_n13,
         oc8051_sfr1_oc8051_ports1_n12, oc8051_sfr1_oc8051_ports1_n11,
         oc8051_sfr1_oc8051_ports1_n10, oc8051_sfr1_oc8051_ports1_n9,
         oc8051_sfr1_oc8051_ports1_n8, oc8051_sfr1_oc8051_ports1_n7,
         oc8051_sfr1_oc8051_ports1_n6, oc8051_sfr1_oc8051_ports1_n5,
         oc8051_sfr1_oc8051_ports1_n4, oc8051_sfr1_oc8051_ports1_n3,
         oc8051_sfr1_oc8051_ports1_n2, oc8051_sfr1_oc8051_ports1_n1,
         oc8051_sfr1_oc8051_ports1_n163, oc8051_sfr1_oc8051_ports1_n162,
         oc8051_sfr1_oc8051_ports1_n161, oc8051_sfr1_oc8051_ports1_n160,
         oc8051_sfr1_oc8051_ports1_n159, oc8051_sfr1_oc8051_ports1_n158,
         oc8051_sfr1_oc8051_ports1_n157, oc8051_sfr1_oc8051_ports1_n156,
         oc8051_sfr1_oc8051_ports1_n155, oc8051_sfr1_oc8051_ports1_n154,
         oc8051_sfr1_oc8051_ports1_n153, oc8051_sfr1_oc8051_ports1_n152,
         oc8051_sfr1_oc8051_ports1_n151, oc8051_sfr1_oc8051_ports1_n150,
         oc8051_sfr1_oc8051_ports1_n149, oc8051_sfr1_oc8051_ports1_n148,
         oc8051_sfr1_oc8051_ports1_n147, oc8051_sfr1_oc8051_ports1_n146,
         oc8051_sfr1_oc8051_ports1_n145, oc8051_sfr1_oc8051_ports1_n144,
         oc8051_sfr1_oc8051_ports1_n143, oc8051_sfr1_oc8051_ports1_n142,
         oc8051_sfr1_oc8051_ports1_n141, oc8051_sfr1_oc8051_ports1_n140,
         oc8051_sfr1_oc8051_ports1_n139, oc8051_sfr1_oc8051_ports1_n138,
         oc8051_sfr1_oc8051_ports1_n137, oc8051_sfr1_oc8051_ports1_n136,
         oc8051_sfr1_oc8051_ports1_n135, oc8051_sfr1_oc8051_ports1_n134,
         oc8051_sfr1_oc8051_ports1_n133, oc8051_sfr1_oc8051_ports1_n132,
         oc8051_sfr1_oc8051_uatr1_n168, oc8051_sfr1_oc8051_uatr1_n166,
         oc8051_sfr1_oc8051_uatr1_n165, oc8051_sfr1_oc8051_uatr1_n164,
         oc8051_sfr1_oc8051_uatr1_n163, oc8051_sfr1_oc8051_uatr1_n162,
         oc8051_sfr1_oc8051_uatr1_n161, oc8051_sfr1_oc8051_uatr1_n160,
         oc8051_sfr1_oc8051_uatr1_n159, oc8051_sfr1_oc8051_uatr1_n158,
         oc8051_sfr1_oc8051_uatr1_n157, oc8051_sfr1_oc8051_uatr1_n156,
         oc8051_sfr1_oc8051_uatr1_n155, oc8051_sfr1_oc8051_uatr1_n154,
         oc8051_sfr1_oc8051_uatr1_n153, oc8051_sfr1_oc8051_uatr1_n152,
         oc8051_sfr1_oc8051_uatr1_n151, oc8051_sfr1_oc8051_uatr1_n150,
         oc8051_sfr1_oc8051_uatr1_n149, oc8051_sfr1_oc8051_uatr1_n148,
         oc8051_sfr1_oc8051_uatr1_n147, oc8051_sfr1_oc8051_uatr1_n146,
         oc8051_sfr1_oc8051_uatr1_n145, oc8051_sfr1_oc8051_uatr1_n144,
         oc8051_sfr1_oc8051_uatr1_n143, oc8051_sfr1_oc8051_uatr1_n142,
         oc8051_sfr1_oc8051_uatr1_n141, oc8051_sfr1_oc8051_uatr1_n140,
         oc8051_sfr1_oc8051_uatr1_n139, oc8051_sfr1_oc8051_uatr1_n138,
         oc8051_sfr1_oc8051_uatr1_n137, oc8051_sfr1_oc8051_uatr1_n136,
         oc8051_sfr1_oc8051_uatr1_n135, oc8051_sfr1_oc8051_uatr1_n134,
         oc8051_sfr1_oc8051_uatr1_n133, oc8051_sfr1_oc8051_uatr1_n132,
         oc8051_sfr1_oc8051_uatr1_n131, oc8051_sfr1_oc8051_uatr1_n130,
         oc8051_sfr1_oc8051_uatr1_n129, oc8051_sfr1_oc8051_uatr1_n128,
         oc8051_sfr1_oc8051_uatr1_n127, oc8051_sfr1_oc8051_uatr1_n126,
         oc8051_sfr1_oc8051_uatr1_n125, oc8051_sfr1_oc8051_uatr1_n124,
         oc8051_sfr1_oc8051_uatr1_n123, oc8051_sfr1_oc8051_uatr1_n122,
         oc8051_sfr1_oc8051_uatr1_n121, oc8051_sfr1_oc8051_uatr1_n120,
         oc8051_sfr1_oc8051_uatr1_n119, oc8051_sfr1_oc8051_uatr1_n118,
         oc8051_sfr1_oc8051_uatr1_n117, oc8051_sfr1_oc8051_uatr1_n116,
         oc8051_sfr1_oc8051_uatr1_n115, oc8051_sfr1_oc8051_uatr1_n114,
         oc8051_sfr1_oc8051_uatr1_n113, oc8051_sfr1_oc8051_uatr1_n112,
         oc8051_sfr1_oc8051_uatr1_n111, oc8051_sfr1_oc8051_uatr1_n110,
         oc8051_sfr1_oc8051_uatr1_n109, oc8051_sfr1_oc8051_uatr1_n108,
         oc8051_sfr1_oc8051_uatr1_n107, oc8051_sfr1_oc8051_uatr1_n106,
         oc8051_sfr1_oc8051_uatr1_n105, oc8051_sfr1_oc8051_uatr1_n104,
         oc8051_sfr1_oc8051_uatr1_n103, oc8051_sfr1_oc8051_uatr1_n102,
         oc8051_sfr1_oc8051_uatr1_n101, oc8051_sfr1_oc8051_uatr1_n100,
         oc8051_sfr1_oc8051_uatr1_n99, oc8051_sfr1_oc8051_uatr1_n98,
         oc8051_sfr1_oc8051_uatr1_n97, oc8051_sfr1_oc8051_uatr1_n96,
         oc8051_sfr1_oc8051_uatr1_n95, oc8051_sfr1_oc8051_uatr1_n94,
         oc8051_sfr1_oc8051_uatr1_n93, oc8051_sfr1_oc8051_uatr1_n92,
         oc8051_sfr1_oc8051_uatr1_n91, oc8051_sfr1_oc8051_uatr1_n90,
         oc8051_sfr1_oc8051_uatr1_n89, oc8051_sfr1_oc8051_uatr1_n88,
         oc8051_sfr1_oc8051_uatr1_n87, oc8051_sfr1_oc8051_uatr1_n86,
         oc8051_sfr1_oc8051_uatr1_n85, oc8051_sfr1_oc8051_uatr1_n84,
         oc8051_sfr1_oc8051_uatr1_n83, oc8051_sfr1_oc8051_uatr1_n82,
         oc8051_sfr1_oc8051_uatr1_n81, oc8051_sfr1_oc8051_uatr1_n80,
         oc8051_sfr1_oc8051_uatr1_n79, oc8051_sfr1_oc8051_uatr1_n78,
         oc8051_sfr1_oc8051_uatr1_n77, oc8051_sfr1_oc8051_uatr1_n76,
         oc8051_sfr1_oc8051_uatr1_n75, oc8051_sfr1_oc8051_uatr1_n74,
         oc8051_sfr1_oc8051_uatr1_n73, oc8051_sfr1_oc8051_uatr1_n72,
         oc8051_sfr1_oc8051_uatr1_n71, oc8051_sfr1_oc8051_uatr1_n70,
         oc8051_sfr1_oc8051_uatr1_n69, oc8051_sfr1_oc8051_uatr1_n68,
         oc8051_sfr1_oc8051_uatr1_n67, oc8051_sfr1_oc8051_uatr1_n66,
         oc8051_sfr1_oc8051_uatr1_n65, oc8051_sfr1_oc8051_uatr1_n64,
         oc8051_sfr1_oc8051_uatr1_n63, oc8051_sfr1_oc8051_uatr1_n62,
         oc8051_sfr1_oc8051_uatr1_n61, oc8051_sfr1_oc8051_uatr1_n60,
         oc8051_sfr1_oc8051_uatr1_n59, oc8051_sfr1_oc8051_uatr1_n58,
         oc8051_sfr1_oc8051_uatr1_n57, oc8051_sfr1_oc8051_uatr1_n56,
         oc8051_sfr1_oc8051_uatr1_n55, oc8051_sfr1_oc8051_uatr1_n54,
         oc8051_sfr1_oc8051_uatr1_n53, oc8051_sfr1_oc8051_uatr1_n52,
         oc8051_sfr1_oc8051_uatr1_n51, oc8051_sfr1_oc8051_uatr1_n50,
         oc8051_sfr1_oc8051_uatr1_n49, oc8051_sfr1_oc8051_uatr1_n48,
         oc8051_sfr1_oc8051_uatr1_n47, oc8051_sfr1_oc8051_uatr1_n46,
         oc8051_sfr1_oc8051_uatr1_n45, oc8051_sfr1_oc8051_uatr1_n44,
         oc8051_sfr1_oc8051_uatr1_n43, oc8051_sfr1_oc8051_uatr1_n42,
         oc8051_sfr1_oc8051_uatr1_n41, oc8051_sfr1_oc8051_uatr1_n40,
         oc8051_sfr1_oc8051_uatr1_n39, oc8051_sfr1_oc8051_uatr1_n38,
         oc8051_sfr1_oc8051_uatr1_n37, oc8051_sfr1_oc8051_uatr1_n36,
         oc8051_sfr1_oc8051_uatr1_n35, oc8051_sfr1_oc8051_uatr1_n34,
         oc8051_sfr1_oc8051_uatr1_n33, oc8051_sfr1_oc8051_uatr1_n32,
         oc8051_sfr1_oc8051_uatr1_n31, oc8051_sfr1_oc8051_uatr1_n30,
         oc8051_sfr1_oc8051_uatr1_n29, oc8051_sfr1_oc8051_uatr1_n28,
         oc8051_sfr1_oc8051_uatr1_n27, oc8051_sfr1_oc8051_uatr1_n26,
         oc8051_sfr1_oc8051_uatr1_n25, oc8051_sfr1_oc8051_uatr1_n24,
         oc8051_sfr1_oc8051_uatr1_n23, oc8051_sfr1_oc8051_uatr1_n22,
         oc8051_sfr1_oc8051_uatr1_n21, oc8051_sfr1_oc8051_uatr1_n20,
         oc8051_sfr1_oc8051_uatr1_n19, oc8051_sfr1_oc8051_uatr1_n18,
         oc8051_sfr1_oc8051_uatr1_n17, oc8051_sfr1_oc8051_uatr1_n16,
         oc8051_sfr1_oc8051_uatr1_n15, oc8051_sfr1_oc8051_uatr1_n14,
         oc8051_sfr1_oc8051_uatr1_n13, oc8051_sfr1_oc8051_uatr1_n12,
         oc8051_sfr1_oc8051_uatr1_n11, oc8051_sfr1_oc8051_uatr1_n10,
         oc8051_sfr1_oc8051_uatr1_n9, oc8051_sfr1_oc8051_uatr1_n8,
         oc8051_sfr1_oc8051_uatr1_n7, oc8051_sfr1_oc8051_uatr1_n6,
         oc8051_sfr1_oc8051_uatr1_n5, oc8051_sfr1_oc8051_uatr1_n4,
         oc8051_sfr1_oc8051_uatr1_n3, oc8051_sfr1_oc8051_uatr1_n2,
         oc8051_sfr1_oc8051_uatr1_n1, oc8051_sfr1_oc8051_uatr1_n254,
         oc8051_sfr1_oc8051_uatr1_n253, oc8051_sfr1_oc8051_uatr1_n252,
         oc8051_sfr1_oc8051_uatr1_n251, oc8051_sfr1_oc8051_uatr1_n250,
         oc8051_sfr1_oc8051_uatr1_n249, oc8051_sfr1_oc8051_uatr1_n248,
         oc8051_sfr1_oc8051_uatr1_n247, oc8051_sfr1_oc8051_uatr1_n246,
         oc8051_sfr1_oc8051_uatr1_n245, oc8051_sfr1_oc8051_uatr1_n244,
         oc8051_sfr1_oc8051_uatr1_n243, oc8051_sfr1_oc8051_uatr1_n242,
         oc8051_sfr1_oc8051_uatr1_n241, oc8051_sfr1_oc8051_uatr1_n240,
         oc8051_sfr1_oc8051_uatr1_n239, oc8051_sfr1_oc8051_uatr1_n238,
         oc8051_sfr1_oc8051_uatr1_n237, oc8051_sfr1_oc8051_uatr1_n236,
         oc8051_sfr1_oc8051_uatr1_n235, oc8051_sfr1_oc8051_uatr1_n234,
         oc8051_sfr1_oc8051_uatr1_n233, oc8051_sfr1_oc8051_uatr1_n232,
         oc8051_sfr1_oc8051_uatr1_n231, oc8051_sfr1_oc8051_uatr1_n230,
         oc8051_sfr1_oc8051_uatr1_n229, oc8051_sfr1_oc8051_uatr1_n228,
         oc8051_sfr1_oc8051_uatr1_n227, oc8051_sfr1_oc8051_uatr1_n226,
         oc8051_sfr1_oc8051_uatr1_n225, oc8051_sfr1_oc8051_uatr1_n224,
         oc8051_sfr1_oc8051_uatr1_n223, oc8051_sfr1_oc8051_uatr1_n222,
         oc8051_sfr1_oc8051_uatr1_n221, oc8051_sfr1_oc8051_uatr1_n220,
         oc8051_sfr1_oc8051_uatr1_n219, oc8051_sfr1_oc8051_uatr1_n218,
         oc8051_sfr1_oc8051_uatr1_n217, oc8051_sfr1_oc8051_uatr1_n216,
         oc8051_sfr1_oc8051_uatr1_n215, oc8051_sfr1_oc8051_uatr1_n214,
         oc8051_sfr1_oc8051_uatr1_n213, oc8051_sfr1_oc8051_uatr1_n212,
         oc8051_sfr1_oc8051_uatr1_n211, oc8051_sfr1_oc8051_uatr1_n210,
         oc8051_sfr1_oc8051_uatr1_n209, oc8051_sfr1_oc8051_uatr1_n208,
         oc8051_sfr1_oc8051_uatr1_n207, oc8051_sfr1_oc8051_uatr1_n206,
         oc8051_sfr1_oc8051_uatr1_n205, oc8051_sfr1_oc8051_uatr1_n204,
         oc8051_sfr1_oc8051_uatr1_n203, oc8051_sfr1_oc8051_uatr1_n202,
         oc8051_sfr1_oc8051_uatr1_n201, oc8051_sfr1_oc8051_uatr1_n200,
         oc8051_sfr1_oc8051_uatr1_n199, oc8051_sfr1_oc8051_uatr1_n198,
         oc8051_sfr1_oc8051_uatr1_n197, oc8051_sfr1_oc8051_uatr1_n196,
         oc8051_sfr1_oc8051_uatr1_n195, oc8051_sfr1_oc8051_uatr1_n194,
         oc8051_sfr1_oc8051_uatr1_n193, oc8051_sfr1_oc8051_uatr1_n192,
         oc8051_sfr1_oc8051_uatr1_n191, oc8051_sfr1_oc8051_uatr1_n190,
         oc8051_sfr1_oc8051_uatr1_n188, oc8051_sfr1_oc8051_uatr1_n187,
         oc8051_sfr1_oc8051_uatr1_n186, oc8051_sfr1_oc8051_uatr1_n185,
         oc8051_sfr1_oc8051_uatr1_n184, oc8051_sfr1_oc8051_uatr1_n183,
         oc8051_sfr1_oc8051_uatr1_n182, oc8051_sfr1_oc8051_uatr1_n181,
         oc8051_sfr1_oc8051_uatr1_n180, oc8051_sfr1_oc8051_uatr1_n269,
         oc8051_sfr1_oc8051_uatr1_smod_clk_re, oc8051_sfr1_oc8051_uatr1_rxd_r,
         oc8051_sfr1_oc8051_uatr1_shift_re, oc8051_sfr1_oc8051_uatr1_rx_sam_0_,
         oc8051_sfr1_oc8051_uatr1_rx_sam_1_,
         oc8051_sfr1_oc8051_uatr1_re_count_0_,
         oc8051_sfr1_oc8051_uatr1_re_count_1_,
         oc8051_sfr1_oc8051_uatr1_re_count_2_,
         oc8051_sfr1_oc8051_uatr1_re_count_3_,
         oc8051_sfr1_oc8051_uatr1_receive, oc8051_sfr1_oc8051_uatr1_n174,
         oc8051_sfr1_oc8051_uatr1_smod_clk_tr,
         oc8051_sfr1_oc8051_uatr1_shift_tr,
         oc8051_sfr1_oc8051_uatr1_tr_count_0_,
         oc8051_sfr1_oc8051_uatr1_tr_count_1_,
         oc8051_sfr1_oc8051_uatr1_tr_count_2_, oc8051_sfr1_oc8051_uatr1_trans,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_6_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_7_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_,
         oc8051_sfr1_oc8051_uatr1_rx_done,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_,
         oc8051_sfr1_oc8051_int1_n204, oc8051_sfr1_oc8051_int1_n203,
         oc8051_sfr1_oc8051_int1_n202, oc8051_sfr1_oc8051_int1_n201,
         oc8051_sfr1_oc8051_int1_n200, oc8051_sfr1_oc8051_int1_n199,
         oc8051_sfr1_oc8051_int1_n198, oc8051_sfr1_oc8051_int1_n197,
         oc8051_sfr1_oc8051_int1_n196, oc8051_sfr1_oc8051_int1_n195,
         oc8051_sfr1_oc8051_int1_n194, oc8051_sfr1_oc8051_int1_n193,
         oc8051_sfr1_oc8051_int1_n192, oc8051_sfr1_oc8051_int1_n191,
         oc8051_sfr1_oc8051_int1_n190, oc8051_sfr1_oc8051_int1_n189,
         oc8051_sfr1_oc8051_int1_n188, oc8051_sfr1_oc8051_int1_n187,
         oc8051_sfr1_oc8051_int1_n186, oc8051_sfr1_oc8051_int1_n185,
         oc8051_sfr1_oc8051_int1_n184, oc8051_sfr1_oc8051_int1_n183,
         oc8051_sfr1_oc8051_int1_n182, oc8051_sfr1_oc8051_int1_n181,
         oc8051_sfr1_oc8051_int1_n180, oc8051_sfr1_oc8051_int1_n179,
         oc8051_sfr1_oc8051_int1_n178, oc8051_sfr1_oc8051_int1_n177,
         oc8051_sfr1_oc8051_int1_n176, oc8051_sfr1_oc8051_int1_n175,
         oc8051_sfr1_oc8051_int1_n174, oc8051_sfr1_oc8051_int1_n173,
         oc8051_sfr1_oc8051_int1_n172, oc8051_sfr1_oc8051_int1_n171,
         oc8051_sfr1_oc8051_int1_n170, oc8051_sfr1_oc8051_int1_n169,
         oc8051_sfr1_oc8051_int1_n168, oc8051_sfr1_oc8051_int1_n167,
         oc8051_sfr1_oc8051_int1_n166, oc8051_sfr1_oc8051_int1_n165,
         oc8051_sfr1_oc8051_int1_n164, oc8051_sfr1_oc8051_int1_n163,
         oc8051_sfr1_oc8051_int1_n162, oc8051_sfr1_oc8051_int1_n161,
         oc8051_sfr1_oc8051_int1_n160, oc8051_sfr1_oc8051_int1_n159,
         oc8051_sfr1_oc8051_int1_n158, oc8051_sfr1_oc8051_int1_n157,
         oc8051_sfr1_oc8051_int1_n156, oc8051_sfr1_oc8051_int1_n155,
         oc8051_sfr1_oc8051_int1_n154, oc8051_sfr1_oc8051_int1_n153,
         oc8051_sfr1_oc8051_int1_n152, oc8051_sfr1_oc8051_int1_n151,
         oc8051_sfr1_oc8051_int1_n150, oc8051_sfr1_oc8051_int1_n149,
         oc8051_sfr1_oc8051_int1_n148, oc8051_sfr1_oc8051_int1_n147,
         oc8051_sfr1_oc8051_int1_n146, oc8051_sfr1_oc8051_int1_n145,
         oc8051_sfr1_oc8051_int1_n144, oc8051_sfr1_oc8051_int1_n143,
         oc8051_sfr1_oc8051_int1_n142, oc8051_sfr1_oc8051_int1_n141,
         oc8051_sfr1_oc8051_int1_n140, oc8051_sfr1_oc8051_int1_n139,
         oc8051_sfr1_oc8051_int1_n138, oc8051_sfr1_oc8051_int1_n137,
         oc8051_sfr1_oc8051_int1_n136, oc8051_sfr1_oc8051_int1_n135,
         oc8051_sfr1_oc8051_int1_n134, oc8051_sfr1_oc8051_int1_n133,
         oc8051_sfr1_oc8051_int1_n132, oc8051_sfr1_oc8051_int1_n131,
         oc8051_sfr1_oc8051_int1_n130, oc8051_sfr1_oc8051_int1_n129,
         oc8051_sfr1_oc8051_int1_n128, oc8051_sfr1_oc8051_int1_n127,
         oc8051_sfr1_oc8051_int1_n126, oc8051_sfr1_oc8051_int1_n125,
         oc8051_sfr1_oc8051_int1_n124, oc8051_sfr1_oc8051_int1_n123,
         oc8051_sfr1_oc8051_int1_n122, oc8051_sfr1_oc8051_int1_n121,
         oc8051_sfr1_oc8051_int1_n120, oc8051_sfr1_oc8051_int1_n119,
         oc8051_sfr1_oc8051_int1_n118, oc8051_sfr1_oc8051_int1_n117,
         oc8051_sfr1_oc8051_int1_n116, oc8051_sfr1_oc8051_int1_n115,
         oc8051_sfr1_oc8051_int1_n114, oc8051_sfr1_oc8051_int1_n113,
         oc8051_sfr1_oc8051_int1_n112, oc8051_sfr1_oc8051_int1_n111,
         oc8051_sfr1_oc8051_int1_n110, oc8051_sfr1_oc8051_int1_n109,
         oc8051_sfr1_oc8051_int1_n108, oc8051_sfr1_oc8051_int1_n107,
         oc8051_sfr1_oc8051_int1_n106, oc8051_sfr1_oc8051_int1_n105,
         oc8051_sfr1_oc8051_int1_n104, oc8051_sfr1_oc8051_int1_n103,
         oc8051_sfr1_oc8051_int1_n102, oc8051_sfr1_oc8051_int1_n101,
         oc8051_sfr1_oc8051_int1_n100, oc8051_sfr1_oc8051_int1_n99,
         oc8051_sfr1_oc8051_int1_n98, oc8051_sfr1_oc8051_int1_n97,
         oc8051_sfr1_oc8051_int1_n96, oc8051_sfr1_oc8051_int1_n95,
         oc8051_sfr1_oc8051_int1_n94, oc8051_sfr1_oc8051_int1_n93,
         oc8051_sfr1_oc8051_int1_n92, oc8051_sfr1_oc8051_int1_n91,
         oc8051_sfr1_oc8051_int1_n90, oc8051_sfr1_oc8051_int1_n89,
         oc8051_sfr1_oc8051_int1_n88, oc8051_sfr1_oc8051_int1_n87,
         oc8051_sfr1_oc8051_int1_n86, oc8051_sfr1_oc8051_int1_n85,
         oc8051_sfr1_oc8051_int1_n84, oc8051_sfr1_oc8051_int1_n83,
         oc8051_sfr1_oc8051_int1_n82, oc8051_sfr1_oc8051_int1_n81,
         oc8051_sfr1_oc8051_int1_n80, oc8051_sfr1_oc8051_int1_n79,
         oc8051_sfr1_oc8051_int1_n78, oc8051_sfr1_oc8051_int1_n77,
         oc8051_sfr1_oc8051_int1_n76, oc8051_sfr1_oc8051_int1_n75,
         oc8051_sfr1_oc8051_int1_n74, oc8051_sfr1_oc8051_int1_n73,
         oc8051_sfr1_oc8051_int1_n72, oc8051_sfr1_oc8051_int1_n71,
         oc8051_sfr1_oc8051_int1_n70, oc8051_sfr1_oc8051_int1_n69,
         oc8051_sfr1_oc8051_int1_n68, oc8051_sfr1_oc8051_int1_n67,
         oc8051_sfr1_oc8051_int1_n66, oc8051_sfr1_oc8051_int1_n65,
         oc8051_sfr1_oc8051_int1_n64, oc8051_sfr1_oc8051_int1_n63,
         oc8051_sfr1_oc8051_int1_n62, oc8051_sfr1_oc8051_int1_n61,
         oc8051_sfr1_oc8051_int1_n60, oc8051_sfr1_oc8051_int1_n59,
         oc8051_sfr1_oc8051_int1_n58, oc8051_sfr1_oc8051_int1_n57,
         oc8051_sfr1_oc8051_int1_n56, oc8051_sfr1_oc8051_int1_n55,
         oc8051_sfr1_oc8051_int1_n54, oc8051_sfr1_oc8051_int1_n53,
         oc8051_sfr1_oc8051_int1_n52, oc8051_sfr1_oc8051_int1_n51,
         oc8051_sfr1_oc8051_int1_n50, oc8051_sfr1_oc8051_int1_n49,
         oc8051_sfr1_oc8051_int1_n48, oc8051_sfr1_oc8051_int1_n47,
         oc8051_sfr1_oc8051_int1_n46, oc8051_sfr1_oc8051_int1_n45,
         oc8051_sfr1_oc8051_int1_n44, oc8051_sfr1_oc8051_int1_n43,
         oc8051_sfr1_oc8051_int1_n42, oc8051_sfr1_oc8051_int1_n41,
         oc8051_sfr1_oc8051_int1_n40, oc8051_sfr1_oc8051_int1_n39,
         oc8051_sfr1_oc8051_int1_n38, oc8051_sfr1_oc8051_int1_n37,
         oc8051_sfr1_oc8051_int1_n36, oc8051_sfr1_oc8051_int1_n35,
         oc8051_sfr1_oc8051_int1_n34, oc8051_sfr1_oc8051_int1_n33,
         oc8051_sfr1_oc8051_int1_n32, oc8051_sfr1_oc8051_int1_n31,
         oc8051_sfr1_oc8051_int1_n30, oc8051_sfr1_oc8051_int1_n29,
         oc8051_sfr1_oc8051_int1_n28, oc8051_sfr1_oc8051_int1_n27,
         oc8051_sfr1_oc8051_int1_n26, oc8051_sfr1_oc8051_int1_n25,
         oc8051_sfr1_oc8051_int1_n24, oc8051_sfr1_oc8051_int1_n23,
         oc8051_sfr1_oc8051_int1_n22, oc8051_sfr1_oc8051_int1_n21,
         oc8051_sfr1_oc8051_int1_n20, oc8051_sfr1_oc8051_int1_n19,
         oc8051_sfr1_oc8051_int1_n18, oc8051_sfr1_oc8051_int1_n17,
         oc8051_sfr1_oc8051_int1_n16, oc8051_sfr1_oc8051_int1_n15,
         oc8051_sfr1_oc8051_int1_n14, oc8051_sfr1_oc8051_int1_n13,
         oc8051_sfr1_oc8051_int1_n12, oc8051_sfr1_oc8051_int1_n3,
         oc8051_sfr1_oc8051_int1_n2, oc8051_sfr1_oc8051_int1_int_vec_2_,
         oc8051_sfr1_oc8051_int1_n265, oc8051_sfr1_oc8051_int1_n264,
         oc8051_sfr1_oc8051_int1_n263, oc8051_sfr1_oc8051_int1_n262,
         oc8051_sfr1_oc8051_int1_n261, oc8051_sfr1_oc8051_int1_n260,
         oc8051_sfr1_oc8051_int1_n259, oc8051_sfr1_oc8051_int1_n258,
         oc8051_sfr1_oc8051_int1_n257, oc8051_sfr1_oc8051_int1_n256,
         oc8051_sfr1_oc8051_int1_n255, oc8051_sfr1_oc8051_int1_n254,
         oc8051_sfr1_oc8051_int1_n253, oc8051_sfr1_oc8051_int1_n252,
         oc8051_sfr1_oc8051_int1_n251, oc8051_sfr1_oc8051_int1_n250,
         oc8051_sfr1_oc8051_int1_n249, oc8051_sfr1_oc8051_int1_n248,
         oc8051_sfr1_oc8051_int1_n247, oc8051_sfr1_oc8051_int1_n246,
         oc8051_sfr1_oc8051_int1_n245, oc8051_sfr1_oc8051_int1_n244,
         oc8051_sfr1_oc8051_int1_n243, oc8051_sfr1_oc8051_int1_n242,
         oc8051_sfr1_oc8051_int1_n241, oc8051_sfr1_oc8051_int1_n240,
         oc8051_sfr1_oc8051_int1_n239, oc8051_sfr1_oc8051_int1_n238,
         oc8051_sfr1_oc8051_int1_n237, oc8051_sfr1_oc8051_int1_n236,
         oc8051_sfr1_oc8051_int1_n235, oc8051_sfr1_oc8051_int1_n234,
         oc8051_sfr1_oc8051_int1_n233, oc8051_sfr1_oc8051_int1_n232,
         oc8051_sfr1_oc8051_int1_n231, oc8051_sfr1_oc8051_int1_n230,
         oc8051_sfr1_oc8051_int1_n229, oc8051_sfr1_oc8051_int1_n228,
         oc8051_sfr1_oc8051_int1_n227, oc8051_sfr1_oc8051_int1_n226,
         oc8051_sfr1_oc8051_int1_n11, oc8051_sfr1_oc8051_int1_n10,
         oc8051_sfr1_oc8051_int1_n9, oc8051_sfr1_oc8051_int1_n8,
         oc8051_sfr1_oc8051_int1_n7, oc8051_sfr1_oc8051_int1_n6,
         oc8051_sfr1_oc8051_int1_n5, oc8051_sfr1_oc8051_int1_n4,
         oc8051_sfr1_oc8051_int1_ie1_buff, oc8051_sfr1_oc8051_int1_ie0_buff,
         oc8051_sfr1_oc8051_int1_tf0_buff, oc8051_sfr1_oc8051_int1_tf1_buff,
         oc8051_sfr1_oc8051_int1_int_lev_0__0_,
         oc8051_sfr1_oc8051_int1_int_lev_1__0_,
         oc8051_sfr1_oc8051_int1_int_dept_0_,
         oc8051_sfr1_oc8051_int1_int_dept_1_,
         oc8051_sfr1_oc8051_int1_isrc_0__0_,
         oc8051_sfr1_oc8051_int1_isrc_0__1_,
         oc8051_sfr1_oc8051_int1_isrc_1__0_,
         oc8051_sfr1_oc8051_int1_isrc_1__1_, oc8051_sfr1_oc8051_int1_int_proc,
         oc8051_sfr1_oc8051_tc1_n164, oc8051_sfr1_oc8051_tc1_n163,
         oc8051_sfr1_oc8051_tc1_n162, oc8051_sfr1_oc8051_tc1_n161,
         oc8051_sfr1_oc8051_tc1_n160, oc8051_sfr1_oc8051_tc1_n159,
         oc8051_sfr1_oc8051_tc1_n158, oc8051_sfr1_oc8051_tc1_n157,
         oc8051_sfr1_oc8051_tc1_n156, oc8051_sfr1_oc8051_tc1_n155,
         oc8051_sfr1_oc8051_tc1_n154, oc8051_sfr1_oc8051_tc1_n153,
         oc8051_sfr1_oc8051_tc1_n152, oc8051_sfr1_oc8051_tc1_n151,
         oc8051_sfr1_oc8051_tc1_n150, oc8051_sfr1_oc8051_tc1_n149,
         oc8051_sfr1_oc8051_tc1_n148, oc8051_sfr1_oc8051_tc1_n147,
         oc8051_sfr1_oc8051_tc1_n146, oc8051_sfr1_oc8051_tc1_n145,
         oc8051_sfr1_oc8051_tc1_n144, oc8051_sfr1_oc8051_tc1_n143,
         oc8051_sfr1_oc8051_tc1_n142, oc8051_sfr1_oc8051_tc1_n141,
         oc8051_sfr1_oc8051_tc1_n140, oc8051_sfr1_oc8051_tc1_n139,
         oc8051_sfr1_oc8051_tc1_n138, oc8051_sfr1_oc8051_tc1_n137,
         oc8051_sfr1_oc8051_tc1_n136, oc8051_sfr1_oc8051_tc1_n135,
         oc8051_sfr1_oc8051_tc1_n134, oc8051_sfr1_oc8051_tc1_n133,
         oc8051_sfr1_oc8051_tc1_n132, oc8051_sfr1_oc8051_tc1_n131,
         oc8051_sfr1_oc8051_tc1_n130, oc8051_sfr1_oc8051_tc1_n129,
         oc8051_sfr1_oc8051_tc1_n128, oc8051_sfr1_oc8051_tc1_n127,
         oc8051_sfr1_oc8051_tc1_n126, oc8051_sfr1_oc8051_tc1_n125,
         oc8051_sfr1_oc8051_tc1_n124, oc8051_sfr1_oc8051_tc1_n123,
         oc8051_sfr1_oc8051_tc1_n122, oc8051_sfr1_oc8051_tc1_n121,
         oc8051_sfr1_oc8051_tc1_n120, oc8051_sfr1_oc8051_tc1_n119,
         oc8051_sfr1_oc8051_tc1_n118, oc8051_sfr1_oc8051_tc1_n117,
         oc8051_sfr1_oc8051_tc1_n116, oc8051_sfr1_oc8051_tc1_n115,
         oc8051_sfr1_oc8051_tc1_n114, oc8051_sfr1_oc8051_tc1_n113,
         oc8051_sfr1_oc8051_tc1_n112, oc8051_sfr1_oc8051_tc1_n111,
         oc8051_sfr1_oc8051_tc1_n110, oc8051_sfr1_oc8051_tc1_n109,
         oc8051_sfr1_oc8051_tc1_n108, oc8051_sfr1_oc8051_tc1_n107,
         oc8051_sfr1_oc8051_tc1_n106, oc8051_sfr1_oc8051_tc1_n105,
         oc8051_sfr1_oc8051_tc1_n104, oc8051_sfr1_oc8051_tc1_n103,
         oc8051_sfr1_oc8051_tc1_n102, oc8051_sfr1_oc8051_tc1_n101,
         oc8051_sfr1_oc8051_tc1_n100, oc8051_sfr1_oc8051_tc1_n99,
         oc8051_sfr1_oc8051_tc1_n98, oc8051_sfr1_oc8051_tc1_n97,
         oc8051_sfr1_oc8051_tc1_n96, oc8051_sfr1_oc8051_tc1_n95,
         oc8051_sfr1_oc8051_tc1_n94, oc8051_sfr1_oc8051_tc1_n93,
         oc8051_sfr1_oc8051_tc1_n92, oc8051_sfr1_oc8051_tc1_n91,
         oc8051_sfr1_oc8051_tc1_n90, oc8051_sfr1_oc8051_tc1_n89,
         oc8051_sfr1_oc8051_tc1_n88, oc8051_sfr1_oc8051_tc1_n87,
         oc8051_sfr1_oc8051_tc1_n86, oc8051_sfr1_oc8051_tc1_n85,
         oc8051_sfr1_oc8051_tc1_n84, oc8051_sfr1_oc8051_tc1_n83,
         oc8051_sfr1_oc8051_tc1_n82, oc8051_sfr1_oc8051_tc1_n81,
         oc8051_sfr1_oc8051_tc1_n80, oc8051_sfr1_oc8051_tc1_n79,
         oc8051_sfr1_oc8051_tc1_n78, oc8051_sfr1_oc8051_tc1_n77,
         oc8051_sfr1_oc8051_tc1_n76, oc8051_sfr1_oc8051_tc1_n75,
         oc8051_sfr1_oc8051_tc1_n74, oc8051_sfr1_oc8051_tc1_n73,
         oc8051_sfr1_oc8051_tc1_n72, oc8051_sfr1_oc8051_tc1_n71,
         oc8051_sfr1_oc8051_tc1_n70, oc8051_sfr1_oc8051_tc1_n69,
         oc8051_sfr1_oc8051_tc1_n68, oc8051_sfr1_oc8051_tc1_n67,
         oc8051_sfr1_oc8051_tc1_n66, oc8051_sfr1_oc8051_tc1_n65,
         oc8051_sfr1_oc8051_tc1_n64, oc8051_sfr1_oc8051_tc1_n63,
         oc8051_sfr1_oc8051_tc1_n62, oc8051_sfr1_oc8051_tc1_n61,
         oc8051_sfr1_oc8051_tc1_n60, oc8051_sfr1_oc8051_tc1_n59,
         oc8051_sfr1_oc8051_tc1_n58, oc8051_sfr1_oc8051_tc1_n57,
         oc8051_sfr1_oc8051_tc1_n56, oc8051_sfr1_oc8051_tc1_n55,
         oc8051_sfr1_oc8051_tc1_n54, oc8051_sfr1_oc8051_tc1_n53,
         oc8051_sfr1_oc8051_tc1_n52, oc8051_sfr1_oc8051_tc1_n51,
         oc8051_sfr1_oc8051_tc1_n50, oc8051_sfr1_oc8051_tc1_n49,
         oc8051_sfr1_oc8051_tc1_n48, oc8051_sfr1_oc8051_tc1_n47,
         oc8051_sfr1_oc8051_tc1_n46, oc8051_sfr1_oc8051_tc1_n45,
         oc8051_sfr1_oc8051_tc1_n44, oc8051_sfr1_oc8051_tc1_n43,
         oc8051_sfr1_oc8051_tc1_n42, oc8051_sfr1_oc8051_tc1_n41,
         oc8051_sfr1_oc8051_tc1_n40, oc8051_sfr1_oc8051_tc1_n39,
         oc8051_sfr1_oc8051_tc1_n38, oc8051_sfr1_oc8051_tc1_n37,
         oc8051_sfr1_oc8051_tc1_n36, oc8051_sfr1_oc8051_tc1_n35,
         oc8051_sfr1_oc8051_tc1_n34, oc8051_sfr1_oc8051_tc1_n33,
         oc8051_sfr1_oc8051_tc1_n32, oc8051_sfr1_oc8051_tc1_n31,
         oc8051_sfr1_oc8051_tc1_n30, oc8051_sfr1_oc8051_tc1_n29,
         oc8051_sfr1_oc8051_tc1_n28, oc8051_sfr1_oc8051_tc1_n27,
         oc8051_sfr1_oc8051_tc1_n26, oc8051_sfr1_oc8051_tc1_n25,
         oc8051_sfr1_oc8051_tc1_n24, oc8051_sfr1_oc8051_tc1_n23,
         oc8051_sfr1_oc8051_tc1_n22, oc8051_sfr1_oc8051_tc1_n21,
         oc8051_sfr1_oc8051_tc1_n20, oc8051_sfr1_oc8051_tc1_n19,
         oc8051_sfr1_oc8051_tc1_n18, oc8051_sfr1_oc8051_tc1_n17,
         oc8051_sfr1_oc8051_tc1_n16, oc8051_sfr1_oc8051_tc1_n15,
         oc8051_sfr1_oc8051_tc1_n14, oc8051_sfr1_oc8051_tc1_n13,
         oc8051_sfr1_oc8051_tc1_n12, oc8051_sfr1_oc8051_tc1_n11,
         oc8051_sfr1_oc8051_tc1_n10, oc8051_sfr1_oc8051_tc1_n9,
         oc8051_sfr1_oc8051_tc1_n8, oc8051_sfr1_oc8051_tc1_n7,
         oc8051_sfr1_oc8051_tc1_n6, oc8051_sfr1_oc8051_tc1_n4,
         oc8051_sfr1_oc8051_tc1_n3, oc8051_sfr1_oc8051_tc1_n2,
         oc8051_sfr1_oc8051_tc1_n1, oc8051_sfr1_oc8051_tc1_n268,
         oc8051_sfr1_oc8051_tc1_n267, oc8051_sfr1_oc8051_tc1_n266,
         oc8051_sfr1_oc8051_tc1_n265, oc8051_sfr1_oc8051_tc1_n264,
         oc8051_sfr1_oc8051_tc1_n263, oc8051_sfr1_oc8051_tc1_n262,
         oc8051_sfr1_oc8051_tc1_n261, oc8051_sfr1_oc8051_tc1_n260,
         oc8051_sfr1_oc8051_tc1_n259, oc8051_sfr1_oc8051_tc1_n258,
         oc8051_sfr1_oc8051_tc1_n257, oc8051_sfr1_oc8051_tc1_n256,
         oc8051_sfr1_oc8051_tc1_n255, oc8051_sfr1_oc8051_tc1_n254,
         oc8051_sfr1_oc8051_tc1_n253, oc8051_sfr1_oc8051_tc1_n252,
         oc8051_sfr1_oc8051_tc1_n251, oc8051_sfr1_oc8051_tc1_n250,
         oc8051_sfr1_oc8051_tc1_n249, oc8051_sfr1_oc8051_tc1_n248,
         oc8051_sfr1_oc8051_tc1_n247, oc8051_sfr1_oc8051_tc1_n246,
         oc8051_sfr1_oc8051_tc1_n245, oc8051_sfr1_oc8051_tc1_n244,
         oc8051_sfr1_oc8051_tc1_n243, oc8051_sfr1_oc8051_tc1_n242,
         oc8051_sfr1_oc8051_tc1_n241, oc8051_sfr1_oc8051_tc1_n240,
         oc8051_sfr1_oc8051_tc1_n239, oc8051_sfr1_oc8051_tc1_n238,
         oc8051_sfr1_oc8051_tc1_n237, oc8051_sfr1_oc8051_tc1_n236,
         oc8051_sfr1_oc8051_tc1_n235, oc8051_sfr1_oc8051_tc1_n234,
         oc8051_sfr1_oc8051_tc1_n233, oc8051_sfr1_oc8051_tc1_n232,
         oc8051_sfr1_oc8051_tc1_n231, oc8051_sfr1_oc8051_tc1_n230,
         oc8051_sfr1_oc8051_tc1_n229, oc8051_sfr1_oc8051_tc1_n228,
         oc8051_sfr1_oc8051_tc1_n227, oc8051_sfr1_oc8051_tc1_n226,
         oc8051_sfr1_oc8051_tc1_n225, oc8051_sfr1_oc8051_tc1_n224,
         oc8051_sfr1_oc8051_tc1_n223, oc8051_sfr1_oc8051_tc1_n222,
         oc8051_sfr1_oc8051_tc1_n221, oc8051_sfr1_oc8051_tc1_n220,
         oc8051_sfr1_oc8051_tc1_n219, oc8051_sfr1_oc8051_tc1_n218,
         oc8051_sfr1_oc8051_tc1_n217, oc8051_sfr1_oc8051_tc1_n216,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_15, oc8051_sfr1_oc8051_tc1_u3_u8_z_14,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_13, oc8051_sfr1_oc8051_tc1_u3_u8_z_12,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_11, oc8051_sfr1_oc8051_tc1_u3_u8_z_10,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_9, oc8051_sfr1_oc8051_tc1_u3_u8_z_8,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_7, oc8051_sfr1_oc8051_tc1_u3_u8_z_6,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_5, oc8051_sfr1_oc8051_tc1_u3_u1_z_15,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_14, oc8051_sfr1_oc8051_tc1_u3_u1_z_13,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_12, oc8051_sfr1_oc8051_tc1_u3_u1_z_11,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_10, oc8051_sfr1_oc8051_tc1_u3_u1_z_9,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_8, oc8051_sfr1_oc8051_tc1_u3_u1_z_7,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_6, oc8051_sfr1_oc8051_tc1_u3_u1_z_5,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_4, oc8051_sfr1_oc8051_tc1_u3_u1_z_3,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_2, oc8051_sfr1_oc8051_tc1_u3_u1_z_1,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_0, oc8051_sfr1_oc8051_tc1_n5,
         oc8051_sfr1_oc8051_tc1_n203, oc8051_sfr1_oc8051_tc1_n202,
         oc8051_sfr1_oc8051_tc1_n201, oc8051_sfr1_oc8051_tc1_n200,
         oc8051_sfr1_oc8051_tc1_n199, oc8051_sfr1_oc8051_tc1_n198,
         oc8051_sfr1_oc8051_tc1_n197, oc8051_sfr1_oc8051_tc1_n196,
         oc8051_sfr1_oc8051_tc1_n192, oc8051_sfr1_oc8051_tc1_n191,
         oc8051_sfr1_oc8051_tc1_n190, oc8051_sfr1_oc8051_tc1_n174,
         oc8051_sfr1_oc8051_tc1_n173, oc8051_sfr1_oc8051_tc1_n172,
         oc8051_sfr1_oc8051_tc1_n171, oc8051_sfr1_oc8051_tc1_n170,
         oc8051_sfr1_oc8051_tc1_n169, oc8051_sfr1_oc8051_tc1_n168,
         oc8051_sfr1_oc8051_tc1_n167, oc8051_sfr1_oc8051_tc1_n166,
         oc8051_sfr1_oc8051_tc1_n165, oc8051_sfr1_oc8051_tc1_n1640,
         oc8051_sfr1_oc8051_tc1_n1630, oc8051_sfr1_oc8051_tc1_n1620,
         oc8051_sfr1_oc8051_tc1_n1610, oc8051_sfr1_oc8051_tc1_n920,
         oc8051_sfr1_oc8051_tc1_n910, oc8051_sfr1_oc8051_tc1_n900,
         oc8051_sfr1_oc8051_tc1_n890, oc8051_sfr1_oc8051_tc1_n880,
         oc8051_sfr1_oc8051_tc1_n870, oc8051_sfr1_oc8051_tc1_n860,
         oc8051_sfr1_oc8051_tc1_n850, oc8051_sfr1_oc8051_tc1_n840,
         oc8051_sfr1_oc8051_tc1_n630, oc8051_sfr1_oc8051_tc1_n620,
         oc8051_sfr1_oc8051_tc1_n610, oc8051_sfr1_oc8051_tc1_n600,
         oc8051_sfr1_oc8051_tc1_n590, oc8051_sfr1_oc8051_tc1_n580,
         oc8051_sfr1_oc8051_tc1_n570, oc8051_sfr1_oc8051_tc1_n560,
         oc8051_sfr1_oc8051_tc1_n550, oc8051_sfr1_oc8051_tc1_n540,
         oc8051_sfr1_oc8051_tc1_n530, oc8051_sfr1_oc8051_tc1_n520,
         oc8051_sfr1_oc8051_tc1_n510, oc8051_sfr1_oc8051_tc1_n500,
         oc8051_sfr1_oc8051_tc1_n490, oc8051_sfr1_oc8051_tc1_n480,
         oc8051_sfr1_oc8051_tc1_n470, oc8051_sfr1_oc8051_tc1_t1_buff,
         oc8051_sfr1_oc8051_tc1_t0_buff, oc8051_sfr1_oc8051_tc21_n139,
         oc8051_sfr1_oc8051_tc21_n138, oc8051_sfr1_oc8051_tc21_n137,
         oc8051_sfr1_oc8051_tc21_n136, oc8051_sfr1_oc8051_tc21_n135,
         oc8051_sfr1_oc8051_tc21_n134, oc8051_sfr1_oc8051_tc21_n133,
         oc8051_sfr1_oc8051_tc21_n132, oc8051_sfr1_oc8051_tc21_n131,
         oc8051_sfr1_oc8051_tc21_n130, oc8051_sfr1_oc8051_tc21_n129,
         oc8051_sfr1_oc8051_tc21_n128, oc8051_sfr1_oc8051_tc21_n127,
         oc8051_sfr1_oc8051_tc21_n126, oc8051_sfr1_oc8051_tc21_n125,
         oc8051_sfr1_oc8051_tc21_n124, oc8051_sfr1_oc8051_tc21_n123,
         oc8051_sfr1_oc8051_tc21_n122, oc8051_sfr1_oc8051_tc21_n121,
         oc8051_sfr1_oc8051_tc21_n120, oc8051_sfr1_oc8051_tc21_n119,
         oc8051_sfr1_oc8051_tc21_n118, oc8051_sfr1_oc8051_tc21_n117,
         oc8051_sfr1_oc8051_tc21_n116, oc8051_sfr1_oc8051_tc21_n115,
         oc8051_sfr1_oc8051_tc21_n114, oc8051_sfr1_oc8051_tc21_n113,
         oc8051_sfr1_oc8051_tc21_n112, oc8051_sfr1_oc8051_tc21_n111,
         oc8051_sfr1_oc8051_tc21_n110, oc8051_sfr1_oc8051_tc21_n109,
         oc8051_sfr1_oc8051_tc21_n108, oc8051_sfr1_oc8051_tc21_n107,
         oc8051_sfr1_oc8051_tc21_n106, oc8051_sfr1_oc8051_tc21_n105,
         oc8051_sfr1_oc8051_tc21_n104, oc8051_sfr1_oc8051_tc21_n103,
         oc8051_sfr1_oc8051_tc21_n102, oc8051_sfr1_oc8051_tc21_n101,
         oc8051_sfr1_oc8051_tc21_n100, oc8051_sfr1_oc8051_tc21_n99,
         oc8051_sfr1_oc8051_tc21_n98, oc8051_sfr1_oc8051_tc21_n97,
         oc8051_sfr1_oc8051_tc21_n96, oc8051_sfr1_oc8051_tc21_n95,
         oc8051_sfr1_oc8051_tc21_n94, oc8051_sfr1_oc8051_tc21_n93,
         oc8051_sfr1_oc8051_tc21_n92, oc8051_sfr1_oc8051_tc21_n91,
         oc8051_sfr1_oc8051_tc21_n90, oc8051_sfr1_oc8051_tc21_n89,
         oc8051_sfr1_oc8051_tc21_n88, oc8051_sfr1_oc8051_tc21_n87,
         oc8051_sfr1_oc8051_tc21_n86, oc8051_sfr1_oc8051_tc21_n85,
         oc8051_sfr1_oc8051_tc21_n84, oc8051_sfr1_oc8051_tc21_n83,
         oc8051_sfr1_oc8051_tc21_n82, oc8051_sfr1_oc8051_tc21_n81,
         oc8051_sfr1_oc8051_tc21_n80, oc8051_sfr1_oc8051_tc21_n79,
         oc8051_sfr1_oc8051_tc21_n78, oc8051_sfr1_oc8051_tc21_n77,
         oc8051_sfr1_oc8051_tc21_n76, oc8051_sfr1_oc8051_tc21_n75,
         oc8051_sfr1_oc8051_tc21_n74, oc8051_sfr1_oc8051_tc21_n73,
         oc8051_sfr1_oc8051_tc21_n72, oc8051_sfr1_oc8051_tc21_n71,
         oc8051_sfr1_oc8051_tc21_n70, oc8051_sfr1_oc8051_tc21_n69,
         oc8051_sfr1_oc8051_tc21_n68, oc8051_sfr1_oc8051_tc21_n67,
         oc8051_sfr1_oc8051_tc21_n66, oc8051_sfr1_oc8051_tc21_n65,
         oc8051_sfr1_oc8051_tc21_n64, oc8051_sfr1_oc8051_tc21_n63,
         oc8051_sfr1_oc8051_tc21_n62, oc8051_sfr1_oc8051_tc21_n61,
         oc8051_sfr1_oc8051_tc21_n60, oc8051_sfr1_oc8051_tc21_n59,
         oc8051_sfr1_oc8051_tc21_n58, oc8051_sfr1_oc8051_tc21_n57,
         oc8051_sfr1_oc8051_tc21_n56, oc8051_sfr1_oc8051_tc21_n55,
         oc8051_sfr1_oc8051_tc21_n54, oc8051_sfr1_oc8051_tc21_n53,
         oc8051_sfr1_oc8051_tc21_n52, oc8051_sfr1_oc8051_tc21_n51,
         oc8051_sfr1_oc8051_tc21_n50, oc8051_sfr1_oc8051_tc21_n49,
         oc8051_sfr1_oc8051_tc21_n48, oc8051_sfr1_oc8051_tc21_n47,
         oc8051_sfr1_oc8051_tc21_n46, oc8051_sfr1_oc8051_tc21_n45,
         oc8051_sfr1_oc8051_tc21_n44, oc8051_sfr1_oc8051_tc21_n43,
         oc8051_sfr1_oc8051_tc21_n42, oc8051_sfr1_oc8051_tc21_n41,
         oc8051_sfr1_oc8051_tc21_n40, oc8051_sfr1_oc8051_tc21_n39,
         oc8051_sfr1_oc8051_tc21_n38, oc8051_sfr1_oc8051_tc21_n37,
         oc8051_sfr1_oc8051_tc21_n36, oc8051_sfr1_oc8051_tc21_n35,
         oc8051_sfr1_oc8051_tc21_n34, oc8051_sfr1_oc8051_tc21_n33,
         oc8051_sfr1_oc8051_tc21_n32, oc8051_sfr1_oc8051_tc21_n31,
         oc8051_sfr1_oc8051_tc21_n30, oc8051_sfr1_oc8051_tc21_n29,
         oc8051_sfr1_oc8051_tc21_n28, oc8051_sfr1_oc8051_tc21_n27,
         oc8051_sfr1_oc8051_tc21_n26, oc8051_sfr1_oc8051_tc21_n25,
         oc8051_sfr1_oc8051_tc21_n24, oc8051_sfr1_oc8051_tc21_n23,
         oc8051_sfr1_oc8051_tc21_n22, oc8051_sfr1_oc8051_tc21_n21,
         oc8051_sfr1_oc8051_tc21_n20, oc8051_sfr1_oc8051_tc21_n19,
         oc8051_sfr1_oc8051_tc21_n18, oc8051_sfr1_oc8051_tc21_n17,
         oc8051_sfr1_oc8051_tc21_n16, oc8051_sfr1_oc8051_tc21_n15,
         oc8051_sfr1_oc8051_tc21_n14, oc8051_sfr1_oc8051_tc21_n13,
         oc8051_sfr1_oc8051_tc21_n12, oc8051_sfr1_oc8051_tc21_n11,
         oc8051_sfr1_oc8051_tc21_n10, oc8051_sfr1_oc8051_tc21_n9,
         oc8051_sfr1_oc8051_tc21_n4, oc8051_sfr1_oc8051_tc21_n3,
         oc8051_sfr1_oc8051_tc21_n2, oc8051_sfr1_oc8051_tc21_n191,
         oc8051_sfr1_oc8051_tc21_n190, oc8051_sfr1_oc8051_tc21_n189,
         oc8051_sfr1_oc8051_tc21_n188, oc8051_sfr1_oc8051_tc21_n187,
         oc8051_sfr1_oc8051_tc21_n186, oc8051_sfr1_oc8051_tc21_n185,
         oc8051_sfr1_oc8051_tc21_n184, oc8051_sfr1_oc8051_tc21_n183,
         oc8051_sfr1_oc8051_tc21_n182, oc8051_sfr1_oc8051_tc21_n181,
         oc8051_sfr1_oc8051_tc21_n180, oc8051_sfr1_oc8051_tc21_n179,
         oc8051_sfr1_oc8051_tc21_n178, oc8051_sfr1_oc8051_tc21_n177,
         oc8051_sfr1_oc8051_tc21_n176, oc8051_sfr1_oc8051_tc21_n175,
         oc8051_sfr1_oc8051_tc21_n174, oc8051_sfr1_oc8051_tc21_n173,
         oc8051_sfr1_oc8051_tc21_n172, oc8051_sfr1_oc8051_tc21_n171,
         oc8051_sfr1_oc8051_tc21_n170, oc8051_sfr1_oc8051_tc21_n169,
         oc8051_sfr1_oc8051_tc21_n168, oc8051_sfr1_oc8051_tc21_n167,
         oc8051_sfr1_oc8051_tc21_n166, oc8051_sfr1_oc8051_tc21_n165,
         oc8051_sfr1_oc8051_tc21_n164, oc8051_sfr1_oc8051_tc21_n163,
         oc8051_sfr1_oc8051_tc21_n162, oc8051_sfr1_oc8051_tc21_n161,
         oc8051_sfr1_oc8051_tc21_n160, oc8051_sfr1_oc8051_tc21_n159,
         oc8051_sfr1_oc8051_tc21_n158, oc8051_sfr1_oc8051_tc21_n157,
         oc8051_sfr1_oc8051_tc21_n156, oc8051_sfr1_oc8051_tc21_n155,
         oc8051_sfr1_oc8051_tc21_n154, oc8051_sfr1_oc8051_tc21_n153,
         oc8051_sfr1_oc8051_tc21_n152, oc8051_sfr1_oc8051_tc21_n151,
         oc8051_sfr1_oc8051_tc21_n150, oc8051_sfr1_oc8051_tc21_n8,
         oc8051_sfr1_oc8051_tc21_n7, oc8051_sfr1_oc8051_tc21_n6,
         oc8051_sfr1_oc8051_tc21_n5, oc8051_sfr1_oc8051_tc21_n1,
         oc8051_sfr1_oc8051_tc21_n220, oc8051_sfr1_oc8051_tc21_t2_r,
         oc8051_sfr1_oc8051_tc21_n217, oc8051_sfr1_oc8051_tc21_t2ex_r,
         oc8051_sfr1_oc8051_tc21_n850, oc8051_sfr1_oc8051_tc21_n840,
         oc8051_sfr1_oc8051_tc21_n830, oc8051_sfr1_oc8051_tc21_n820,
         oc8051_sfr1_oc8051_tc21_n810, oc8051_sfr1_oc8051_tc21_n800,
         oc8051_sfr1_oc8051_tc21_n790, oc8051_sfr1_oc8051_tc21_n780,
         oc8051_sfr1_oc8051_tc21_n770, oc8051_sfr1_oc8051_tc21_n760,
         oc8051_sfr1_oc8051_tc21_n750, oc8051_sfr1_oc8051_tc21_n740,
         oc8051_sfr1_oc8051_tc21_n730, oc8051_sfr1_oc8051_tc21_n720,
         oc8051_sfr1_oc8051_tc21_n710, oc8051_sfr1_oc8051_tc21_n700,
         oc8051_sfr1_oc8051_tc21_n690, oc8051_sfr1_oc8051_tc21_tc2_event,
         oc8051_sfr1_oc8051_tc21_neg_trans, oc8051_sfr1_oc8051_tc21_tf2_set;
  wire   [7:0] op1_n;
  wire   [2:0] op1_cur;
  wire   [2:0] ram_rd_sel;
  wire   [2:0] ram_wr_sel;
  wire   [2:0] src_sel1;
  wire   [1:0] src_sel2;
  wire   [3:0] alu_op;
  wire   [1:0] psw_set;
  wire   [1:0] cy_sel;
  wire   [2:0] pc_wr_sel;
  wire   [1:0] comp_sel;
  wire   [1:0] wr_sfr;
  wire   [2:0] mem_act;
  wire   [7:0] src1;
  wire   [7:0] src2;
  wire   [7:0] src3;
  wire   [7:0] des_acc;
  wire   [7:0] sub_result;
  wire   [7:0] des2;
  wire   [7:0] rd_addr;
  wire   [7:0] ram_data;
  wire   [7:0] wr_addr;
  wire   [7:0] wr_dat;
  wire   [7:0] acc;
  wire   [7:0] ram_out;
  wire   [15:0] pc;
  wire   [7:0] op2_n;
  wire   [7:0] op3_n;
  wire   [7:0] dptr_hi;
  wire   [7:0] dptr_lo;
  wire   [7:0] ri;
  wire   [1:0] bank_sel;
  wire   [7:0] sfr_out;
  wire   [5:0] int_src;
  wire   [7:0] sp_w;
  wire   [7:0] sp;
  wire   [2:0] oc8051_decoder1_ram_rd_sel_r;
  wire   [7:0] oc8051_decoder1_op;
  wire   [1:3] oc8051_alu1_add_1_root_add_173_2_carry;
  wire   [0:3] oc8051_alu1_sub_1_root_sub_189_2_b_not;
  wire   [7:0] oc8051_alu1_des_acc_1;
  wire   [15:0] oc8051_alu1_dec;
  wire   [15:0] oc8051_alu1_inc;
  wire   [7:0] oc8051_alu1_divsrc2;
  wire   [7:0] oc8051_alu1_divsrc1;
  wire   [7:0] oc8051_alu1_mulsrc2;
  wire   [7:0] oc8051_alu1_mulsrc1;
  wire   [13:0] oc8051_alu1_oc8051_mul1_tmp_mul;
  wire   [9:2] oc8051_alu1_oc8051_mul1_mul_result1;
  wire   [8:0] oc8051_alu1_oc8051_div1_sub0;
  wire   [8:0] oc8051_alu1_oc8051_div1_sub1;
  wire   [7:0] oc8051_alu1_oc8051_div1_tmp_rem;
  wire   [8:2] oc8051_alu1_oc8051_div1_sub_98_carry;
  wire   [7:1] oc8051_alu1_oc8051_div1_sub_94_b_not;
  wire   [8:2] oc8051_alu1_oc8051_div1_sub_94_carry;
  wire   [15:2] oc8051_alu1_add_204_carry;
  wire   [7:0] oc8051_ram_top1_wr_data_m;
  wire   [7:0] oc8051_ram_top1_rd_data_m;
  wire   [7:0] oc8051_ram_top1_wr_data_r;
  wire   [7:0] oc8051_alu_src_sel1_op3_r;
  wire   [7:0] oc8051_alu_src_sel1_op1_r;
  wire   [7:0] oc8051_memory_interface1_pcs_result;
  wire   [7:0] oc8051_memory_interface1_op2_buff;
  wire   [7:0] oc8051_memory_interface1_op3_buff;
  wire   [7:0] oc8051_memory_interface1_op3;
  wire   [7:0] oc8051_memory_interface1_op2;
  wire   [7:0] oc8051_memory_interface1_imm2_r;
  wire   [7:0] oc8051_memory_interface1_imm_r;
  wire   [7:0] oc8051_memory_interface1_ri_r;
  wire   [4:0] oc8051_memory_interface1_rn_r;
  wire   [7:0] oc8051_sfr1_rcap2h;
  wire   [7:0] oc8051_sfr1_rcap2l;
  wire   [7:0] oc8051_sfr1_th2;
  wire   [7:0] oc8051_sfr1_tl2;
  wire   [7:0] oc8051_sfr1_th1;
  wire   [7:0] oc8051_sfr1_tl1;
  wire   [7:0] oc8051_sfr1_th0;
  wire   [7:0] oc8051_sfr1_tl0;
  wire   [7:0] oc8051_sfr1_tmod;
  wire   [7:0] oc8051_sfr1_sbuf;
  wire   [7:0] oc8051_sfr1_pcon;
  wire   [7:0] oc8051_sfr1_oc8051_sp1_sp_t;
  wire   [7:2] oc8051_sfr1_oc8051_sp1_add_102_s2_carry;
  wire   [15:2] oc8051_sfr1_oc8051_tc1_r372_carry;
  wire   [7:2] oc8051_sfr1_oc8051_tc1_add_220_carry;
  wire   [7:2] oc8051_sfr1_oc8051_tc1_r364_carry;
  wire   [15:2] oc8051_sfr1_oc8051_tc1_r360_carry;
  wire   [15:2] oc8051_sfr1_oc8051_tc21_r320_carry;
  assign wbi_cyc_o = wbi_stb_o;
  assign wbd_stb_o = wbd_cyc_o;

  TIELO_X1M_A12TS u7 ( .Y(n_logic0_) );
  TIEHI_X1M_A12TS u8 ( .Y(wbi_stb_o) );
  NOR2_X0P5A_A12TS u9 ( .A(wr_ind), .B(n2), .Y(n_5_net_) );
  AND2_X0P5M_A12TS u10 ( .A(pc_wr), .B(comp_wait), .Y(n_3_net_) );
  AOI2XB1_X0P5M_A12TS u11 ( .A1N(wr_ind), .A0(wr_addr[7]), .B0(n2), .Y(
        n_0_net_) );
  INV_X0P5B_A12TS u12 ( .A(wr_o), .Y(n2) );
  INV_X0P5B_A12TS oc8051_decoder1_u472 ( .A(oc8051_decoder1_state_1_), .Y(
        oc8051_decoder1_n317) );
  INV_X0P5B_A12TS oc8051_decoder1_u471 ( .A(oc8051_decoder1_state_0_), .Y(
        oc8051_decoder1_n316) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u470 ( .A(oc8051_decoder1_n317), .B(
        oc8051_decoder1_n316), .Y(oc8051_decoder1_n303) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u469 ( .A(oc8051_decoder1_n303), .B(
        wait_data), .Y(rd) );
  INV_X0P5B_A12TS oc8051_decoder1_u468 ( .A(mem_wait), .Y(oc8051_decoder1_n435) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u467 ( .A(rd), .B(oc8051_decoder1_n435), 
        .Y(oc8051_decoder1_n318) );
  INV_X0P5B_A12TS oc8051_decoder1_u466 ( .A(op1_n[0]), .Y(oc8051_decoder1_n301) );
  OR2_X0P5M_A12TS oc8051_decoder1_u465 ( .A(rd), .B(mem_wait), .Y(
        oc8051_decoder1_n439) );
  INV_X0P5B_A12TS oc8051_decoder1_u464 ( .A(oc8051_decoder1_op[0]), .Y(
        oc8051_decoder1_n302) );
  INV_X0P5B_A12TS oc8051_decoder1_u463 ( .A(op1_n[1]), .Y(oc8051_decoder1_n304) );
  INV_X0P5B_A12TS oc8051_decoder1_u462 ( .A(oc8051_decoder1_op[1]), .Y(
        oc8051_decoder1_n305) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u461 ( .A0(oc8051_decoder1_n318), .A1(
        oc8051_decoder1_n304), .B0(oc8051_decoder1_n439), .B1(
        oc8051_decoder1_n305), .Y(op1_cur[1]) );
  INV_X0P5B_A12TS oc8051_decoder1_u460 ( .A(op1_cur[1]), .Y(
        oc8051_decoder1_n22) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u459 ( .A(op1_cur[0]), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n25) );
  INV_X0P5B_A12TS oc8051_decoder1_u458 ( .A(oc8051_decoder1_op[3]), .Y(
        oc8051_decoder1_n309) );
  INV_X0P5B_A12TS oc8051_decoder1_u457 ( .A(op1_n[3]), .Y(oc8051_decoder1_n308) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u456 ( .A(oc8051_decoder1_n309), .B(
        oc8051_decoder1_n308), .S0(rd), .Y(oc8051_decoder1_n440) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u455 ( .A(oc8051_decoder1_n440), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n69) );
  INV_X0P5B_A12TS oc8051_decoder1_u454 ( .A(op1_n[2]), .Y(oc8051_decoder1_n306) );
  INV_X0P5B_A12TS oc8051_decoder1_u453 ( .A(oc8051_decoder1_op[2]), .Y(
        oc8051_decoder1_n307) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u452 ( .A0(oc8051_decoder1_n318), .A1(
        oc8051_decoder1_n306), .B0(oc8051_decoder1_n439), .B1(
        oc8051_decoder1_n307), .Y(op1_cur[2]) );
  INV_X0P5B_A12TS oc8051_decoder1_u451 ( .A(op1_cur[2]), .Y(
        oc8051_decoder1_n131) );
  INV_X0P5B_A12TS oc8051_decoder1_u450 ( .A(oc8051_decoder1_op[7]), .Y(
        oc8051_decoder1_n315) );
  INV_X0P5B_A12TS oc8051_decoder1_u449 ( .A(op1_n[7]), .Y(oc8051_decoder1_n314) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u448 ( .A(oc8051_decoder1_n315), .B(
        oc8051_decoder1_n314), .S0(rd), .Y(oc8051_decoder1_n438) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u447 ( .A(oc8051_decoder1_n438), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n185) );
  INV_X0P5B_A12TS oc8051_decoder1_u446 ( .A(oc8051_decoder1_n185), .Y(
        oc8051_decoder1_n54) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u445 ( .A(oc8051_decoder1_n69), .B(
        oc8051_decoder1_n131), .C(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n334) );
  INV_X0P5B_A12TS oc8051_decoder1_u444 ( .A(oc8051_decoder1_n334), .Y(
        oc8051_decoder1_n224) );
  AND3_X0P5M_A12TS oc8051_decoder1_u443 ( .A(rd), .B(oc8051_decoder1_n25), .C(
        oc8051_decoder1_n224), .Y(oc8051_decoder1_n432) );
  INV_X0P5B_A12TS oc8051_decoder1_u442 ( .A(oc8051_decoder1_op[4]), .Y(
        oc8051_decoder1_n310) );
  INV_X0P5B_A12TS oc8051_decoder1_u441 ( .A(op1_n[4]), .Y(oc8051_decoder1_n300) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u440 ( .A(oc8051_decoder1_n310), .B(
        oc8051_decoder1_n300), .S0(rd), .Y(oc8051_decoder1_n437) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u439 ( .A(oc8051_decoder1_n437), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n82) );
  INV_X0P5B_A12TS oc8051_decoder1_u438 ( .A(oc8051_decoder1_n82), .Y(
        oc8051_decoder1_n165) );
  INV_X0P5B_A12TS oc8051_decoder1_u437 ( .A(oc8051_decoder1_op[5]), .Y(
        oc8051_decoder1_n312) );
  INV_X0P5B_A12TS oc8051_decoder1_u436 ( .A(op1_n[5]), .Y(oc8051_decoder1_n311) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u435 ( .A(oc8051_decoder1_n312), .B(
        oc8051_decoder1_n311), .S0(rd), .Y(oc8051_decoder1_n436) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u434 ( .A(oc8051_decoder1_n436), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n71) );
  INV_X0P5B_A12TS oc8051_decoder1_u433 ( .A(oc8051_decoder1_n71), .Y(
        oc8051_decoder1_n161) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u432 ( .A(oc8051_decoder1_n165), .B(
        oc8051_decoder1_n161), .Y(oc8051_decoder1_n59) );
  INV_X0P5B_A12TS oc8051_decoder1_u431 ( .A(op1_cur[0]), .Y(
        oc8051_decoder1_n137) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u430 ( .A(oc8051_decoder1_n71), .B(
        oc8051_decoder1_n137), .Y(oc8051_decoder1_n55) );
  INV_X0P5B_A12TS oc8051_decoder1_u429 ( .A(oc8051_decoder1_op[6]), .Y(
        oc8051_decoder1_n313) );
  INV_X0P5B_A12TS oc8051_decoder1_u428 ( .A(op1_n[6]), .Y(oc8051_decoder1_n299) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u427 ( .A(oc8051_decoder1_n313), .B(
        oc8051_decoder1_n299), .S0(rd), .Y(oc8051_decoder1_n434) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u426 ( .A(oc8051_decoder1_n434), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n21) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u425 ( .A(oc8051_decoder1_n21), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n431) );
  INV_X0P5B_A12TS oc8051_decoder1_u424 ( .A(oc8051_decoder1_n21), .Y(
        oc8051_decoder1_n14) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u423 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n275) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u422 ( .A(oc8051_decoder1_n431), .B(
        oc8051_decoder1_n275), .Y(oc8051_decoder1_n141) );
  INV_X0P5B_A12TS oc8051_decoder1_u421 ( .A(oc8051_decoder1_n141), .Y(
        oc8051_decoder1_n118) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u420 ( .A(oc8051_decoder1_n432), .B(
        oc8051_decoder1_n59), .C(oc8051_decoder1_n55), .D(oc8051_decoder1_n118), .Y(oc8051_decoder1_n1804) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u419 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n225) );
  INV_X0P5B_A12TS oc8051_decoder1_u418 ( .A(oc8051_decoder1_n225), .Y(
        oc8051_decoder1_n139) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u417 ( .A0(oc8051_decoder1_n21), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n139), .Y(
        oc8051_decoder1_n433) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u416 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n432), .C0(
        oc8051_decoder1_n433), .Y(oc8051_decoder1_n1805) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u415 ( .A(oc8051_decoder1_n431), .B(
        oc8051_decoder1_n432), .Y(oc8051_decoder1_n1806) );
  INV_X0P5B_A12TS oc8051_decoder1_u414 ( .A(oc8051_decoder1_alu_op_0_), .Y(
        oc8051_decoder1_n124) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u413 ( .A(wait_data), .B(
        oc8051_decoder1_n124), .Y(alu_op[0]) );
  INV_X0P5B_A12TS oc8051_decoder1_u412 ( .A(oc8051_decoder1_alu_op_1_), .Y(
        oc8051_decoder1_n145) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u411 ( .A(wait_data), .B(
        oc8051_decoder1_n145), .Y(alu_op[1]) );
  NOR2B_X0P5M_A12TS oc8051_decoder1_u410 ( .AN(oc8051_decoder1_alu_op_2_), .B(
        wait_data), .Y(alu_op[2]) );
  INV_X0P5B_A12TS oc8051_decoder1_u409 ( .A(oc8051_decoder1_alu_op_3_), .Y(
        oc8051_decoder1_n379) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u408 ( .A(wait_data), .B(
        oc8051_decoder1_n379), .Y(alu_op[3]) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u407 ( .A(op1_cur[1]), .B(
        oc8051_decoder1_n137), .Y(oc8051_decoder1_n193) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u406 ( .A(oc8051_decoder1_n71), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n375) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u405 ( .A(oc8051_decoder1_n375), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n52) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u404 ( .A0(oc8051_decoder1_n161), .A1(
        oc8051_decoder1_n193), .B0(oc8051_decoder1_n52), .Y(
        oc8051_decoder1_n430) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u403 ( .A(op1_cur[1]), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n66) );
  INV_X0P5B_A12TS oc8051_decoder1_u402 ( .A(oc8051_decoder1_n66), .Y(
        oc8051_decoder1_n425) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u401 ( .A(oc8051_decoder1_n69), .B(
        oc8051_decoder1_n131), .Y(oc8051_decoder1_n36) );
  INV_X0P5B_A12TS oc8051_decoder1_u400 ( .A(oc8051_decoder1_n36), .Y(
        oc8051_decoder1_n90) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u399 ( .A(oc8051_decoder1_n425), .B(
        oc8051_decoder1_n90), .Y(oc8051_decoder1_n257) );
  INV_X0P5B_A12TS oc8051_decoder1_u398 ( .A(oc8051_decoder1_n257), .Y(
        oc8051_decoder1_n75) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u397 ( .A(oc8051_decoder1_n75), .B(
        oc8051_decoder1_n137), .Y(oc8051_decoder1_n270) );
  INV_X0P5B_A12TS oc8051_decoder1_u396 ( .A(oc8051_decoder1_n270), .Y(
        oc8051_decoder1_n109) );
  INV_X0P5B_A12TS oc8051_decoder1_u395 ( .A(oc8051_decoder1_n59), .Y(
        oc8051_decoder1_n53) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u394 ( .A(oc8051_decoder1_n53), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n283) );
  INV_X0P5B_A12TS oc8051_decoder1_u393 ( .A(oc8051_decoder1_n283), .Y(
        oc8051_decoder1_n221) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u392 ( .A0(oc8051_decoder1_n224), .A1(
        oc8051_decoder1_n430), .B0(oc8051_decoder1_n109), .B1(
        oc8051_decoder1_n221), .Y(oc8051_decoder1_n428) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u391 ( .A(oc8051_decoder1_n53), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n115) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u390 ( .A(oc8051_decoder1_n137), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n50) );
  INV_X0P5B_A12TS oc8051_decoder1_u389 ( .A(oc8051_decoder1_n50), .Y(
        oc8051_decoder1_n178) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u388 ( .A(oc8051_decoder1_n90), .B(
        oc8051_decoder1_n185), .C(oc8051_decoder1_n178), .Y(
        oc8051_decoder1_n322) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u387 ( .A(oc8051_decoder1_n115), .B(
        oc8051_decoder1_n322), .Y(oc8051_decoder1_n85) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u386 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n58) );
  INV_X0P5B_A12TS oc8051_decoder1_u385 ( .A(oc8051_decoder1_n58), .Y(
        oc8051_decoder1_n42) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u384 ( .A(oc8051_decoder1_n42), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n236) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u383 ( .A(oc8051_decoder1_n236), .B(
        oc8051_decoder1_n322), .Y(oc8051_decoder1_n84) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u382 ( .A(oc8051_decoder1_n85), .B(
        oc8051_decoder1_n84), .Y(oc8051_decoder1_n92) );
  INV_X0P5B_A12TS oc8051_decoder1_u381 ( .A(oc8051_decoder1_n92), .Y(
        oc8051_decoder1_n117) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u380 ( .A(oc8051_decoder1_n165), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n265) );
  INV_X0P5B_A12TS oc8051_decoder1_u379 ( .A(oc8051_decoder1_n265), .Y(
        oc8051_decoder1_n156) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u378 ( .A(oc8051_decoder1_n156), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n226) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u377 ( .A(oc8051_decoder1_n226), .B(
        oc8051_decoder1_n322), .Y(oc8051_decoder1_n83) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u376 ( .A(oc8051_decoder1_n117), .B(
        oc8051_decoder1_n83), .Y(oc8051_decoder1_n112) );
  INV_X0P5B_A12TS oc8051_decoder1_u375 ( .A(wait_data), .Y(
        oc8051_decoder1_n125) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u374 ( .A(oc8051_decoder1_n125), .B(
        oc8051_decoder1_n303), .Y(oc8051_decoder1_n33) );
  INV_X0P5B_A12TS oc8051_decoder1_u373 ( .A(oc8051_decoder1_n33), .Y(
        oc8051_decoder1_n5) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u372 ( .A(oc8051_decoder1_n316), .B(
        oc8051_decoder1_n125), .C(oc8051_decoder1_state_1_), .Y(
        oc8051_decoder1_n30) );
  INV_X0P5B_A12TS oc8051_decoder1_u371 ( .A(oc8051_decoder1_n30), .Y(
        oc8051_decoder1_n111) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u370 ( .A0(oc8051_decoder1_n85), .A1(
        oc8051_decoder1_n83), .B0(oc8051_decoder1_n111), .Y(
        oc8051_decoder1_n429) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u369 ( .A0(oc8051_decoder1_n428), .A1(
        oc8051_decoder1_n112), .B0(oc8051_decoder1_n5), .C0(
        oc8051_decoder1_n429), .Y(bit_addr_o) );
  INV_X0P5B_A12TS oc8051_decoder1_u368 ( .A(oc8051_decoder1_n322), .Y(
        oc8051_decoder1_n427) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u367 ( .A(oc8051_decoder1_n427), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n29) );
  INV_X0P5B_A12TS oc8051_decoder1_u366 ( .A(oc8051_decoder1_n29), .Y(
        oc8051_decoder1_n81) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u365 ( .A(oc8051_decoder1_n111), .B(
        oc8051_decoder1_n81), .Y(comp_sel[0]) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u364 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n156), .Y(oc8051_decoder1_n11) );
  INV_X0P5B_A12TS oc8051_decoder1_u363 ( .A(oc8051_decoder1_n11), .Y(
        oc8051_decoder1_n61) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u362 ( .A(oc8051_decoder1_n427), .B(
        oc8051_decoder1_n61), .Y(oc8051_decoder1_n99) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u361 ( .A(oc8051_decoder1_n111), .B(
        oc8051_decoder1_n33), .Y(oc8051_decoder1_n426) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u360 ( .A(oc8051_decoder1_n71), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n105) );
  OAI222_X0P5M_A12TS oc8051_decoder1_u359 ( .A0(oc8051_decoder1_n30), .A1(
        oc8051_decoder1_n99), .B0(oc8051_decoder1_n112), .B1(
        oc8051_decoder1_n426), .C0(comp_sel[0]), .C1(oc8051_decoder1_n105), 
        .Y(comp_sel[1]) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u358 ( .A(oc8051_decoder1_n317), .B(
        oc8051_decoder1_n125), .C(oc8051_decoder1_state_0_), .Y(
        oc8051_decoder1_n277) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u357 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n132) );
  INV_X0P5B_A12TS oc8051_decoder1_u356 ( .A(oc8051_decoder1_n132), .Y(
        oc8051_decoder1_n281) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u355 ( .A(op1_cur[0]), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n23) );
  INV_X0P5B_A12TS oc8051_decoder1_u354 ( .A(oc8051_decoder1_n23), .Y(
        oc8051_decoder1_n244) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u353 ( .A(oc8051_decoder1_n54), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n155) );
  INV_X0P5B_A12TS oc8051_decoder1_u352 ( .A(oc8051_decoder1_n155), .Y(
        oc8051_decoder1_n40) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u351 ( .A(oc8051_decoder1_n21), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n48) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u350 ( .A(oc8051_decoder1_n132), .B(
        oc8051_decoder1_n48), .Y(oc8051_decoder1_n164) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u349 ( .A0(oc8051_decoder1_n105), .A1(
        oc8051_decoder1_n22), .A2(oc8051_decoder1_n164), .B0(
        oc8051_decoder1_n425), .B1(oc8051_decoder1_n137), .Y(
        oc8051_decoder1_n411) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u348 ( .A(oc8051_decoder1_n221), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n104) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u347 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n411), .B0(oc8051_decoder1_n25), .C0(
        oc8051_decoder1_n104), .Y(oc8051_decoder1_n410) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u346 ( .A0(oc8051_decoder1_n281), .A1(
        oc8051_decoder1_n161), .B0(oc8051_decoder1_n244), .B1(
        oc8051_decoder1_n40), .C0(oc8051_decoder1_n410), .Y(
        oc8051_decoder1_n386) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u345 ( .A0(oc8051_decoder1_n156), .A1(
        oc8051_decoder1_n50), .B0(oc8051_decoder1_n59), .Y(oc8051_decoder1_n24) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u344 ( .A(op1_cur[2]), .B(
        oc8051_decoder1_n69), .Y(oc8051_decoder1_n26) );
  INV_X0P5B_A12TS oc8051_decoder1_u343 ( .A(oc8051_decoder1_n26), .Y(
        oc8051_decoder1_n67) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u342 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n24), .A2(oc8051_decoder1_n67), .B0(
        oc8051_decoder1_state_1_), .Y(oc8051_decoder1_n387) );
  INV_X0P5B_A12TS oc8051_decoder1_u341 ( .A(oc8051_decoder1_n69), .Y(
        oc8051_decoder1_n9) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u340 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n265), .Y(oc8051_decoder1_n186) );
  INV_X0P5B_A12TS oc8051_decoder1_u339 ( .A(oc8051_decoder1_n186), .Y(
        oc8051_decoder1_n373) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u338 ( .A0(oc8051_decoder1_n59), .A1(
        oc8051_decoder1_n21), .B0(oc8051_decoder1_n373), .Y(
        oc8051_decoder1_n409) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u337 ( .A(oc8051_decoder1_n61), .B(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n98) );
  INV_X0P5B_A12TS oc8051_decoder1_u336 ( .A(oc8051_decoder1_n98), .Y(
        oc8051_decoder1_n353) );
  INV_X0P5B_A12TS oc8051_decoder1_u335 ( .A(oc8051_decoder1_n25), .Y(
        oc8051_decoder1_n44) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u334 ( .A0(oc8051_decoder1_n9), .A1(
        oc8051_decoder1_n54), .A2(oc8051_decoder1_n409), .B0(
        oc8051_decoder1_n353), .B1(oc8051_decoder1_n44), .Y(
        oc8051_decoder1_n404) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u333 ( .A0(oc8051_decoder1_n386), .A1(
        oc8051_decoder1_n36), .B0(oc8051_decoder1_n387), .C0(
        oc8051_decoder1_n404), .Y(oc8051_decoder1_n385) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u332 ( .A(oc8051_decoder1_n277), .B(
        oc8051_decoder1_n385), .Y(istb) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u331 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n18) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u330 ( .A0(oc8051_decoder1_n82), .A1(
        oc8051_decoder1_n21), .B0(oc8051_decoder1_n18), .Y(
        oc8051_decoder1_n251) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u329 ( .A(oc8051_decoder1_n251), .B(
        oc8051_decoder1_n161), .S0(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n380) );
  INV_X0P5B_A12TS oc8051_decoder1_u328 ( .A(oc8051_decoder1_n105), .Y(
        oc8051_decoder1_n47) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u327 ( .A(oc8051_decoder1_n185), .B(
        oc8051_decoder1_n47), .Y(oc8051_decoder1_n138) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u326 ( .A0(oc8051_decoder1_n138), .A1(
        oc8051_decoder1_n178), .B0(oc8051_decoder1_n40), .Y(
        oc8051_decoder1_n381) );
  INV_X0P5B_A12TS oc8051_decoder1_u325 ( .A(oc8051_decoder1_n193), .Y(
        oc8051_decoder1_n8) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u324 ( .A(oc8051_decoder1_n165), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n136) );
  INV_X0P5B_A12TS oc8051_decoder1_u323 ( .A(oc8051_decoder1_n136), .Y(
        oc8051_decoder1_n154) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u322 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n375), .B0(op1_cur[1]), .Y(oc8051_decoder1_n384) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u321 ( .A0(oc8051_decoder1_n8), .A1(
        oc8051_decoder1_n186), .B0(oc8051_decoder1_n154), .B1(
        oc8051_decoder1_n14), .C0(oc8051_decoder1_n384), .Y(
        oc8051_decoder1_n382) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u320 ( .A(oc8051_decoder1_n54), .B(
        op1_cur[1]), .Y(oc8051_decoder1_n245) );
  INV_X0P5B_A12TS oc8051_decoder1_u319 ( .A(oc8051_decoder1_n245), .Y(
        oc8051_decoder1_n142) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u318 ( .A(oc8051_decoder1_n9), .B(
        op1_cur[2]), .C(oc8051_decoder1_n142), .Y(oc8051_decoder1_n383) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u317 ( .A0(oc8051_decoder1_n380), .A1(
        oc8051_decoder1_n67), .A2(oc8051_decoder1_n381), .B0(
        oc8051_decoder1_n382), .B1(oc8051_decoder1_n383), .Y(
        oc8051_decoder1_n377) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u316 ( .A(oc8051_decoder1_n125), .B(
        oc8051_decoder1_n33), .Y(oc8051_decoder1_n144) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u315 ( .A(oc8051_decoder1_n139), .B(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n49) );
  INV_X0P5B_A12TS oc8051_decoder1_u314 ( .A(oc8051_decoder1_n49), .Y(
        oc8051_decoder1_n176) );
  INV_X0P5B_A12TS oc8051_decoder1_u313 ( .A(oc8051_decoder1_n144), .Y(
        oc8051_decoder1_n126) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u312 ( .A(oc8051_decoder1_n126), .B(
        oc8051_decoder1_n9), .Y(oc8051_decoder1_n166) );
  INV_X0P5B_A12TS oc8051_decoder1_u311 ( .A(oc8051_decoder1_n166), .Y(
        oc8051_decoder1_n330) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u310 ( .A(oc8051_decoder1_n176), .B(
        oc8051_decoder1_n330), .Y(oc8051_decoder1_n182) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u309 ( .A(oc8051_decoder1_n330), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n119) );
  OA22_X0P5M_A12TS oc8051_decoder1_u308 ( .A0(oc8051_decoder1_n251), .A1(
        oc8051_decoder1_n119), .B0(oc8051_decoder1_n379), .B1(
        oc8051_decoder1_n125), .Y(oc8051_decoder1_n378) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u307 ( .A0(oc8051_decoder1_n377), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n182), .C0(
        oc8051_decoder1_n378), .Y(oc8051_decoder1_n388) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u306 ( .A(oc8051_decoder1_n90), .B(
        op1_cur[1]), .Y(oc8051_decoder1_n355) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u305 ( .A(oc8051_decoder1_n244), .B(
        oc8051_decoder1_n281), .Y(oc8051_decoder1_n150) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u304 ( .A(oc8051_decoder1_n21), .B(
        oc8051_decoder1_n53), .Y(oc8051_decoder1_n217) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u303 ( .A(oc8051_decoder1_n257), .B(
        oc8051_decoder1_n136), .Y(oc8051_decoder1_n376) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u302 ( .A(oc8051_decoder1_n109), .B(
        oc8051_decoder1_n376), .S0(oc8051_decoder1_n21), .Y(
        oc8051_decoder1_n374) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u301 ( .A(oc8051_decoder1_n375), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n326) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u300 ( .A(oc8051_decoder1_n90), .B(
        oc8051_decoder1_n40), .Y(oc8051_decoder1_n157) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u299 ( .A(oc8051_decoder1_n326), .B(
        oc8051_decoder1_n157), .Y(oc8051_decoder1_n20) );
  AOI2XB1_X0P5M_A12TS oc8051_decoder1_u298 ( .A1N(oc8051_decoder1_n217), .A0(
        oc8051_decoder1_n374), .B0(oc8051_decoder1_n20), .Y(
        oc8051_decoder1_n351) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u297 ( .A0(oc8051_decoder1_n155), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n71), .B1(
        oc8051_decoder1_n48), .Y(oc8051_decoder1_n367) );
  INV_X0P5B_A12TS oc8051_decoder1_u296 ( .A(oc8051_decoder1_n367), .Y(
        oc8051_decoder1_n201) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u295 ( .A(oc8051_decoder1_n67), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n37) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u294 ( .A0(oc8051_decoder1_n201), .A1(
        oc8051_decoder1_n131), .B0(oc8051_decoder1_n37), .C0(
        oc8051_decoder1_n373), .Y(oc8051_decoder1_n369) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u293 ( .A(oc8051_decoder1_n40), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n370) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u292 ( .A0(oc8051_decoder1_n185), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n14), .B1(op1_cur[0]), .Y(
        oc8051_decoder1_n371) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u291 ( .A(oc8051_decoder1_n59), .B(
        oc8051_decoder1_n165), .S0(oc8051_decoder1_n137), .Y(
        oc8051_decoder1_n372) );
  INV_X0P5B_A12TS oc8051_decoder1_u290 ( .A(oc8051_decoder1_n157), .Y(
        oc8051_decoder1_n6) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u289 ( .A(oc8051_decoder1_n6), .B(
        op1_cur[1]), .Y(oc8051_decoder1_n350) );
  INV_X0P5B_A12TS oc8051_decoder1_u288 ( .A(oc8051_decoder1_n350), .Y(
        oc8051_decoder1_n146) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u287 ( .A0(oc8051_decoder1_n369), .A1(
        oc8051_decoder1_n370), .A2(oc8051_decoder1_n371), .B0(
        oc8051_decoder1_n372), .B1(oc8051_decoder1_n146), .Y(
        oc8051_decoder1_n368) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u286 ( .A0(oc8051_decoder1_n355), .A1(
        oc8051_decoder1_n150), .B0(oc8051_decoder1_n351), .C0(
        oc8051_decoder1_n368), .Y(oc8051_decoder1_n366) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u285 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n366), .B0(oc8051_decoder1_n330), .B1(
        oc8051_decoder1_n367), .Y(oc8051_decoder1_n365) );
  AO1B2_X0P5M_A12TS oc8051_decoder1_u284 ( .B0(psw_set[0]), .B1(wait_data), 
        .A0N(oc8051_decoder1_n365), .Y(oc8051_decoder1_n389) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u283 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n356) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u282 ( .A(oc8051_decoder1_n281), .B(
        oc8051_decoder1_n47), .Y(oc8051_decoder1_n292) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u281 ( .A(oc8051_decoder1_n292), .B(
        oc8051_decoder1_n166), .Y(oc8051_decoder1_n128) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u280 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n40), .A2(oc8051_decoder1_n330), .B0(
        oc8051_decoder1_n128), .Y(oc8051_decoder1_n357) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u279 ( .A(oc8051_decoder1_n281), .B(
        oc8051_decoder1_n42), .Y(oc8051_decoder1_n202) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u278 ( .A(oc8051_decoder1_n217), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n13) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u277 ( .A0(oc8051_decoder1_n155), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n202), .C0(
        oc8051_decoder1_n13), .Y(oc8051_decoder1_n362) );
  INV_X0P5B_A12TS oc8051_decoder1_u276 ( .A(oc8051_decoder1_n356), .Y(
        oc8051_decoder1_n70) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u275 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n40), .B0(oc8051_decoder1_n176), .C0(op1_cur[1]), .Y(
        oc8051_decoder1_n364) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u274 ( .A0(oc8051_decoder1_n25), .A1(
        oc8051_decoder1_n292), .B0(oc8051_decoder1_n326), .B1(
        oc8051_decoder1_n48), .C0(oc8051_decoder1_n364), .Y(
        oc8051_decoder1_n363) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u273 ( .A0(oc8051_decoder1_n178), .A1(
        oc8051_decoder1_n362), .B0(oc8051_decoder1_n70), .B1(
        oc8051_decoder1_n185), .C0(oc8051_decoder1_n363), .Y(
        oc8051_decoder1_n360) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u272 ( .A(oc8051_decoder1_n50), .B(
        oc8051_decoder1_n157), .C(oc8051_decoder1_n265), .Y(
        oc8051_decoder1_n279) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u271 ( .A0(oc8051_decoder1_n47), .A1(
        op1_cur[0]), .A2(oc8051_decoder1_n146), .B0(oc8051_decoder1_n279), .Y(
        oc8051_decoder1_n361) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u270 ( .A0(oc8051_decoder1_n360), .A1(
        oc8051_decoder1_n26), .B0(oc8051_decoder1_n270), .B1(
        oc8051_decoder1_n356), .C0(oc8051_decoder1_n361), .Y(
        oc8051_decoder1_n359) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u269 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n359), .B0(src_sel2[0]), .B1(wait_data), .Y(
        oc8051_decoder1_n358) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u268 ( .A0(oc8051_decoder1_n119), .A1(
        oc8051_decoder1_n356), .B0(oc8051_decoder1_n357), .C0(
        oc8051_decoder1_n358), .Y(oc8051_decoder1_n390) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u267 ( .A(op1_cur[2]), .B(
        oc8051_decoder1_n69), .C(oc8051_decoder1_n54), .Y(oc8051_decoder1_n116) );
  INV_X0P5B_A12TS oc8051_decoder1_u266 ( .A(oc8051_decoder1_n116), .Y(
        oc8051_decoder1_n293) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u265 ( .A(oc8051_decoder1_n126), .B(
        oc8051_decoder1_n293), .Y(oc8051_decoder1_n212) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u264 ( .A0(oc8051_decoder1_n155), .A1(
        oc8051_decoder1_n166), .B0(oc8051_decoder1_n50), .B1(
        oc8051_decoder1_n212), .Y(oc8051_decoder1_n347) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u263 ( .A0(oc8051_decoder1_n137), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n55), .Y(
        oc8051_decoder1_n262) );
  INV_X0P5B_A12TS oc8051_decoder1_u262 ( .A(oc8051_decoder1_n262), .Y(
        oc8051_decoder1_n349) );
  INV_X0P5B_A12TS oc8051_decoder1_u261 ( .A(oc8051_decoder1_n355), .Y(
        oc8051_decoder1_n16) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u260 ( .A(oc8051_decoder1_n265), .B(
        oc8051_decoder1_n155), .C(oc8051_decoder1_n26), .Y(
        oc8051_decoder1_n287) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u259 ( .A(oc8051_decoder1_n67), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n27) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u258 ( .A(oc8051_decoder1_n27), .B(
        oc8051_decoder1_n14), .C(oc8051_decoder1_n82), .Y(oc8051_decoder1_n354) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u257 ( .A0(oc8051_decoder1_n353), .A1(
        oc8051_decoder1_n16), .B0(oc8051_decoder1_n287), .C0(
        oc8051_decoder1_n354), .Y(oc8051_decoder1_n352) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u256 ( .A0(oc8051_decoder1_n349), .A1(
        oc8051_decoder1_n350), .B0(oc8051_decoder1_n351), .C0(
        oc8051_decoder1_n352), .Y(oc8051_decoder1_n348) );
  AOI222_X0P5M_A12TS oc8051_decoder1_u255 ( .A0(cy_sel[0]), .A1(wait_data), 
        .B0(oc8051_decoder1_n156), .B1(oc8051_decoder1_n347), .C0(
        oc8051_decoder1_n126), .C1(oc8051_decoder1_n348), .Y(
        oc8051_decoder1_n342) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u254 ( .A(oc8051_decoder1_n47), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n211) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u253 ( .A0(op1_cur[1]), .A1(
        oc8051_decoder1_n225), .B0(oc8051_decoder1_n211), .C0(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n344) );
  INV_X0P5B_A12TS oc8051_decoder1_u252 ( .A(oc8051_decoder1_n212), .Y(
        oc8051_decoder1_n273) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u251 ( .A(oc8051_decoder1_n166), .B(
        oc8051_decoder1_n82), .C(oc8051_decoder1_n48), .Y(oc8051_decoder1_n345) );
  INV_X0P5B_A12TS oc8051_decoder1_u250 ( .A(oc8051_decoder1_n182), .Y(
        oc8051_decoder1_n346) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u249 ( .A0(oc8051_decoder1_n344), .A1(
        oc8051_decoder1_n273), .B0(oc8051_decoder1_n345), .C0(
        oc8051_decoder1_n346), .Y(oc8051_decoder1_n343) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u248 ( .A(oc8051_decoder1_n342), .B(
        oc8051_decoder1_n343), .Y(oc8051_decoder1_n391) );
  INV_X0P5B_A12TS oc8051_decoder1_u247 ( .A(oc8051_decoder1_n27), .Y(
        oc8051_decoder1_n189) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u246 ( .A(oc8051_decoder1_n44), .B(
        oc8051_decoder1_n61), .C(oc8051_decoder1_n293), .Y(
        oc8051_decoder1_n114) );
  INV_X0P5B_A12TS oc8051_decoder1_u245 ( .A(oc8051_decoder1_n115), .Y(
        oc8051_decoder1_n341) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u244 ( .A(oc8051_decoder1_n9), .B(
        oc8051_decoder1_n54), .C(oc8051_decoder1_n341), .Y(
        oc8051_decoder1_n113) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u243 ( .A(oc8051_decoder1_n341), .B(
        oc8051_decoder1_n54), .C(oc8051_decoder1_n25), .D(op1_cur[2]), .Y(
        oc8051_decoder1_n340) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u242 ( .A(oc8051_decoder1_n114), .B(
        oc8051_decoder1_n113), .C(oc8051_decoder1_n340), .Y(
        oc8051_decoder1_n339) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u241 ( .A(oc8051_decoder1_n224), .B(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n325) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u240 ( .A(op1_cur[0]), .B(op1_cur[1]), .C(
        oc8051_decoder1_n224), .Y(oc8051_decoder1_n102) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u239 ( .A0(oc8051_decoder1_n325), .A1(
        oc8051_decoder1_n226), .B0(oc8051_decoder1_n102), .B1(
        oc8051_decoder1_n236), .Y(oc8051_decoder1_n291) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u238 ( .A0(oc8051_decoder1_n275), .A1(
        oc8051_decoder1_n189), .B0(oc8051_decoder1_n339), .C0(
        oc8051_decoder1_n291), .Y(oc8051_decoder1_n335) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u237 ( .A(src_sel2[1]), .B(wait_data), .Y(
        oc8051_decoder1_n336) );
  INV_X0P5B_A12TS oc8051_decoder1_u236 ( .A(oc8051_decoder1_n226), .Y(
        oc8051_decoder1_n207) );
  INV_X0P5B_A12TS oc8051_decoder1_u235 ( .A(oc8051_decoder1_n48), .Y(
        oc8051_decoder1_n135) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u234 ( .A(oc8051_decoder1_n135), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n12) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u233 ( .A0(oc8051_decoder1_n98), .A1(
        oc8051_decoder1_n12), .B0(oc8051_decoder1_n166), .Y(
        oc8051_decoder1_n338) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u232 ( .A0(oc8051_decoder1_n207), .A1(
        oc8051_decoder1_n178), .A2(oc8051_decoder1_n273), .B0(
        oc8051_decoder1_n338), .Y(oc8051_decoder1_n337) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u231 ( .A0(oc8051_decoder1_n335), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n336), .C0(
        oc8051_decoder1_n337), .Y(oc8051_decoder1_n392) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u230 ( .A0(oc8051_decoder1_n115), .A1(
        oc8051_decoder1_n193), .A2(oc8051_decoder1_n334), .B0(
        oc8051_decoder1_n114), .Y(oc8051_decoder1_n332) );
  INV_X0P5B_A12TS oc8051_decoder1_u229 ( .A(oc8051_decoder1_n102), .Y(
        oc8051_decoder1_n269) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u228 ( .A0(oc8051_decoder1_n8), .A1(
        oc8051_decoder1_n224), .B0(oc8051_decoder1_n269), .Y(
        oc8051_decoder1_n324) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u227 ( .A0(oc8051_decoder1_n82), .A1(
        oc8051_decoder1_n225), .B0(oc8051_decoder1_n236), .C0(
        oc8051_decoder1_n324), .Y(oc8051_decoder1_n333) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u226 ( .A0(oc8051_decoder1_n189), .A1(
        oc8051_decoder1_n207), .B0(oc8051_decoder1_n332), .C0(
        oc8051_decoder1_n333), .Y(oc8051_decoder1_n327) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u225 ( .A(oc8051_decoder1_n225), .B(
        oc8051_decoder1_n212), .Y(oc8051_decoder1_n331) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u224 ( .A0(op1_cur[1]), .A1(
        oc8051_decoder1_n44), .B0(oc8051_decoder1_n82), .C0(
        oc8051_decoder1_n331), .Y(oc8051_decoder1_n328) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u223 ( .A0(oc8051_decoder1_n54), .A1(
        oc8051_decoder1_n226), .B0(oc8051_decoder1_n49), .Y(
        oc8051_decoder1_n197) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u222 ( .A0(oc8051_decoder1_n330), .A1(
        oc8051_decoder1_n197), .B0(cy_sel[1]), .B1(wait_data), .Y(
        oc8051_decoder1_n329) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u221 ( .A0(oc8051_decoder1_n327), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n328), .C0(
        oc8051_decoder1_n329), .Y(oc8051_decoder1_n393) );
  INV_X0P5B_A12TS oc8051_decoder1_u220 ( .A(oc8051_decoder1_n326), .Y(
        oc8051_decoder1_n320) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u219 ( .A(oc8051_decoder1_n47), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n181) );
  INV_X0P5B_A12TS oc8051_decoder1_u218 ( .A(oc8051_decoder1_n181), .Y(
        oc8051_decoder1_n219) );
  INV_X0P5B_A12TS oc8051_decoder1_u217 ( .A(oc8051_decoder1_n325), .Y(
        oc8051_decoder1_n60) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u216 ( .A(oc8051_decoder1_n219), .B(
        oc8051_decoder1_n60), .Y(oc8051_decoder1_n78) );
  OA22_X0P5M_A12TS oc8051_decoder1_u215 ( .A0(oc8051_decoder1_n225), .A1(
        oc8051_decoder1_n324), .B0(oc8051_decoder1_n105), .B1(
        oc8051_decoder1_n102), .Y(oc8051_decoder1_n323) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u214 ( .A0(oc8051_decoder1_n219), .A1(
        oc8051_decoder1_n322), .B0(oc8051_decoder1_n78), .C0(
        oc8051_decoder1_n323), .Y(oc8051_decoder1_n321) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u213 ( .A0(oc8051_decoder1_n273), .A1(
        oc8051_decoder1_n320), .A2(oc8051_decoder1_n70), .B0(
        oc8051_decoder1_n126), .B1(oc8051_decoder1_n321), .Y(
        oc8051_decoder1_n319) );
  AO1B2_X0P5M_A12TS oc8051_decoder1_u212 ( .B0(src_sel3), .B1(wait_data), 
        .A0N(oc8051_decoder1_n319), .Y(oc8051_decoder1_n394) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u211 ( .A(wait_data), .B(mem_wait), .Y(
        oc8051_decoder1_n296) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u210 ( .A0(oc8051_decoder1_n296), .A1(
        oc8051_decoder1_n316), .B0(oc8051_decoder1_n317), .C0(
        oc8051_decoder1_n318), .Y(oc8051_decoder1_n395) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u209 ( .A(oc8051_decoder1_n314), .B(
        oc8051_decoder1_n315), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n396) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u208 ( .A(oc8051_decoder1_n299), .B(
        oc8051_decoder1_n313), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n397) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u207 ( .A(oc8051_decoder1_n311), .B(
        oc8051_decoder1_n312), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n398) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u206 ( .A(oc8051_decoder1_n300), .B(
        oc8051_decoder1_n310), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n399) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u205 ( .A(oc8051_decoder1_n308), .B(
        oc8051_decoder1_n309), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n400) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u204 ( .A(oc8051_decoder1_n306), .B(
        oc8051_decoder1_n307), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n401) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u203 ( .A(oc8051_decoder1_n304), .B(
        oc8051_decoder1_n305), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n402) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u202 ( .A(oc8051_decoder1_n301), .B(
        oc8051_decoder1_n302), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n403) );
  XOR2_X0P5M_A12TS oc8051_decoder1_u201 ( .A(op1_n[7]), .B(op1_n[5]), .Y(
        oc8051_decoder1_n298) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u200 ( .A0(oc8051_decoder1_n298), .A1(
        oc8051_decoder1_n299), .A2(op1_n[1]), .B0(op1_n[2]), .B1(
        oc8051_decoder1_n300), .Y(oc8051_decoder1_n297) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u199 ( .A(oc8051_decoder1_state_0_), .B(
        oc8051_decoder1_n297), .Y(oc8051_decoder1_n295) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u198 ( .A(oc8051_decoder1_state_0_), .B(
        oc8051_decoder1_n295), .S0(oc8051_decoder1_n296), .Y(
        oc8051_decoder1_n294) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u197 ( .A0(mem_wait), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n294), .Y(
        oc8051_decoder1_n405) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u196 ( .A(oc8051_decoder1_n293), .B(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n180) );
  INV_X0P5B_A12TS oc8051_decoder1_u195 ( .A(oc8051_decoder1_n52), .Y(
        oc8051_decoder1_n68) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u194 ( .A(oc8051_decoder1_n68), .B(
        oc8051_decoder1_n293), .C(oc8051_decoder1_n82), .D(oc8051_decoder1_n22), .Y(oc8051_decoder1_n122) );
  OA21_X0P5M_A12TS oc8051_decoder1_u193 ( .A0(oc8051_decoder1_n180), .A1(
        oc8051_decoder1_n181), .B0(oc8051_decoder1_n122), .Y(
        oc8051_decoder1_n255) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u192 ( .A(oc8051_decoder1_n277), .B(
        oc8051_decoder1_n255), .Y(oc8051_decoder1_n228) );
  INV_X0P5B_A12TS oc8051_decoder1_u191 ( .A(oc8051_decoder1_n228), .Y(
        oc8051_decoder1_n229) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u190 ( .A(oc8051_decoder1_n219), .B(
        oc8051_decoder1_n44), .C(oc8051_decoder1_n273), .Y(
        oc8051_decoder1_n213) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u189 ( .A0(oc8051_decoder1_n408), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n229), .C0(
        oc8051_decoder1_n213), .Y(oc8051_decoder1_n412) );
  INV_X0P5B_A12TS oc8051_decoder1_u188 ( .A(oc8051_decoder1_n292), .Y(
        oc8051_decoder1_n290) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u187 ( .A0(oc8051_decoder1_n290), .A1(
        oc8051_decoder1_n36), .B0(oc8051_decoder1_n291), .C0(
        oc8051_decoder1_n126), .Y(oc8051_decoder1_n288) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u186 ( .A0(oc8051_decoder1_n61), .A1(
        op1_cur[1]), .A2(oc8051_decoder1_n273), .B0(oc8051_decoder1_n228), .Y(
        oc8051_decoder1_n289) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u185 ( .A0(oc8051_decoder1_n406), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n288), .C0(
        oc8051_decoder1_n289), .Y(oc8051_decoder1_n413) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u184 ( .A0(oc8051_decoder1_n42), .A1(
        oc8051_decoder1_n16), .B0(oc8051_decoder1_n75), .Y(
        oc8051_decoder1_n284) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u183 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n23), .B0(oc8051_decoder1_n104), .Y(
        oc8051_decoder1_n190) );
  INV_X0P5B_A12TS oc8051_decoder1_u182 ( .A(oc8051_decoder1_n190), .Y(
        oc8051_decoder1_n286) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u181 ( .A0(oc8051_decoder1_n286), .A1(
        oc8051_decoder1_n189), .B0(oc8051_decoder1_n287), .C0(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n285) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u180 ( .A0(oc8051_decoder1_n284), .A1(
        oc8051_decoder1_n14), .A2(oc8051_decoder1_n137), .B0(
        oc8051_decoder1_n285), .Y(oc8051_decoder1_n278) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u179 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n131), .B0(oc8051_decoder1_n69), .Y(
        oc8051_decoder1_n41) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u178 ( .A(oc8051_decoder1_n283), .B(
        oc8051_decoder1_n12), .C(oc8051_decoder1_n41), .Y(oc8051_decoder1_n282) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u177 ( .A0(oc8051_decoder1_n281), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n40), .B1(
        oc8051_decoder1_n265), .C0(oc8051_decoder1_n282), .Y(
        oc8051_decoder1_n280) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u176 ( .A0(oc8051_decoder1_n278), .A1(
        oc8051_decoder1_n279), .A2(oc8051_decoder1_n280), .B0(
        oc8051_decoder1_n126), .Y(oc8051_decoder1_n271) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u175 ( .A0(oc8051_decoder1_n50), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n47), .Y(
        oc8051_decoder1_n274) );
  AND4_X0P5M_A12TS oc8051_decoder1_u174 ( .A(oc8051_decoder1_n42), .B(
        oc8051_decoder1_n224), .C(oc8051_decoder1_n14), .D(oc8051_decoder1_n25), .Y(oc8051_decoder1_n276) );
  INV_X0P5B_A12TS oc8051_decoder1_u173 ( .A(oc8051_decoder1_n277), .Y(
        oc8051_decoder1_n183) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u172 ( .A0(oc8051_decoder1_n275), .A1(
        oc8051_decoder1_n269), .B0(oc8051_decoder1_n276), .C0(
        oc8051_decoder1_n183), .Y(oc8051_decoder1_n267) );
  INV_X0P5B_A12TS oc8051_decoder1_u171 ( .A(oc8051_decoder1_n267), .Y(
        oc8051_decoder1_n241) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u170 ( .A0(oc8051_decoder1_n273), .A1(
        oc8051_decoder1_n14), .A2(oc8051_decoder1_n274), .B0(
        oc8051_decoder1_n241), .Y(oc8051_decoder1_n272) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u169 ( .A0(oc8051_decoder1_n407), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n271), .C0(
        oc8051_decoder1_n272), .Y(oc8051_decoder1_n414) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u168 ( .A(oc8051_decoder1_n165), .B(
        oc8051_decoder1_n90), .C(oc8051_decoder1_n44), .Y(oc8051_decoder1_n200) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u167 ( .A0(oc8051_decoder1_n270), .A1(
        oc8051_decoder1_n226), .B0(oc8051_decoder1_n200), .Y(
        oc8051_decoder1_n218) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u166 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n111), .B0(oc8051_decoder1_n218), .Y(
        oc8051_decoder1_n230) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u165 ( .A0(oc8051_decoder1_n219), .A1(
        oc8051_decoder1_n269), .A2(oc8051_decoder1_n126), .B0(src_sel1[2]), 
        .B1(wait_data), .Y(oc8051_decoder1_n268) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u164 ( .A(oc8051_decoder1_n267), .B(
        oc8051_decoder1_n230), .C(oc8051_decoder1_n268), .Y(
        oc8051_decoder1_n415) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u163 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n185), .B0(oc8051_decoder1_n161), .Y(
        oc8051_decoder1_n266) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u162 ( .A(oc8051_decoder1_n265), .B(
        oc8051_decoder1_n266), .S0(oc8051_decoder1_n164), .Y(
        oc8051_decoder1_n252) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u161 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n185), .B1(
        oc8051_decoder1_n50), .Y(oc8051_decoder1_n259) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u160 ( .A(oc8051_decoder1_n154), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n264) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u159 ( .A(oc8051_decoder1_n217), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n38) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u158 ( .A0(oc8051_decoder1_n137), .A1(
        oc8051_decoder1_n165), .B0(oc8051_decoder1_n38), .Y(
        oc8051_decoder1_n250) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u157 ( .A(oc8051_decoder1_n264), .B(
        oc8051_decoder1_n250), .S0(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n263) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u156 ( .A0(oc8051_decoder1_n135), .A1(
        oc8051_decoder1_n262), .B0(oc8051_decoder1_n263), .Y(
        oc8051_decoder1_n261) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u155 ( .A(oc8051_decoder1_n252), .B(
        oc8051_decoder1_n261), .S0(oc8051_decoder1_n22), .Y(
        oc8051_decoder1_n260) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u154 ( .A0(oc8051_decoder1_n90), .A1(
        oc8051_decoder1_n259), .A2(oc8051_decoder1_n207), .B0(
        oc8051_decoder1_n260), .B1(oc8051_decoder1_n67), .Y(
        oc8051_decoder1_n258) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u153 ( .A0(oc8051_decoder1_n11), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n257), .C0(
        oc8051_decoder1_n258), .Y(oc8051_decoder1_n256) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u152 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n256), .B0(oc8051_decoder1_n241), .Y(
        oc8051_decoder1_n253) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u151 ( .A(oc8051_decoder1_state_1_), .B(
        oc8051_decoder1_n125), .C(oc8051_decoder1_state_0_), .Y(
        oc8051_decoder1_n184) );
  NAND3B_X0P5M_A12TS oc8051_decoder1_u150 ( .AN(oc8051_decoder1_n180), .B(
        oc8051_decoder1_n82), .C(oc8051_decoder1_n21), .Y(oc8051_decoder1_n101) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u149 ( .A0(oc8051_decoder1_n184), .A1(
        oc8051_decoder1_n101), .B0(oc8051_decoder1_n255), .B1(
        oc8051_decoder1_n30), .C0(oc8051_decoder1_n229), .Y(
        oc8051_decoder1_n203) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u148 ( .A0(src_sel1[1]), .A1(wait_data), 
        .B0(oc8051_decoder1_n203), .Y(oc8051_decoder1_n254) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u147 ( .A0(oc8051_decoder1_n166), .A1(
        oc8051_decoder1_n252), .B0(oc8051_decoder1_n253), .C0(
        oc8051_decoder1_n254), .Y(oc8051_decoder1_n416) );
  OAI222_X0P5M_A12TS oc8051_decoder1_u146 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n132), .B0(oc8051_decoder1_n54), .B1(
        oc8051_decoder1_n251), .C0(oc8051_decoder1_n156), .C1(
        oc8051_decoder1_n155), .Y(oc8051_decoder1_n237) );
  INV_X0P5B_A12TS oc8051_decoder1_u145 ( .A(oc8051_decoder1_n237), .Y(
        oc8051_decoder1_n247) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u144 ( .A(oc8051_decoder1_n25), .B(
        oc8051_decoder1_n186), .Y(oc8051_decoder1_n249) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u143 ( .A(oc8051_decoder1_n249), .B(
        oc8051_decoder1_n250), .S0(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n248) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u142 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n247), .B0(oc8051_decoder1_n48), .B1(
        oc8051_decoder1_n23), .C0(oc8051_decoder1_n248), .Y(
        oc8051_decoder1_n242) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u141 ( .A(oc8051_decoder1_n154), .B(
        oc8051_decoder1_n38), .S0(op1_cur[1]), .Y(oc8051_decoder1_n246) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u140 ( .A0(op1_cur[0]), .A1(
        oc8051_decoder1_n156), .B0(oc8051_decoder1_n244), .B1(
        oc8051_decoder1_n245), .C0(oc8051_decoder1_n246), .Y(
        oc8051_decoder1_n243) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u139 ( .A(oc8051_decoder1_n242), .B(
        oc8051_decoder1_n243), .S0(oc8051_decoder1_n131), .Y(
        oc8051_decoder1_n240) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u138 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n69), .A2(oc8051_decoder1_n240), .B0(
        oc8051_decoder1_n241), .Y(oc8051_decoder1_n238) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u137 ( .A0(src_sel1[0]), .A1(wait_data), 
        .B0(oc8051_decoder1_n203), .Y(oc8051_decoder1_n239) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u136 ( .A0(oc8051_decoder1_n166), .A1(
        oc8051_decoder1_n237), .B0(oc8051_decoder1_n238), .C0(
        oc8051_decoder1_n239), .Y(oc8051_decoder1_n417) );
  INV_X0P5B_A12TS oc8051_decoder1_u135 ( .A(oc8051_decoder1_n211), .Y(
        oc8051_decoder1_n222) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u134 ( .A(oc8051_decoder1_n126), .B(
        oc8051_decoder1_n60), .C(oc8051_decoder1_n222), .Y(
        oc8051_decoder1_n231) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u133 ( .A(oc8051_decoder1_n226), .B(
        oc8051_decoder1_n181), .Y(oc8051_decoder1_n108) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u132 ( .A0(oc8051_decoder1_n189), .A1(
        oc8051_decoder1_n108), .B0(oc8051_decoder1_n221), .B1(
        oc8051_decoder1_n67), .Y(oc8051_decoder1_n234) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u131 ( .A0(oc8051_decoder1_n11), .A1(
        oc8051_decoder1_n211), .A2(oc8051_decoder1_n236), .B0(
        oc8051_decoder1_n212), .Y(oc8051_decoder1_n235) );
  OAI21B_X0P5M_A12TS oc8051_decoder1_u130 ( .A0(oc8051_decoder1_n234), .A1(
        oc8051_decoder1_n144), .B0N(oc8051_decoder1_n235), .Y(
        oc8051_decoder1_n233) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u129 ( .A0(oc8051_decoder1_n233), .A1(
        op1_cur[1]), .B0(wait_data), .B1(oc8051_decoder1_ram_wr_sel_1_), .Y(
        oc8051_decoder1_n232) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u128 ( .A(oc8051_decoder1_n229), .B(
        oc8051_decoder1_n230), .C(oc8051_decoder1_n231), .D(
        oc8051_decoder1_n232), .Y(oc8051_decoder1_n418) );
  INV_X0P5B_A12TS oc8051_decoder1_u127 ( .A(oc8051_decoder1_ram_wr_sel_0_), 
        .Y(oc8051_decoder1_n28) );
  AND4_X0P5M_A12TS oc8051_decoder1_u126 ( .A(oc8051_decoder1_n207), .B(
        oc8051_decoder1_n90), .C(oc8051_decoder1_n185), .D(oc8051_decoder1_n22), .Y(oc8051_decoder1_n227) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u125 ( .A0(oc8051_decoder1_n218), .A1(
        oc8051_decoder1_n227), .B0(oc8051_decoder1_n111), .C0(
        oc8051_decoder1_n228), .Y(oc8051_decoder1_n188) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u124 ( .A0(oc8051_decoder1_n115), .A1(
        oc8051_decoder1_n225), .A2(oc8051_decoder1_n226), .B0(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n223) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u123 ( .A0(oc8051_decoder1_n222), .A1(
        oc8051_decoder1_n223), .B0(oc8051_decoder1_n137), .C0(
        oc8051_decoder1_n224), .Y(oc8051_decoder1_n214) );
  AO22_X0P5M_A12TS oc8051_decoder1_u122 ( .A0(oc8051_decoder1_n69), .A1(
        oc8051_decoder1_n221), .B0(oc8051_decoder1_n108), .B1(
        oc8051_decoder1_n189), .Y(oc8051_decoder1_n220) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u121 ( .A0(oc8051_decoder1_n54), .A1(
        oc8051_decoder1_n41), .A2(oc8051_decoder1_n219), .B0(
        oc8051_decoder1_n44), .B1(oc8051_decoder1_n220), .Y(
        oc8051_decoder1_n215) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u120 ( .A0(oc8051_decoder1_n60), .A1(
        oc8051_decoder1_n61), .B0(oc8051_decoder1_n75), .B1(
        oc8051_decoder1_n217), .C0(oc8051_decoder1_n218), .Y(
        oc8051_decoder1_n216) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u119 ( .A(oc8051_decoder1_n214), .B(
        oc8051_decoder1_n114), .C(oc8051_decoder1_n215), .D(
        oc8051_decoder1_n216), .Y(oc8051_decoder1_n209) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u118 ( .A0(oc8051_decoder1_n211), .A1(
        oc8051_decoder1_n25), .A2(oc8051_decoder1_n212), .B0(
        oc8051_decoder1_n213), .Y(oc8051_decoder1_n210) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u117 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n209), .B0(oc8051_decoder1_n210), .Y(
        oc8051_decoder1_n208) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u116 ( .A0(oc8051_decoder1_n28), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n188), .C0(
        oc8051_decoder1_n208), .Y(oc8051_decoder1_n419) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u115 ( .A0(oc8051_decoder1_n135), .A1(
        oc8051_decoder1_n161), .B0(oc8051_decoder1_n207), .B1(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n206) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u114 ( .A0(oc8051_decoder1_n90), .A1(
        oc8051_decoder1_n206), .B0(oc8051_decoder1_n101), .Y(
        oc8051_decoder1_n205) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u113 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n205), .B0(psw_set[1]), .B1(wait_data), .Y(
        oc8051_decoder1_n204) );
  NAND2B_X0P5M_A12TS oc8051_decoder1_u112 ( .AN(oc8051_decoder1_n203), .B(
        oc8051_decoder1_n204), .Y(oc8051_decoder1_n420) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u111 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n47), .C0(
        oc8051_decoder1_n44), .Y(oc8051_decoder1_n198) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u110 ( .A(oc8051_decoder1_n201), .B(
        oc8051_decoder1_n202), .C(oc8051_decoder1_n41), .D(oc8051_decoder1_n13), .Y(oc8051_decoder1_n199) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u109 ( .A0(oc8051_decoder1_n116), .A1(
        oc8051_decoder1_n198), .B0(oc8051_decoder1_n199), .C0(
        oc8051_decoder1_n200), .Y(oc8051_decoder1_n191) );
  INV_X0P5B_A12TS oc8051_decoder1_u108 ( .A(oc8051_decoder1_n197), .Y(
        oc8051_decoder1_n196) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u107 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n13), .B0(oc8051_decoder1_n196), .B1(
        oc8051_decoder1_n193), .Y(oc8051_decoder1_n195) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u106 ( .A0(oc8051_decoder1_n176), .A1(
        oc8051_decoder1_n178), .B0(oc8051_decoder1_n195), .C0(
        oc8051_decoder1_n90), .Y(oc8051_decoder1_n194) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u105 ( .A0(oc8051_decoder1_n193), .A1(
        oc8051_decoder1_n157), .A2(oc8051_decoder1_n82), .B0(
        oc8051_decoder1_n194), .Y(oc8051_decoder1_n192) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u104 ( .A0(oc8051_decoder1_n189), .A1(
        oc8051_decoder1_n190), .B0(oc8051_decoder1_n191), .C0(
        oc8051_decoder1_n192), .Y(oc8051_decoder1_n187) );
  INV_X0P5B_A12TS oc8051_decoder1_u103 ( .A(oc8051_decoder1_wr), .Y(
        oc8051_decoder1_n1) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u102 ( .A0(oc8051_decoder1_n187), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n1), .B1(
        oc8051_decoder1_n125), .C0(oc8051_decoder1_n188), .Y(
        oc8051_decoder1_n421) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u101 ( .A(oc8051_decoder1_n185), .B(
        oc8051_decoder1_n18), .C(oc8051_decoder1_n186), .Y(
        oc8051_decoder1_n151) );
  INV_X0P5B_A12TS oc8051_decoder1_u100 ( .A(oc8051_decoder1_n184), .Y(
        oc8051_decoder1_n110) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u99 ( .A(oc8051_decoder1_n110), .B(
        oc8051_decoder1_n183), .C(oc8051_decoder1_n111), .Y(
        oc8051_decoder1_n123) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u98 ( .A0(oc8051_decoder1_n180), .A1(
        oc8051_decoder1_n123), .A2(oc8051_decoder1_n181), .B0(
        oc8051_decoder1_n182), .Y(oc8051_decoder1_n179) );
  INV_X0P5B_A12TS oc8051_decoder1_u97 ( .A(oc8051_decoder1_n179), .Y(
        oc8051_decoder1_n167) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u96 ( .A0(op1_cur[0]), .A1(
        oc8051_decoder1_n105), .B0(oc8051_decoder1_n59), .Y(
        oc8051_decoder1_n147) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u95 ( .A0(oc8051_decoder1_n132), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n105), .B1(
        oc8051_decoder1_n155), .Y(oc8051_decoder1_n177) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u94 ( .A0(op1_cur[1]), .A1(
        oc8051_decoder1_n176), .B0(oc8051_decoder1_n177), .B1(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n175) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u93 ( .A0(oc8051_decoder1_n175), .A1(
        oc8051_decoder1_n151), .A2(oc8051_decoder1_n150), .B0(
        oc8051_decoder1_n26), .Y(oc8051_decoder1_n171) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u92 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n23), .B0(oc8051_decoder1_n11), .Y(
        oc8051_decoder1_n174) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u91 ( .A0(oc8051_decoder1_n6), .A1(
        oc8051_decoder1_n137), .A2(oc8051_decoder1_n53), .B0(
        oc8051_decoder1_n75), .B1(oc8051_decoder1_n174), .Y(
        oc8051_decoder1_n173) );
  INV_X0P5B_A12TS oc8051_decoder1_u90 ( .A(oc8051_decoder1_n173), .Y(
        oc8051_decoder1_n172) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u89 ( .A0(oc8051_decoder1_n147), .A1(
        oc8051_decoder1_n146), .B0(oc8051_decoder1_n171), .C0(
        oc8051_decoder1_n172), .Y(oc8051_decoder1_n170) );
  INV_X0P5B_A12TS oc8051_decoder1_u88 ( .A(oc8051_decoder1_n170), .Y(
        oc8051_decoder1_n169) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u87 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n169), .B0(oc8051_decoder1_alu_op_2_), .B1(wait_data), 
        .Y(oc8051_decoder1_n168) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u86 ( .A0(oc8051_decoder1_n166), .A1(
        oc8051_decoder1_n151), .B0(oc8051_decoder1_n167), .C0(
        oc8051_decoder1_n168), .Y(oc8051_decoder1_n422) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u85 ( .A(oc8051_decoder1_n137), .B(
        oc8051_decoder1_n82), .S0(oc8051_decoder1_n14), .Y(
        oc8051_decoder1_n159) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u84 ( .A0(oc8051_decoder1_n156), .A1(
        oc8051_decoder1_n54), .B0(oc8051_decoder1_n165), .Y(
        oc8051_decoder1_n162) );
  INV_X0P5B_A12TS oc8051_decoder1_u83 ( .A(oc8051_decoder1_n164), .Y(
        oc8051_decoder1_n163) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u82 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n162), .S0(oc8051_decoder1_n163), .Y(
        oc8051_decoder1_n160) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u81 ( .A0(oc8051_decoder1_n141), .A1(
        oc8051_decoder1_n75), .A2(oc8051_decoder1_n159), .B0(
        oc8051_decoder1_n160), .B1(oc8051_decoder1_n41), .Y(
        oc8051_decoder1_n158) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u80 ( .A0(oc8051_decoder1_n58), .A1(
        oc8051_decoder1_n157), .A2(oc8051_decoder1_n50), .B0(
        oc8051_decoder1_n158), .Y(oc8051_decoder1_n148) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u79 ( .A0(oc8051_decoder1_n47), .A1(
        oc8051_decoder1_n155), .B0(oc8051_decoder1_n156), .B1(
        oc8051_decoder1_n132), .Y(oc8051_decoder1_n153) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u78 ( .A0(oc8051_decoder1_n153), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n154), .B1(
        oc8051_decoder1_n40), .Y(oc8051_decoder1_n152) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u77 ( .A0(oc8051_decoder1_n150), .A1(
        oc8051_decoder1_n151), .A2(oc8051_decoder1_n152), .B0(
        oc8051_decoder1_n37), .Y(oc8051_decoder1_n149) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u76 ( .A0(oc8051_decoder1_n146), .A1(
        oc8051_decoder1_n147), .B0(oc8051_decoder1_n148), .C0(
        oc8051_decoder1_n149), .Y(oc8051_decoder1_n143) );
  OAI222_X0P5M_A12TS oc8051_decoder1_u75 ( .A0(oc8051_decoder1_n123), .A1(
        oc8051_decoder1_n122), .B0(oc8051_decoder1_n143), .B1(
        oc8051_decoder1_n144), .C0(oc8051_decoder1_n125), .C1(
        oc8051_decoder1_n145), .Y(oc8051_decoder1_n423) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u74 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n138), .B1(op1_cur[0]), .C0(
        oc8051_decoder1_n142), .Y(oc8051_decoder1_n140) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u73 ( .A0(oc8051_decoder1_n139), .A1(
        op1_cur[1]), .B0(oc8051_decoder1_n140), .C0(oc8051_decoder1_n141), .Y(
        oc8051_decoder1_n129) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u72 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n138), .Y(
        oc8051_decoder1_n133) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u71 ( .A0(oc8051_decoder1_n135), .A1(
        oc8051_decoder1_n136), .B0(oc8051_decoder1_n42), .B1(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n134) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u70 ( .A(oc8051_decoder1_n132), .B(
        op1_cur[1]), .C(oc8051_decoder1_n133), .D(oc8051_decoder1_n134), .Y(
        oc8051_decoder1_n130) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u69 ( .A(oc8051_decoder1_n129), .B(
        oc8051_decoder1_n130), .S0(oc8051_decoder1_n131), .Y(
        oc8051_decoder1_n127) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u68 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n69), .A2(oc8051_decoder1_n127), .B0(
        oc8051_decoder1_n128), .Y(oc8051_decoder1_n120) );
  OA22_X0P5M_A12TS oc8051_decoder1_u67 ( .A0(oc8051_decoder1_n122), .A1(
        oc8051_decoder1_n123), .B0(oc8051_decoder1_n124), .B1(
        oc8051_decoder1_n125), .Y(oc8051_decoder1_n121) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u66 ( .A0(oc8051_decoder1_n118), .A1(
        oc8051_decoder1_n119), .B0(oc8051_decoder1_n120), .C0(
        oc8051_decoder1_n121), .Y(oc8051_decoder1_n424) );
  INV_X0P5B_A12TS oc8051_decoder1_u65 ( .A(wb_rst_i), .Y(oc8051_decoder1_n444)
         );
  NAND2_X0P5A_A12TS oc8051_decoder1_u64 ( .A(oc8051_decoder1_n117), .B(
        oc8051_decoder1_n33), .Y(oc8051_decoder1_n106) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u63 ( .A(oc8051_decoder1_n115), .B(
        oc8051_decoder1_n116), .Y(oc8051_decoder1_n72) );
  NAND3B_X0P5M_A12TS oc8051_decoder1_u62 ( .AN(oc8051_decoder1_n72), .B(
        oc8051_decoder1_n113), .C(oc8051_decoder1_n114), .Y(
        oc8051_decoder1_n96) );
  INV_X0P5B_A12TS oc8051_decoder1_u61 ( .A(oc8051_decoder1_n112), .Y(
        oc8051_decoder1_n94) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u60 ( .A0(oc8051_decoder1_n96), .A1(
        oc8051_decoder1_n94), .B0(oc8051_decoder1_n111), .Y(
        oc8051_decoder1_n107) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u59 ( .A(oc8051_decoder1_n68), .B(
        oc8051_decoder1_n75), .C(oc8051_decoder1_n110), .Y(oc8051_decoder1_n34) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u58 ( .A(oc8051_decoder1_n108), .B(
        oc8051_decoder1_n33), .C(oc8051_decoder1_n109), .Y(oc8051_decoder1_n89) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u57 ( .A(oc8051_decoder1_n106), .B(
        oc8051_decoder1_n107), .C(oc8051_decoder1_n34), .D(oc8051_decoder1_n89), .Y(pc_wr_sel[0]) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u56 ( .A(oc8051_decoder1_n59), .B(
        oc8051_decoder1_n105), .Y(oc8051_decoder1_n7) );
  INV_X0P5B_A12TS oc8051_decoder1_u55 ( .A(oc8051_decoder1_n104), .Y(
        oc8051_decoder1_n103) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u54 ( .A(oc8051_decoder1_n103), .B(
        oc8051_decoder1_n75), .Y(oc8051_decoder1_n87) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u53 ( .A0(oc8051_decoder1_n7), .A1(
        oc8051_decoder1_n14), .A2(oc8051_decoder1_n102), .B0(
        oc8051_decoder1_n87), .Y(oc8051_decoder1_n63) );
  INV_X0P5B_A12TS oc8051_decoder1_u52 ( .A(oc8051_decoder1_n63), .Y(
        oc8051_decoder1_n100) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u51 ( .A0(oc8051_decoder1_n5), .A1(
        oc8051_decoder1_n100), .B0(oc8051_decoder1_n29), .B1(
        oc8051_decoder1_n30), .C0(oc8051_decoder1_n101), .Y(
        oc8051_decoder1_n441) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u50 ( .A(oc8051_decoder1_n78), .B(
        oc8051_decoder1_n87), .C(oc8051_decoder1_n29), .Y(oc8051_decoder1_n93)
         );
  OAI21_X0P5M_A12TS oc8051_decoder1_u49 ( .A0(oc8051_decoder1_n98), .A1(
        oc8051_decoder1_n69), .B0(oc8051_decoder1_n99), .Y(oc8051_decoder1_n97) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u48 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n81), .B0(oc8051_decoder1_n96), .C0(
        oc8051_decoder1_n97), .Y(oc8051_decoder1_n95) );
  INV_X0P5B_A12TS oc8051_decoder1_u47 ( .A(oc8051_decoder1_n95), .Y(
        oc8051_decoder1_n86) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u46 ( .A(oc8051_decoder1_n93), .B(
        oc8051_decoder1_n86), .C(oc8051_decoder1_n94), .Y(oc8051_decoder1_n91)
         );
  OAI22_X0P5M_A12TS oc8051_decoder1_u45 ( .A0(oc8051_decoder1_n91), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n5), .B1(oc8051_decoder1_n92), .Y(pc_wr_sel[1]) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u44 ( .A(oc8051_decoder1_n90), .B(
        oc8051_decoder1_n33), .C(oc8051_decoder1_n44), .Y(oc8051_decoder1_n88)
         );
  OAI211_X0P5M_A12TS oc8051_decoder1_u43 ( .A0(oc8051_decoder1_n30), .A1(
        oc8051_decoder1_n87), .B0(oc8051_decoder1_n88), .C0(
        oc8051_decoder1_n89), .Y(pc_wr_sel[2]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u42 ( .A(oc8051_decoder1_n85), .B(
        oc8051_decoder1_n86), .Y(oc8051_decoder1_n79) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u41 ( .A0(oc8051_decoder1_n81), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n83), .C0(
        oc8051_decoder1_n84), .Y(oc8051_decoder1_n80) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u40 ( .A(oc8051_decoder1_n79), .B(
        oc8051_decoder1_n80), .S0(eq), .Y(oc8051_decoder1_n76) );
  INV_X0P5B_A12TS oc8051_decoder1_u39 ( .A(oc8051_decoder1_n78), .Y(
        oc8051_decoder1_n77) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u38 ( .A0(oc8051_decoder1_n68), .A1(
        oc8051_decoder1_n75), .B0(oc8051_decoder1_n76), .C0(
        oc8051_decoder1_n77), .Y(oc8051_decoder1_n73) );
  INV_X0P5B_A12TS oc8051_decoder1_u37 ( .A(pc_wr_sel[2]), .Y(
        oc8051_decoder1_n74) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u36 ( .A0(oc8051_decoder1_n73), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n34), .C0(
        oc8051_decoder1_n74), .Y(pc_wr) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u35 ( .A0(oc8051_decoder1_n70), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n67), .C0(
        oc8051_decoder1_n72), .Y(oc8051_decoder1_n64) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u34 ( .A0(oc8051_decoder1_n67), .A1(
        oc8051_decoder1_n21), .B0(oc8051_decoder1_n68), .B1(
        oc8051_decoder1_n69), .Y(oc8051_decoder1_n65) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u33 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n64), .B0(oc8051_decoder1_n65), .B1(
        oc8051_decoder1_n66), .Y(oc8051_decoder1_n62) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u32 ( .A0(oc8051_decoder1_n60), .A1(
        oc8051_decoder1_n61), .B0(oc8051_decoder1_n62), .C0(
        oc8051_decoder1_n63), .Y(oc8051_decoder1_n56) );
  AO21_X0P5M_A12TS oc8051_decoder1_u31 ( .A0(oc8051_decoder1_n58), .A1(
        oc8051_decoder1_n59), .B0(comp_sel[0]), .Y(oc8051_decoder1_n57) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u30 ( .A0(oc8051_decoder1_n5), .A1(
        oc8051_decoder1_n56), .B0(oc8051_decoder1_n57), .C0(
        oc8051_decoder1_n34), .Y(oc8051_decoder1_ram_rd_sel_0_) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u29 ( .A0(oc8051_decoder1_n53), .A1(
        op1_cur[0]), .B0(oc8051_decoder1_n54), .C0(oc8051_decoder1_n55), .Y(
        oc8051_decoder1_n15) );
  INV_X0P5B_A12TS oc8051_decoder1_u28 ( .A(oc8051_decoder1_n15), .Y(
        oc8051_decoder1_n51) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u27 ( .A0(oc8051_decoder1_n21), .A1(
        oc8051_decoder1_n22), .A2(oc8051_decoder1_n51), .B0(
        oc8051_decoder1_n52), .Y(oc8051_decoder1_n45) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u26 ( .A0(oc8051_decoder1_n47), .A1(
        oc8051_decoder1_n48), .B0(oc8051_decoder1_n49), .C0(
        oc8051_decoder1_n50), .Y(oc8051_decoder1_n46) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u25 ( .A0(oc8051_decoder1_n8), .A1(
        oc8051_decoder1_n40), .B0(oc8051_decoder1_n45), .C0(
        oc8051_decoder1_n46), .Y(oc8051_decoder1_n35) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u24 ( .A0(oc8051_decoder1_n42), .A1(
        oc8051_decoder1_n26), .B0(oc8051_decoder1_n27), .C0(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n43) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u23 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n41), .A2(oc8051_decoder1_n42), .B0(
        oc8051_decoder1_n43), .B1(oc8051_decoder1_n44), .Y(oc8051_decoder1_n39) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u22 ( .A0(oc8051_decoder1_n35), .A1(
        oc8051_decoder1_n36), .B0(oc8051_decoder1_n37), .B1(
        oc8051_decoder1_n38), .C0(oc8051_decoder1_n39), .Y(oc8051_decoder1_n32) );
  AOI21B_X0P5M_A12TS oc8051_decoder1_u21 ( .A0(oc8051_decoder1_n32), .A1(
        oc8051_decoder1_n33), .B0N(oc8051_decoder1_n34), .Y(
        oc8051_decoder1_n31) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u20 ( .A0(oc8051_decoder1_n29), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n31), .Y(
        oc8051_decoder1_ram_rd_sel_1_) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u19 ( .A(oc8051_decoder1_ram_rd_sel_0_), 
        .B(oc8051_decoder1_ram_rd_sel_r[0]), .S0(wait_data), .Y(ram_rd_sel[0])
         );
  MXT2_X0P5M_A12TS oc8051_decoder1_u18 ( .A(oc8051_decoder1_ram_rd_sel_1_), 
        .B(oc8051_decoder1_ram_rd_sel_r[1]), .S0(wait_data), .Y(ram_rd_sel[1])
         );
  MXT2_X0P5M_A12TS oc8051_decoder1_u17 ( .A(oc8051_decoder1_n441), .B(
        oc8051_decoder1_ram_rd_sel_r[2]), .S0(wait_data), .Y(ram_rd_sel[2]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u16 ( .A(wait_data), .B(oc8051_decoder1_n28), .Y(ram_wr_sel[0]) );
  NOR2B_X0P5M_A12TS oc8051_decoder1_u15 ( .AN(oc8051_decoder1_ram_wr_sel_1_), 
        .B(wait_data), .Y(ram_wr_sel[1]) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u14 ( .A0(oc8051_decoder1_n25), .A1(
        oc8051_decoder1_n26), .A2(oc8051_decoder1_n11), .B0(
        oc8051_decoder1_n27), .Y(oc8051_decoder1_n17) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u13 ( .A0(oc8051_decoder1_n21), .A1(
        oc8051_decoder1_n22), .A2(oc8051_decoder1_n23), .B0(
        oc8051_decoder1_n24), .Y(oc8051_decoder1_n19) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u12 ( .A0(oc8051_decoder1_n17), .A1(
        oc8051_decoder1_n18), .A2(oc8051_decoder1_n19), .B0(
        oc8051_decoder1_n20), .Y(oc8051_decoder1_n2) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u11 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n15), .C(oc8051_decoder1_n16), .Y(oc8051_decoder1_n3)
         );
  NAND3_X0P5A_A12TS oc8051_decoder1_u10 ( .A(oc8051_decoder1_n11), .B(
        oc8051_decoder1_n12), .C(oc8051_decoder1_n13), .Y(oc8051_decoder1_n10)
         );
  AOI32_X0P5M_A12TS oc8051_decoder1_u9 ( .A0(oc8051_decoder1_n6), .A1(
        oc8051_decoder1_n7), .A2(oc8051_decoder1_n8), .B0(oc8051_decoder1_n9), 
        .B1(oc8051_decoder1_n10), .Y(oc8051_decoder1_n4) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u8 ( .A(wait_data), .B(oc8051_decoder1_n1), 
        .Y(wr_o) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u7 ( .A(wait_data), .B(oc8051_decoder1_n407), .Y(wr_sfr[0]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u6 ( .A(wait_data), .B(oc8051_decoder1_n406), .Y(wr_sfr[1]) );
  AOI31_X2M_A12TS oc8051_decoder1_u5 ( .A0(oc8051_decoder1_n2), .A1(
        oc8051_decoder1_n3), .A2(oc8051_decoder1_n4), .B0(oc8051_decoder1_n5), 
        .Y(rmw) );
  OAI22_X2M_A12TS oc8051_decoder1_u4 ( .A0(oc8051_decoder1_n318), .A1(
        oc8051_decoder1_n301), .B0(oc8051_decoder1_n439), .B1(
        oc8051_decoder1_n302), .Y(op1_cur[0]) );
  NOR2_X1M_A12TS oc8051_decoder1_u3 ( .A(wait_data), .B(oc8051_decoder1_n408), 
        .Y(ram_wr_sel[2]) );
  DFFRPQN_X1M_A12TS oc8051_decoder1_ram_wr_sel_reg_2_ ( .D(
        oc8051_decoder1_n412), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_decoder1_n408) );
  DFFRPQN_X1M_A12TS oc8051_decoder1_wr_sfr_reg_0_ ( .D(oc8051_decoder1_n414), 
        .CK(wb_clk_i), .R(wb_rst_i), .QN(oc8051_decoder1_n407) );
  DFFRPQN_X1M_A12TS oc8051_decoder1_wr_sfr_reg_1_ ( .D(oc8051_decoder1_n413), 
        .CK(wb_clk_i), .R(wb_rst_i), .QN(oc8051_decoder1_n406) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel3_reg ( .D(oc8051_decoder1_n394), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel3) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel1_reg_0_ ( .D(oc8051_decoder1_n417), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel1[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel1_reg_1_ ( .D(oc8051_decoder1_n416), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel1[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel1_reg_2_ ( .D(oc8051_decoder1_n415), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel1[2]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_psw_set_reg_1_ ( .D(oc8051_decoder1_n420), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(psw_set[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel2_reg_0_ ( .D(oc8051_decoder1_n390), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel2[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel2_reg_1_ ( .D(oc8051_decoder1_n392), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel2[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_psw_set_reg_0_ ( .D(oc8051_decoder1_n389), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(psw_set[0]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_state_reg_0_ ( .D(oc8051_decoder1_n405), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(oc8051_decoder1_state_0_)
         );
  DFFRPQ_X1M_A12TS oc8051_decoder1_cy_sel_reg_0_ ( .D(oc8051_decoder1_n391), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(cy_sel[0]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_state_reg_1_ ( .D(oc8051_decoder1_n395), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(oc8051_decoder1_state_1_)
         );
  DFFRPQ_X1M_A12TS oc8051_decoder1_cy_sel_reg_1_ ( .D(oc8051_decoder1_n393), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(cy_sel[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_wr_sel_reg_1_ ( .D(oc8051_decoder1_n418), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_ram_wr_sel_1_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_2_ ( .D(oc8051_decoder1_n422), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_2_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_3_ ( .D(oc8051_decoder1_n388), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_3_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_0_ ( .D(oc8051_decoder1_n424), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_0_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_1_ ( .D(oc8051_decoder1_n423), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_1_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_wr_reg ( .D(oc8051_decoder1_n421), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_wr) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_wr_sel_reg_0_ ( .D(oc8051_decoder1_n419), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_ram_wr_sel_0_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_7_ ( .D(oc8051_decoder1_n396), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[7]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_6_ ( .D(oc8051_decoder1_n397), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[6]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_5_ ( .D(oc8051_decoder1_n398), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[5]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_4_ ( .D(oc8051_decoder1_n399), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[4]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_3_ ( .D(oc8051_decoder1_n400), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[3]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_2_ ( .D(oc8051_decoder1_n401), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[2]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_1_ ( .D(oc8051_decoder1_n402), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_0_ ( .D(oc8051_decoder1_n403), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_rd_sel_r_reg_0_ ( .D(
        oc8051_decoder1_ram_rd_sel_0_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_decoder1_ram_rd_sel_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_rd_sel_r_reg_1_ ( .D(
        oc8051_decoder1_ram_rd_sel_1_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_decoder1_ram_rd_sel_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_rd_sel_r_reg_2_ ( .D(
        oc8051_decoder1_n441), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_decoder1_ram_rd_sel_r[2]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_mem_act_reg_1_ ( .D(oc8051_decoder1_n1805), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(mem_act[1]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_mem_act_reg_0_ ( .D(oc8051_decoder1_n1804), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(mem_act[0]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_mem_act_reg_2_ ( .D(oc8051_decoder1_n1806), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(mem_act[2]) );
  INV_X0P5B_A12TS oc8051_alu1_u297 ( .A(alu_op[2]), .Y(oc8051_alu1_n220) );
  AND2_X0P5M_A12TS oc8051_alu1_u296 ( .A(alu_op[3]), .B(oc8051_alu1_n220), .Y(
        oc8051_alu1_n205) );
  INV_X0P5B_A12TS oc8051_alu1_u295 ( .A(alu_op[0]), .Y(oc8051_alu1_n221) );
  AND2_X0P5M_A12TS oc8051_alu1_u294 ( .A(alu_op[1]), .B(oc8051_alu1_n221), .Y(
        oc8051_alu1_n206) );
  NAND2_X0P5A_A12TS oc8051_alu1_u293 ( .A(oc8051_alu1_n205), .B(
        oc8051_alu1_n206), .Y(oc8051_alu1_n42) );
  INV_X0P5B_A12TS oc8051_alu1_u292 ( .A(src1[7]), .Y(oc8051_alu1_n87) );
  INV_X0P5B_A12TS oc8051_alu1_u291 ( .A(src1[1]), .Y(oc8051_alu1_n195) );
  AND2_X0P5M_A12TS oc8051_alu1_u290 ( .A(alu_op[3]), .B(alu_op[2]), .Y(
        oc8051_alu1_n214) );
  NOR2_X0P5A_A12TS oc8051_alu1_u289 ( .A(alu_op[1]), .B(alu_op[0]), .Y(
        oc8051_alu1_n208) );
  NAND2_X0P5A_A12TS oc8051_alu1_u288 ( .A(oc8051_alu1_n214), .B(
        oc8051_alu1_n208), .Y(oc8051_alu1_n46) );
  INV_X0P5B_A12TS oc8051_alu1_u287 ( .A(oc8051_alu1_n46), .Y(oc8051_alu1_n142)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_u286 ( .A(oc8051_alu1_n221), .B(alu_op[1]), .Y(
        oc8051_alu1_n216) );
  NAND2_X0P5A_A12TS oc8051_alu1_u285 ( .A(oc8051_alu1_n214), .B(
        oc8051_alu1_n216), .Y(oc8051_alu1_n139) );
  INV_X0P5B_A12TS oc8051_alu1_u284 ( .A(oc8051_alu1_n139), .Y(oc8051_alu1_n53)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_u283 ( .A(oc8051_alu1_n142), .B(oc8051_alu1_n53), .Y(oc8051_alu1_n109) );
  NOR2_X0P5A_A12TS oc8051_alu1_u282 ( .A(oc8051_alu1_n220), .B(alu_op[3]), .Y(
        oc8051_alu1_n207) );
  NAND2_X0P5A_A12TS oc8051_alu1_u281 ( .A(oc8051_alu1_n216), .B(
        oc8051_alu1_n207), .Y(oc8051_alu1_n111) );
  INV_X0P5B_A12TS oc8051_alu1_u280 ( .A(oc8051_alu1_n111), .Y(oc8051_alu1_n52)
         );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u279 ( .A0(src1[2]), .A1(src1[1]), .B0(
        src1[3]), .C0(srcac), .Y(oc8051_alu1_n117) );
  NOR2_X0P5A_A12TS oc8051_alu1_u278 ( .A(alu_op[3]), .B(alu_op[2]), .Y(
        oc8051_alu1_n204) );
  NAND2_X0P5A_A12TS oc8051_alu1_u277 ( .A(oc8051_alu1_n204), .B(
        oc8051_alu1_n208), .Y(oc8051_alu1_n43) );
  AO1B2_X0P5M_A12TS oc8051_alu1_u276 ( .B0(oc8051_alu1_n52), .B1(
        oc8051_alu1_n117), .A0N(oc8051_alu1_n43), .Y(oc8051_alu1_n172) );
  NOR2_X0P5A_A12TS oc8051_alu1_u275 ( .A(oc8051_alu1_n111), .B(
        oc8051_alu1_n117), .Y(oc8051_alu1_n50) );
  OAI21_X0P5M_A12TS oc8051_alu1_u274 ( .A0(oc8051_alu1_n172), .A1(
        oc8051_alu1_n50), .B0(src1[0]), .Y(oc8051_alu1_n219) );
  OAI221_X0P5M_A12TS oc8051_alu1_u273 ( .A0(oc8051_alu1_n42), .A1(
        oc8051_alu1_n87), .B0(oc8051_alu1_n195), .B1(oc8051_alu1_n109), .C0(
        oc8051_alu1_n219), .Y(oc8051_alu1_n197) );
  NAND2_X0P5A_A12TS oc8051_alu1_u272 ( .A(oc8051_alu1_n204), .B(
        oc8051_alu1_n216), .Y(oc8051_alu1_n23) );
  INV_X0P5B_A12TS oc8051_alu1_u271 ( .A(oc8051_alu1_n23), .Y(oc8051_alu1_n223)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_u270 ( .A(oc8051_alu1_n206), .B(
        oc8051_alu1_n207), .Y(oc8051_alu1_n40) );
  INV_X0P5B_A12TS oc8051_alu1_u269 ( .A(oc8051_alu1_n40), .Y(oc8051_alu1_n224)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_u268 ( .A(oc8051_alu1_n205), .B(
        oc8051_alu1_n208), .Y(oc8051_alu1_n122) );
  NAND2_X0P5A_A12TS oc8051_alu1_u267 ( .A(oc8051_alu1_n205), .B(
        oc8051_alu1_n216), .Y(oc8051_alu1_n12) );
  OAI21_X0P5M_A12TS oc8051_alu1_u266 ( .A0(src2[0]), .A1(oc8051_alu1_n122), 
        .B0(oc8051_alu1_n12), .Y(oc8051_alu1_n215) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u265 ( .A(oc8051_alu1_n224), .B(
        oc8051_alu1_n215), .S0(src1[0]), .Y(oc8051_alu1_n209) );
  AND3_X0P5M_A12TS oc8051_alu1_u264 ( .A(oc8051_alu1_n206), .B(alu_cy), .C(
        oc8051_alu1_n214), .Y(oc8051_alu1_n138) );
  NAND2_X0P5A_A12TS oc8051_alu1_u263 ( .A(oc8051_alu1_dec[0]), .B(
        oc8051_alu1_n138), .Y(oc8051_alu1_n210) );
  INV_X0P5B_A12TS oc8051_alu1_u262 ( .A(alu_cy), .Y(
        oc8051_alu1_sub_1_root_sub_189_2_carry_0_) );
  AND3_X0P5M_A12TS oc8051_alu1_u261 ( .A(oc8051_alu1_n206), .B(
        oc8051_alu1_sub_1_root_sub_189_2_carry_0_), .C(oc8051_alu1_n214), .Y(
        oc8051_alu1_n137) );
  NAND2_X0P5A_A12TS oc8051_alu1_u260 ( .A(oc8051_alu1_inc[0]), .B(
        oc8051_alu1_n137), .Y(oc8051_alu1_n211) );
  AND2_X0P5M_A12TS oc8051_alu1_u259 ( .A(alu_op[1]), .B(alu_op[0]), .Y(
        oc8051_alu1_n201) );
  NAND2_X0P5A_A12TS oc8051_alu1_u258 ( .A(oc8051_alu1_n214), .B(
        oc8051_alu1_n201), .Y(oc8051_alu1_n136) );
  INV_X0P5B_A12TS oc8051_alu1_u257 ( .A(oc8051_alu1_n136), .Y(oc8051_alu1_n79)
         );
  INV_X0P5B_A12TS oc8051_alu1_u256 ( .A(oc8051_alu1_n12), .Y(oc8051_alu1_n48)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_u255 ( .A(oc8051_alu1_n79), .B(oc8051_alu1_n48), 
        .Y(oc8051_alu1_n247) );
  INV_X0P5B_A12TS oc8051_alu1_u254 ( .A(oc8051_alu1_n247), .Y(oc8051_alu1_n103) );
  NAND2_X0P5A_A12TS oc8051_alu1_u253 ( .A(oc8051_alu1_n201), .B(
        oc8051_alu1_n207), .Y(oc8051_alu1_n124) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u252 ( .A(oc8051_alu1_n122), .B(
        oc8051_alu1_n124), .S0(src1[0]), .Y(oc8051_alu1_n213) );
  OAI21_X0P5M_A12TS oc8051_alu1_u251 ( .A0(oc8051_alu1_n103), .A1(
        oc8051_alu1_n213), .B0(src2[0]), .Y(oc8051_alu1_n212) );
  NAND4_X0P5A_A12TS oc8051_alu1_u250 ( .A(oc8051_alu1_n209), .B(
        oc8051_alu1_n210), .C(oc8051_alu1_n211), .D(oc8051_alu1_n212), .Y(
        oc8051_alu1_n107) );
  AOI21_X0P5M_A12TS oc8051_alu1_u249 ( .A0(oc8051_alu1_add4_0_), .A1(
        oc8051_alu1_n223), .B0(oc8051_alu1_n107), .Y(oc8051_alu1_n198) );
  NAND2_X0P5A_A12TS oc8051_alu1_u248 ( .A(oc8051_alu1_n207), .B(
        oc8051_alu1_n208), .Y(oc8051_alu1_n113) );
  INV_X0P5B_A12TS oc8051_alu1_u247 ( .A(oc8051_alu1_n113), .Y(oc8051_alu1_n222) );
  NAND2_X0P5A_A12TS oc8051_alu1_u246 ( .A(oc8051_alu1_n206), .B(
        oc8051_alu1_n204), .Y(oc8051_alu1_n22) );
  INV_X0P5B_A12TS oc8051_alu1_u245 ( .A(oc8051_alu1_n22), .Y(oc8051_alu1_n49)
         );
  AOI22_X0P5M_A12TS oc8051_alu1_u244 ( .A0(oc8051_alu1_divsrc1[0]), .A1(
        oc8051_alu1_n222), .B0(sub_result[0]), .B1(oc8051_alu1_n49), .Y(
        oc8051_alu1_n199) );
  AND2_X0P5M_A12TS oc8051_alu1_u243 ( .A(oc8051_alu1_n205), .B(
        oc8051_alu1_n201), .Y(oc8051_alu1_n33) );
  NAND2_X0P5A_A12TS oc8051_alu1_u242 ( .A(oc8051_alu1_n201), .B(
        oc8051_alu1_n204), .Y(oc8051_alu1_n112) );
  INV_X0P5B_A12TS oc8051_alu1_u241 ( .A(oc8051_alu1_n112), .Y(oc8051_alu1_n225) );
  AOI22_X0P5M_A12TS oc8051_alu1_u240 ( .A0(oc8051_alu1_n33), .A1(alu_cy), .B0(
        oc8051_alu1_mulsrc1[0]), .B1(oc8051_alu1_n225), .Y(oc8051_alu1_n200)
         );
  NAND4B_X0P5M_A12TS oc8051_alu1_u239 ( .AN(oc8051_alu1_n197), .B(
        oc8051_alu1_n198), .C(oc8051_alu1_n199), .D(oc8051_alu1_n200), .Y(
        oc8051_alu1_n2130) );
  OAI21_X0P5M_A12TS oc8051_alu1_u238 ( .A0(src2[1]), .A1(oc8051_alu1_n122), 
        .B0(oc8051_alu1_n12), .Y(oc8051_alu1_n196) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u237 ( .A(oc8051_alu1_n196), .B(
        oc8051_alu1_n224), .S0(oc8051_alu1_n195), .Y(oc8051_alu1_n190) );
  NAND2_X0P5A_A12TS oc8051_alu1_u236 ( .A(oc8051_alu1_dec[1]), .B(
        oc8051_alu1_n138), .Y(oc8051_alu1_n191) );
  NAND2_X0P5A_A12TS oc8051_alu1_u235 ( .A(oc8051_alu1_inc[1]), .B(
        oc8051_alu1_n137), .Y(oc8051_alu1_n192) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u234 ( .A(oc8051_alu1_n124), .B(
        oc8051_alu1_n122), .S0(oc8051_alu1_n195), .Y(oc8051_alu1_n194) );
  OAI21_X0P5M_A12TS oc8051_alu1_u233 ( .A0(oc8051_alu1_n103), .A1(
        oc8051_alu1_n194), .B0(src2[1]), .Y(oc8051_alu1_n193) );
  NAND4_X0P5A_A12TS oc8051_alu1_u232 ( .A(oc8051_alu1_n190), .B(
        oc8051_alu1_n191), .C(oc8051_alu1_n192), .D(oc8051_alu1_n193), .Y(
        oc8051_alu1_n106) );
  AOI21_X0P5M_A12TS oc8051_alu1_u231 ( .A0(oc8051_alu1_add4_1_), .A1(
        oc8051_alu1_n223), .B0(oc8051_alu1_n106), .Y(oc8051_alu1_n186) );
  AOI22_X0P5M_A12TS oc8051_alu1_u230 ( .A0(oc8051_alu1_divsrc1[1]), .A1(
        oc8051_alu1_n222), .B0(sub_result[1]), .B1(oc8051_alu1_n49), .Y(
        oc8051_alu1_n187) );
  INV_X0P5B_A12TS oc8051_alu1_u229 ( .A(oc8051_alu1_n109), .Y(oc8051_alu1_n152) );
  AOI22_X0P5M_A12TS oc8051_alu1_u228 ( .A0(src1[2]), .A1(oc8051_alu1_n152), 
        .B0(oc8051_alu1_mulsrc1[1]), .B1(oc8051_alu1_n225), .Y(
        oc8051_alu1_n188) );
  INV_X0P5B_A12TS oc8051_alu1_u227 ( .A(oc8051_alu1_n42), .Y(oc8051_alu1_n47)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_u226 ( .A(oc8051_alu1_n33), .B(oc8051_alu1_n47), 
        .Y(oc8051_alu1_n110) );
  INV_X0P5B_A12TS oc8051_alu1_u225 ( .A(oc8051_alu1_n110), .Y(oc8051_alu1_n143) );
  AOI222_X0P5M_A12TS oc8051_alu1_u224 ( .A0(oc8051_alu1_n195), .A1(
        oc8051_alu1_n50), .B0(src1[0]), .B1(oc8051_alu1_n143), .C0(src1[1]), 
        .C1(oc8051_alu1_n172), .Y(oc8051_alu1_n189) );
  NAND4_X0P5A_A12TS oc8051_alu1_u223 ( .A(oc8051_alu1_n186), .B(
        oc8051_alu1_n187), .C(oc8051_alu1_n188), .D(oc8051_alu1_n189), .Y(
        oc8051_alu1_n2140) );
  OAI21_X0P5M_A12TS oc8051_alu1_u222 ( .A0(src2[2]), .A1(oc8051_alu1_n122), 
        .B0(oc8051_alu1_n12), .Y(oc8051_alu1_n185) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u221 ( .A(oc8051_alu1_n224), .B(
        oc8051_alu1_n185), .S0(src1[2]), .Y(oc8051_alu1_n180) );
  NAND2_X0P5A_A12TS oc8051_alu1_u220 ( .A(oc8051_alu1_dec[2]), .B(
        oc8051_alu1_n138), .Y(oc8051_alu1_n181) );
  NAND2_X0P5A_A12TS oc8051_alu1_u219 ( .A(oc8051_alu1_inc[2]), .B(
        oc8051_alu1_n137), .Y(oc8051_alu1_n182) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u218 ( .A(oc8051_alu1_n122), .B(
        oc8051_alu1_n124), .S0(src1[2]), .Y(oc8051_alu1_n184) );
  OAI21_X0P5M_A12TS oc8051_alu1_u217 ( .A0(oc8051_alu1_n103), .A1(
        oc8051_alu1_n184), .B0(src2[2]), .Y(oc8051_alu1_n183) );
  NAND4_X0P5A_A12TS oc8051_alu1_u216 ( .A(oc8051_alu1_n180), .B(
        oc8051_alu1_n181), .C(oc8051_alu1_n182), .D(oc8051_alu1_n183), .Y(
        oc8051_alu1_n105) );
  AOI21_X0P5M_A12TS oc8051_alu1_u215 ( .A0(oc8051_alu1_add4_2_), .A1(
        oc8051_alu1_n223), .B0(oc8051_alu1_n105), .Y(oc8051_alu1_n173) );
  AOI22_X0P5M_A12TS oc8051_alu1_u214 ( .A0(oc8051_alu1_divsrc1[2]), .A1(
        oc8051_alu1_n222), .B0(sub_result[2]), .B1(oc8051_alu1_n49), .Y(
        oc8051_alu1_n177) );
  AOI22_X0P5M_A12TS oc8051_alu1_u213 ( .A0(oc8051_alu1_n152), .A1(src1[3]), 
        .B0(oc8051_alu1_mulsrc1[2]), .B1(oc8051_alu1_n225), .Y(
        oc8051_alu1_n178) );
  AOI222_X0P5M_A12TS oc8051_alu1_u212 ( .A0(oc8051_alu1_n1510), .A1(
        oc8051_alu1_n50), .B0(src1[1]), .B1(oc8051_alu1_n143), .C0(src1[2]), 
        .C1(oc8051_alu1_n172), .Y(oc8051_alu1_n179) );
  NAND4_X0P5A_A12TS oc8051_alu1_u211 ( .A(oc8051_alu1_n173), .B(
        oc8051_alu1_n177), .C(oc8051_alu1_n178), .D(oc8051_alu1_n179), .Y(
        oc8051_alu1_n2150) );
  AOI22_X0P5M_A12TS oc8051_alu1_u210 ( .A0(sub_result[3]), .A1(oc8051_alu1_n49), .B0(oc8051_alu1_add4_3_), .B1(oc8051_alu1_n223), .Y(oc8051_alu1_n168) );
  AOI22_X0P5M_A12TS oc8051_alu1_u209 ( .A0(oc8051_alu1_mulsrc1[3]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc1[3]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n169) );
  AOI22_X0P5M_A12TS oc8051_alu1_u208 ( .A0(oc8051_alu1_n1520), .A1(
        oc8051_alu1_n50), .B0(src1[4]), .B1(oc8051_alu1_n152), .Y(
        oc8051_alu1_n170) );
  NAND2_X0P5A_A12TS oc8051_alu1_u207 ( .A(oc8051_alu1_n244), .B(
        oc8051_alu1_n243), .Y(oc8051_alu1_n176) );
  AOI221_X0P5M_A12TS oc8051_alu1_u206 ( .A0(oc8051_alu1_n172), .A1(src1[3]), 
        .B0(src1[2]), .B1(oc8051_alu1_n143), .C0(oc8051_alu1_n176), .Y(
        oc8051_alu1_n171) );
  NAND4_X0P5A_A12TS oc8051_alu1_u205 ( .A(oc8051_alu1_n168), .B(
        oc8051_alu1_n169), .C(oc8051_alu1_n170), .D(oc8051_alu1_n171), .Y(
        oc8051_alu1_n2160) );
  INV_X0P5B_A12TS oc8051_alu1_u204 ( .A(src2[4]), .Y(oc8051_alu1_n15) );
  INV_X0P5B_A12TS oc8051_alu1_u203 ( .A(src1[4]), .Y(oc8051_alu1_n102) );
  NOR2_X0P5A_A12TS oc8051_alu1_u202 ( .A(oc8051_alu1_n15), .B(oc8051_alu1_n102), .Y(oc8051_alu1_n160) );
  INV_X0P5B_A12TS oc8051_alu1_u201 ( .A(oc8051_alu1_n160), .Y(oc8051_alu1_n16)
         );
  OAI21_X0P5M_A12TS oc8051_alu1_u200 ( .A0(src2[4]), .A1(src1[4]), .B0(
        oc8051_alu1_n16), .Y(oc8051_alu1_n167) );
  INV_X0P5B_A12TS oc8051_alu1_u199 ( .A(oc8051_alu1_sub4_4_), .Y(
        oc8051_alu1_n55) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u198 ( .A(oc8051_alu1_n167), .B(
        oc8051_alu1_n55), .Y(sub_result[4]) );
  OAI221_X0P5M_A12TS oc8051_alu1_u197 ( .A0(oc8051_alu1_n122), .A1(
        oc8051_alu1_n167), .B0(src1[4]), .B1(oc8051_alu1_n40), .C0(
        oc8051_alu1_n236), .Y(oc8051_alu1_n104) );
  AOI21_X0P5M_A12TS oc8051_alu1_u196 ( .A0(sub_result[4]), .A1(oc8051_alu1_n49), .B0(oc8051_alu1_n104), .Y(oc8051_alu1_n162) );
  AOI22_X0P5M_A12TS oc8051_alu1_u195 ( .A0(oc8051_alu1_mulsrc1[4]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc1[4]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n163) );
  AOI22_X0P5M_A12TS oc8051_alu1_u194 ( .A0(oc8051_alu1_n1770), .A1(
        oc8051_alu1_n52), .B0(src1[5]), .B1(oc8051_alu1_n152), .Y(
        oc8051_alu1_n164) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u193 ( .A(oc8051_alu1_add4_4_), .B(
        oc8051_alu1_n167), .Y(oc8051_alu1_n166) );
  OAI21_X0P5M_A12TS oc8051_alu1_u192 ( .A0(alu_cy), .A1(oc8051_alu1_n136), 
        .B0(oc8051_alu1_n43), .Y(oc8051_alu1_n61) );
  NOR2_X0P5A_A12TS oc8051_alu1_u191 ( .A(oc8051_alu1_n61), .B(oc8051_alu1_n48), 
        .Y(oc8051_alu1_n125) );
  INV_X0P5B_A12TS oc8051_alu1_u190 ( .A(oc8051_alu1_n125), .Y(oc8051_alu1_n149) );
  AOI222_X0P5M_A12TS oc8051_alu1_u189 ( .A0(oc8051_alu1_n143), .A1(src1[3]), 
        .B0(oc8051_alu1_n223), .B1(oc8051_alu1_n166), .C0(src1[4]), .C1(
        oc8051_alu1_n149), .Y(oc8051_alu1_n165) );
  NAND4_X0P5A_A12TS oc8051_alu1_u188 ( .A(oc8051_alu1_n162), .B(
        oc8051_alu1_n163), .C(oc8051_alu1_n164), .D(oc8051_alu1_n165), .Y(
        oc8051_alu1_n2170) );
  NAND2_X0P5A_A12TS oc8051_alu1_u187 ( .A(src2[5]), .B(src1[5]), .Y(
        oc8051_alu1_n18) );
  OAI21_X0P5M_A12TS oc8051_alu1_u186 ( .A0(src2[5]), .A1(src1[5]), .B0(
        oc8051_alu1_n18), .Y(oc8051_alu1_n159) );
  NAND2_X0P5A_A12TS oc8051_alu1_u185 ( .A(oc8051_alu1_n15), .B(src1[4]), .Y(
        oc8051_alu1_n161) );
  AOI22_X0P5M_A12TS oc8051_alu1_u184 ( .A0(oc8051_alu1_n102), .A1(src2[4]), 
        .B0(oc8051_alu1_n55), .B1(oc8051_alu1_n161), .Y(oc8051_alu1_n153) );
  XOR2_X0P5M_A12TS oc8051_alu1_u183 ( .A(oc8051_alu1_n159), .B(
        oc8051_alu1_n153), .Y(sub_result[5]) );
  OAI221_X0P5M_A12TS oc8051_alu1_u182 ( .A0(oc8051_alu1_n122), .A1(
        oc8051_alu1_n159), .B0(src1[5]), .B1(oc8051_alu1_n40), .C0(
        oc8051_alu1_n227), .Y(oc8051_alu1_n100) );
  AOI21_X0P5M_A12TS oc8051_alu1_u181 ( .A0(sub_result[5]), .A1(oc8051_alu1_n49), .B0(oc8051_alu1_n100), .Y(oc8051_alu1_n154) );
  AOI22_X0P5M_A12TS oc8051_alu1_u180 ( .A0(oc8051_alu1_mulsrc1[5]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc1[5]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n155) );
  AOI22_X0P5M_A12TS oc8051_alu1_u179 ( .A0(oc8051_alu1_n1780), .A1(
        oc8051_alu1_n52), .B0(src1[6]), .B1(oc8051_alu1_n152), .Y(
        oc8051_alu1_n156) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u178 ( .A0(src2[4]), .A1(src1[4]), .B0(
        oc8051_alu1_add4_4_), .C0(oc8051_alu1_n160), .Y(oc8051_alu1_n151) );
  XOR2_X0P5M_A12TS oc8051_alu1_u177 ( .A(oc8051_alu1_n151), .B(
        oc8051_alu1_n159), .Y(oc8051_alu1_n158) );
  AOI222_X0P5M_A12TS oc8051_alu1_u176 ( .A0(src1[4]), .A1(oc8051_alu1_n143), 
        .B0(oc8051_alu1_n158), .B1(oc8051_alu1_n223), .C0(src1[5]), .C1(
        oc8051_alu1_n149), .Y(oc8051_alu1_n157) );
  NAND4_X0P5A_A12TS oc8051_alu1_u175 ( .A(oc8051_alu1_n154), .B(
        oc8051_alu1_n155), .C(oc8051_alu1_n156), .D(oc8051_alu1_n157), .Y(
        oc8051_alu1_n2180) );
  INV_X0P5B_A12TS oc8051_alu1_u174 ( .A(src2[5]), .Y(oc8051_alu1_n17) );
  CGENI_X1M_A12TS oc8051_alu1_u173 ( .A(src1[5]), .B(oc8051_alu1_n17), .CI(
        oc8051_alu1_n153), .CON(oc8051_alu1_n131) );
  INV_X0P5B_A12TS oc8051_alu1_u172 ( .A(src1[6]), .Y(oc8051_alu1_n19) );
  XOR2_X0P5M_A12TS oc8051_alu1_u171 ( .A(src2[6]), .B(oc8051_alu1_n19), .Y(
        oc8051_alu1_n150) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u170 ( .A(oc8051_alu1_n131), .B(
        oc8051_alu1_n150), .Y(sub_result[6]) );
  OAI221_X0P5M_A12TS oc8051_alu1_u169 ( .A0(oc8051_alu1_n122), .A1(
        oc8051_alu1_n150), .B0(src1[6]), .B1(oc8051_alu1_n40), .C0(
        oc8051_alu1_n217), .Y(oc8051_alu1_n97) );
  AOI21_X0P5M_A12TS oc8051_alu1_u168 ( .A0(oc8051_alu1_n49), .A1(sub_result[6]), .B0(oc8051_alu1_n97), .Y(oc8051_alu1_n144) );
  AOI22_X0P5M_A12TS oc8051_alu1_u167 ( .A0(oc8051_alu1_mulsrc1[6]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc1[6]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n145) );
  AOI22_X0P5M_A12TS oc8051_alu1_u166 ( .A0(oc8051_alu1_n1790), .A1(
        oc8051_alu1_n52), .B0(oc8051_alu1_n152), .B1(src1[7]), .Y(
        oc8051_alu1_n146) );
  INV_X0P5B_A12TS oc8051_alu1_u165 ( .A(src1[5]), .Y(oc8051_alu1_n99) );
  AO21A1AI2_X0P5M_A12TS oc8051_alu1_u164 ( .A0(oc8051_alu1_n17), .A1(
        oc8051_alu1_n99), .B0(oc8051_alu1_n151), .C0(oc8051_alu1_n18), .Y(
        oc8051_alu1_n126) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u163 ( .A(oc8051_alu1_n126), .B(
        oc8051_alu1_n150), .Y(oc8051_alu1_n148) );
  AOI222_X0P5M_A12TS oc8051_alu1_u161 ( .A0(src1[5]), .A1(oc8051_alu1_n143), 
        .B0(oc8051_alu1_n148), .B1(oc8051_alu1_n223), .C0(src1[6]), .C1(
        oc8051_alu1_n149), .Y(oc8051_alu1_n147) );
  NAND4_X0P5A_A12TS oc8051_alu1_u158 ( .A(oc8051_alu1_n144), .B(
        oc8051_alu1_n145), .C(oc8051_alu1_n146), .D(oc8051_alu1_n147), .Y(
        oc8051_alu1_n2190) );
  AOI22_X0P5M_A12TS oc8051_alu1_u157 ( .A0(src1[6]), .A1(oc8051_alu1_n143), 
        .B0(oc8051_alu1_n1800), .B1(oc8051_alu1_n52), .Y(oc8051_alu1_n140) );
  AOI22_X0P5M_A12TS oc8051_alu1_u156 ( .A0(oc8051_alu1_n142), .A1(src1[0]), 
        .B0(oc8051_alu1_mulsrc1[7]), .B1(oc8051_alu1_n225), .Y(
        oc8051_alu1_n141) );
  OAI211_X0P5M_A12TS oc8051_alu1_u155 ( .A0(
        oc8051_alu1_sub_1_root_sub_189_2_carry_0_), .A1(oc8051_alu1_n139), 
        .B0(oc8051_alu1_n140), .C0(oc8051_alu1_n141), .Y(oc8051_alu1_n118) );
  INV_X0P5B_A12TS oc8051_alu1_u154 ( .A(oc8051_alu1_n124), .Y(oc8051_alu1_n45)
         );
  INV_X0P5B_A12TS oc8051_alu1_u153 ( .A(oc8051_alu1_n122), .Y(oc8051_alu1_n39)
         );
  MXIT2_X0P5M_A12TS oc8051_alu1_u152 ( .A(oc8051_alu1_n45), .B(oc8051_alu1_n39), .S0(oc8051_alu1_n87), .Y(oc8051_alu1_n135) );
  NOR2_X0P5A_A12TS oc8051_alu1_u151 ( .A(oc8051_alu1_n136), .B(
        oc8051_alu1_sub_1_root_sub_189_2_carry_0_), .Y(oc8051_alu1_n62) );
  NOR2_X0P5A_A12TS oc8051_alu1_u150 ( .A(oc8051_alu1_n48), .B(oc8051_alu1_n62), 
        .Y(oc8051_alu1_n13) );
  NAND2_X0P5A_A12TS oc8051_alu1_u149 ( .A(oc8051_alu1_n135), .B(
        oc8051_alu1_n13), .Y(oc8051_alu1_n133) );
  NOR2_X0P5A_A12TS oc8051_alu1_u148 ( .A(oc8051_alu1_n87), .B(oc8051_alu1_n122), .Y(oc8051_alu1_n134) );
  INV_X0P5B_A12TS oc8051_alu1_u146 ( .A(src2[7]), .Y(oc8051_alu1_n114) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u145 ( .A(oc8051_alu1_n133), .B(
        oc8051_alu1_n134), .S0(oc8051_alu1_n114), .Y(oc8051_alu1_n132) );
  AND3_X0P5M_A12TS oc8051_alu1_u144 ( .A(oc8051_alu1_n203), .B(
        oc8051_alu1_n202), .C(oc8051_alu1_n132), .Y(oc8051_alu1_n94) );
  INV_X0P5B_A12TS oc8051_alu1_u143 ( .A(oc8051_alu1_n131), .Y(oc8051_alu1_n129) );
  NOR2_X0P5A_A12TS oc8051_alu1_u142 ( .A(oc8051_alu1_n131), .B(oc8051_alu1_n19), .Y(oc8051_alu1_n130) );
  INV_X0P5B_A12TS oc8051_alu1_u141 ( .A(src2[6]), .Y(oc8051_alu1_n20) );
  OAI22_X0P5M_A12TS oc8051_alu1_u140 ( .A0(src1[6]), .A1(oc8051_alu1_n129), 
        .B0(oc8051_alu1_n130), .B1(oc8051_alu1_n20), .Y(oc8051_alu1_n28) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u139 ( .A(oc8051_alu1_n28), .B(
        oc8051_alu1_n114), .Y(oc8051_alu1_n128) );
  NAND2_X0P5A_A12TS oc8051_alu1_u138 ( .A(oc8051_alu1_n128), .B(
        oc8051_alu1_n87), .Y(oc8051_alu1_n51) );
  OAI21_X0P5M_A12TS oc8051_alu1_u137 ( .A0(oc8051_alu1_n87), .A1(
        oc8051_alu1_n128), .B0(oc8051_alu1_n51), .Y(sub_result[7]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u136 ( .A0(oc8051_alu1_divsrc1[7]), .A1(
        oc8051_alu1_n222), .B0(oc8051_alu1_n49), .B1(sub_result[7]), .Y(
        oc8051_alu1_n119) );
  AND2_X0P5M_A12TS oc8051_alu1_u135 ( .A(oc8051_alu1_n126), .B(src1[6]), .Y(
        oc8051_alu1_n127) );
  OAI22_X0P5M_A12TS oc8051_alu1_u134 ( .A0(src1[6]), .A1(oc8051_alu1_n126), 
        .B0(src2[6]), .B1(oc8051_alu1_n127), .Y(oc8051_alu1_n26) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u133 ( .A(oc8051_alu1_n26), .B(
        oc8051_alu1_n114), .Y(oc8051_alu1_n115) );
  AO1B2_X0P5M_A12TS oc8051_alu1_u131 ( .B0(oc8051_alu1_n223), .B1(
        oc8051_alu1_n115), .A0N(oc8051_alu1_n125), .Y(oc8051_alu1_n121) );
  NOR2_X0P5A_A12TS oc8051_alu1_u130 ( .A(oc8051_alu1_n115), .B(oc8051_alu1_n23), .Y(oc8051_alu1_n123) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u129 ( .A(oc8051_alu1_n121), .B(
        oc8051_alu1_n123), .S0(oc8051_alu1_n87), .Y(oc8051_alu1_n120) );
  NAND4B_X0P5M_A12TS oc8051_alu1_u128 ( .AN(oc8051_alu1_n118), .B(
        oc8051_alu1_n94), .C(oc8051_alu1_n119), .D(oc8051_alu1_n120), .Y(
        oc8051_alu1_n2200) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u127 ( .AN(oc8051_alu1_n3), .B(
        oc8051_alu1_n117), .Y(oc8051_alu1_u3_u2_z_0) );
  NOR2_X0P5A_A12TS oc8051_alu1_u126 ( .A(alu_cy), .B(oc8051_alu1_u3_u2_z_0), 
        .Y(oc8051_alu1_n116) );
  AO21A1AI2_X0P5M_A12TS oc8051_alu1_u125 ( .A0(oc8051_alu1_n19), .A1(
        oc8051_alu1_n99), .B0(oc8051_alu1_n87), .C0(oc8051_alu1_n116), .Y(
        oc8051_alu1_u3_u1_z_2) );
  OAI22_X0P5M_A12TS oc8051_alu1_u124 ( .A0(oc8051_alu1_n114), .A1(
        oc8051_alu1_n26), .B0(oc8051_alu1_n87), .B1(oc8051_alu1_n115), .Y(
        oc8051_alu1_addc_1_) );
  NAND4_X0P5A_A12TS oc8051_alu1_u123 ( .A(oc8051_alu1_n111), .B(
        oc8051_alu1_n112), .C(oc8051_alu1_n23), .D(oc8051_alu1_n113), .Y(
        oc8051_alu1_n108) );
  NAND4B_X0P5M_A12TS oc8051_alu1_u122 ( .AN(oc8051_alu1_n108), .B(
        oc8051_alu1_n43), .C(oc8051_alu1_n109), .D(oc8051_alu1_n110), .Y(
        oc8051_alu1_n174) );
  AO22_X0P5M_A12TS oc8051_alu1_u121 ( .A0(oc8051_alu1_n240), .A1(
        oc8051_alu1_n107), .B0(oc8051_alu1_n174), .B1(src1[0]), .Y(wr_dat[0])
         );
  AO22_X0P5M_A12TS oc8051_alu1_u120 ( .A0(oc8051_alu1_n240), .A1(
        oc8051_alu1_n106), .B0(oc8051_alu1_n174), .B1(src1[1]), .Y(wr_dat[1])
         );
  AO22_X0P5M_A12TS oc8051_alu1_u119 ( .A0(oc8051_alu1_n240), .A1(
        oc8051_alu1_n105), .B0(oc8051_alu1_n174), .B1(src1[2]), .Y(wr_dat[2])
         );
  INV_X0P5B_A12TS oc8051_alu1_u117 ( .A(oc8051_alu1_n175), .Y(wr_dat[3]) );
  INV_X0P5B_A12TS oc8051_alu1_u116 ( .A(oc8051_alu1_n240), .Y(oc8051_alu1_n32)
         );
  INV_X0P5B_A12TS oc8051_alu1_u115 ( .A(oc8051_alu1_n104), .Y(oc8051_alu1_n101) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u114 ( .A0(oc8051_alu1_n48), .A1(
        oc8051_alu1_sub_1_root_sub_189_2_carry_0_), .B0(oc8051_alu1_n103), 
        .C0(oc8051_alu1_n174), .Y(oc8051_alu1_n95) );
  INV_X0P5B_A12TS oc8051_alu1_u113 ( .A(oc8051_alu1_n100), .Y(oc8051_alu1_n98)
         );
  INV_X0P5B_A12TS oc8051_alu1_u112 ( .A(oc8051_alu1_n97), .Y(oc8051_alu1_n96)
         );
  AOI22_X0P5M_A12TS oc8051_alu1_u111 ( .A0(oc8051_alu1_inc[8]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[8]), .B1(oc8051_alu1_n138), .Y(
        oc8051_alu1_n89) );
  AOI22_X0P5M_A12TS oc8051_alu1_u110 ( .A0(src1[0]), .A1(oc8051_alu1_n79), 
        .B0(oc8051_alu1_n1340), .B1(oc8051_alu1_n223), .Y(oc8051_alu1_n90) );
  AOI22_X0P5M_A12TS oc8051_alu1_u109 ( .A0(oc8051_alu1_mulsrc2[0]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc2[0]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n92) );
  INV_X0P5B_A12TS oc8051_alu1_u108 ( .A(oc8051_alu1_n43), .Y(oc8051_alu1_n56)
         );
  AOI22_X0P5M_A12TS oc8051_alu1_u107 ( .A0(oc8051_alu1_n56), .A1(src2[0]), 
        .B0(oc8051_alu1_n33), .B1(src1[4]), .Y(oc8051_alu1_n93) );
  NAND4_X0P5A_A12TS oc8051_alu1_u106 ( .A(oc8051_alu1_n89), .B(oc8051_alu1_n90), .C(oc8051_alu1_n92), .D(oc8051_alu1_n93), .Y(des2[0]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u105 ( .A0(oc8051_alu1_inc[9]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[9]), .B1(oc8051_alu1_n138), .Y(
        oc8051_alu1_n84) );
  AOI22_X0P5M_A12TS oc8051_alu1_u104 ( .A0(src1[1]), .A1(oc8051_alu1_n79), 
        .B0(oc8051_alu1_n1350), .B1(oc8051_alu1_n223), .Y(oc8051_alu1_n85) );
  AOI22_X0P5M_A12TS oc8051_alu1_u103 ( .A0(oc8051_alu1_mulsrc2[1]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc2[1]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n86) );
  AOI22_X0P5M_A12TS oc8051_alu1_u102 ( .A0(oc8051_alu1_n56), .A1(src2[1]), 
        .B0(oc8051_alu1_n33), .B1(src1[5]), .Y(oc8051_alu1_n88) );
  NAND4_X0P5A_A12TS oc8051_alu1_u99 ( .A(oc8051_alu1_n84), .B(oc8051_alu1_n85), 
        .C(oc8051_alu1_n86), .D(oc8051_alu1_n88), .Y(des2[1]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u98 ( .A0(oc8051_alu1_inc[10]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[10]), .B1(oc8051_alu1_n138), 
        .Y(oc8051_alu1_n80) );
  AOI22_X0P5M_A12TS oc8051_alu1_u97 ( .A0(src1[2]), .A1(oc8051_alu1_n79), .B0(
        oc8051_alu1_n1360), .B1(oc8051_alu1_n223), .Y(oc8051_alu1_n81) );
  AOI22_X0P5M_A12TS oc8051_alu1_u96 ( .A0(oc8051_alu1_mulsrc2[2]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc2[2]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n82) );
  AOI22_X0P5M_A12TS oc8051_alu1_u95 ( .A0(oc8051_alu1_n56), .A1(src2[2]), .B0(
        oc8051_alu1_n33), .B1(src1[6]), .Y(oc8051_alu1_n83) );
  NAND4_X0P5A_A12TS oc8051_alu1_u94 ( .A(oc8051_alu1_n80), .B(oc8051_alu1_n81), 
        .C(oc8051_alu1_n82), .D(oc8051_alu1_n83), .Y(des2[2]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u93 ( .A0(oc8051_alu1_inc[11]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[11]), .B1(oc8051_alu1_n138), 
        .Y(oc8051_alu1_n75) );
  AOI22_X0P5M_A12TS oc8051_alu1_u92 ( .A0(oc8051_alu1_n79), .A1(src1[3]), .B0(
        oc8051_alu1_n1370), .B1(oc8051_alu1_n223), .Y(oc8051_alu1_n76) );
  AOI22_X0P5M_A12TS oc8051_alu1_u91 ( .A0(oc8051_alu1_mulsrc2[3]), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divsrc2[3]), .B1(oc8051_alu1_n222), 
        .Y(oc8051_alu1_n77) );
  AOI22_X0P5M_A12TS oc8051_alu1_u90 ( .A0(oc8051_alu1_n56), .A1(src2[3]), .B0(
        oc8051_alu1_n33), .B1(src1[7]), .Y(oc8051_alu1_n78) );
  NAND4_X0P5A_A12TS oc8051_alu1_u89 ( .A(oc8051_alu1_n75), .B(oc8051_alu1_n76), 
        .C(oc8051_alu1_n77), .D(oc8051_alu1_n78), .Y(des2[3]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u88 ( .A0(oc8051_alu1_inc[12]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[12]), .B1(oc8051_alu1_n138), 
        .Y(oc8051_alu1_n71) );
  AOI22_X0P5M_A12TS oc8051_alu1_u87 ( .A0(oc8051_alu1_divsrc2[4]), .A1(
        oc8051_alu1_n222), .B0(oc8051_alu1_n1380), .B1(oc8051_alu1_n223), .Y(
        oc8051_alu1_n72) );
  AOI22_X0P5M_A12TS oc8051_alu1_u86 ( .A0(oc8051_alu1_n33), .A1(src1[0]), .B0(
        oc8051_alu1_mulsrc2[4]), .B1(oc8051_alu1_n225), .Y(oc8051_alu1_n73) );
  AOI22_X0P5M_A12TS oc8051_alu1_u85 ( .A0(src2[4]), .A1(oc8051_alu1_n61), .B0(
        oc8051_alu1_n62), .B1(src1[4]), .Y(oc8051_alu1_n74) );
  NAND4_X0P5A_A12TS oc8051_alu1_u84 ( .A(oc8051_alu1_n71), .B(oc8051_alu1_n72), 
        .C(oc8051_alu1_n73), .D(oc8051_alu1_n74), .Y(des2[4]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u83 ( .A0(oc8051_alu1_inc[13]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[13]), .B1(oc8051_alu1_n138), 
        .Y(oc8051_alu1_n67) );
  AOI22_X0P5M_A12TS oc8051_alu1_u82 ( .A0(oc8051_alu1_divsrc2[5]), .A1(
        oc8051_alu1_n222), .B0(oc8051_alu1_n1390), .B1(oc8051_alu1_n223), .Y(
        oc8051_alu1_n68) );
  AOI22_X0P5M_A12TS oc8051_alu1_u81 ( .A0(src1[1]), .A1(oc8051_alu1_n33), .B0(
        oc8051_alu1_mulsrc2[5]), .B1(oc8051_alu1_n225), .Y(oc8051_alu1_n69) );
  AOI22_X0P5M_A12TS oc8051_alu1_u80 ( .A0(src2[5]), .A1(oc8051_alu1_n61), .B0(
        oc8051_alu1_n62), .B1(src1[5]), .Y(oc8051_alu1_n70) );
  NAND4_X0P5A_A12TS oc8051_alu1_u79 ( .A(oc8051_alu1_n67), .B(oc8051_alu1_n68), 
        .C(oc8051_alu1_n69), .D(oc8051_alu1_n70), .Y(des2[5]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u77 ( .A0(oc8051_alu1_inc[14]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[14]), .B1(oc8051_alu1_n138), 
        .Y(oc8051_alu1_n63) );
  AOI22_X0P5M_A12TS oc8051_alu1_u76 ( .A0(oc8051_alu1_divsrc2[6]), .A1(
        oc8051_alu1_n222), .B0(oc8051_alu1_n1400), .B1(oc8051_alu1_n223), .Y(
        oc8051_alu1_n64) );
  AOI22_X0P5M_A12TS oc8051_alu1_u75 ( .A0(src1[2]), .A1(oc8051_alu1_n33), .B0(
        oc8051_alu1_mulsrc2[6]), .B1(oc8051_alu1_n225), .Y(oc8051_alu1_n65) );
  AOI22_X0P5M_A12TS oc8051_alu1_u74 ( .A0(src2[6]), .A1(oc8051_alu1_n61), .B0(
        oc8051_alu1_n62), .B1(src1[6]), .Y(oc8051_alu1_n66) );
  NAND4_X0P5A_A12TS oc8051_alu1_u73 ( .A(oc8051_alu1_n63), .B(oc8051_alu1_n64), 
        .C(oc8051_alu1_n65), .D(oc8051_alu1_n66), .Y(des2[6]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u72 ( .A0(oc8051_alu1_inc[15]), .A1(
        oc8051_alu1_n137), .B0(oc8051_alu1_dec[15]), .B1(oc8051_alu1_n138), 
        .Y(oc8051_alu1_n57) );
  AOI22_X0P5M_A12TS oc8051_alu1_u71 ( .A0(oc8051_alu1_divsrc2[7]), .A1(
        oc8051_alu1_n222), .B0(oc8051_alu1_n1410), .B1(oc8051_alu1_n223), .Y(
        oc8051_alu1_n58) );
  AOI22_X0P5M_A12TS oc8051_alu1_u70 ( .A0(oc8051_alu1_n33), .A1(src1[3]), .B0(
        oc8051_alu1_mulsrc2[7]), .B1(oc8051_alu1_n225), .Y(oc8051_alu1_n59) );
  AOI22_X0P5M_A12TS oc8051_alu1_u69 ( .A0(src2[7]), .A1(oc8051_alu1_n61), .B0(
        oc8051_alu1_n62), .B1(src1[7]), .Y(oc8051_alu1_n60) );
  NAND4_X0P5A_A12TS oc8051_alu1_u68 ( .A(oc8051_alu1_n57), .B(oc8051_alu1_n58), 
        .C(oc8051_alu1_n59), .D(oc8051_alu1_n60), .Y(des2[7]) );
  AOI222_X0P5M_A12TS oc8051_alu1_u67 ( .A0(oc8051_alu1_n55), .A1(
        oc8051_alu1_n49), .B0(oc8051_alu1_n56), .B1(srcac), .C0(
        oc8051_alu1_add4_4_), .C1(oc8051_alu1_n223), .Y(oc8051_alu1_n54) );
  INV_X0P5B_A12TS oc8051_alu1_u66 ( .A(oc8051_alu1_n54), .Y(desac) );
  AOI22_X0P5M_A12TS oc8051_alu1_u65 ( .A0(oc8051_alu1_n1810), .A1(
        oc8051_alu1_n52), .B0(src1[0]), .B1(oc8051_alu1_n53), .Y(
        oc8051_alu1_n29) );
  AO1B2_X0P5M_A12TS oc8051_alu1_u64 ( .B0(oc8051_alu1_n28), .B1(src2[7]), 
        .A0N(oc8051_alu1_n51), .Y(oc8051_alu1_n27) );
  AOI22_X0P5M_A12TS oc8051_alu1_u63 ( .A0(oc8051_alu1_n49), .A1(
        oc8051_alu1_n27), .B0(oc8051_alu1_n3), .B1(oc8051_alu1_n50), .Y(
        oc8051_alu1_n30) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u62 ( .A(oc8051_alu1_n47), .B(oc8051_alu1_n48), 
        .S0(bit_out), .Y(oc8051_alu1_n35) );
  NAND2_X0P5A_A12TS oc8051_alu1_u61 ( .A(oc8051_alu1_n122), .B(oc8051_alu1_n46), .Y(oc8051_alu1_n44) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u60 ( .A(oc8051_alu1_n44), .B(oc8051_alu1_n45), 
        .S0(bit_out), .Y(oc8051_alu1_n41) );
  NAND4_X0P5A_A12TS oc8051_alu1_u59 ( .A(oc8051_alu1_n41), .B(oc8051_alu1_n42), 
        .C(oc8051_alu1_n43), .D(oc8051_alu1_n12), .Y(oc8051_alu1_n37) );
  AO1B2_X0P5M_A12TS oc8051_alu1_u58 ( .B0(oc8051_alu1_n39), .B1(bit_out), 
        .A0N(oc8051_alu1_n40), .Y(oc8051_alu1_n38) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u57 ( .A(oc8051_alu1_n37), .B(oc8051_alu1_n38), 
        .S0(oc8051_alu1_sub_1_root_sub_189_2_carry_0_), .Y(oc8051_alu1_n36) );
  NAND2_X0P5A_A12TS oc8051_alu1_u56 ( .A(oc8051_alu1_n35), .B(oc8051_alu1_n36), 
        .Y(oc8051_alu1_n34) );
  AOI221_X0P5M_A12TS oc8051_alu1_u55 ( .A0(oc8051_alu1_n33), .A1(src1[7]), 
        .B0(oc8051_alu1_n223), .B1(oc8051_alu1_addc_1_), .C0(oc8051_alu1_n34), 
        .Y(oc8051_alu1_n31) );
  AOI31_X0P5M_A12TS oc8051_alu1_u54 ( .A0(oc8051_alu1_n29), .A1(
        oc8051_alu1_n30), .A2(oc8051_alu1_n31), .B0(oc8051_alu1_n32), .Y(descy) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u53 ( .A(oc8051_alu1_n27), .B(oc8051_alu1_n28), 
        .Y(oc8051_alu1_n21) );
  XOR2_X0P5M_A12TS oc8051_alu1_u52 ( .A(oc8051_alu1_n26), .B(
        oc8051_alu1_addc_1_), .Y(oc8051_alu1_n24) );
  AOI22_X0P5M_A12TS oc8051_alu1_u51 ( .A0(oc8051_alu1_mulov), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_divov), .B1(oc8051_alu1_n222), .Y(
        oc8051_alu1_n25) );
  OAI221_X0P5M_A12TS oc8051_alu1_u50 ( .A0(oc8051_alu1_n21), .A1(
        oc8051_alu1_n22), .B0(oc8051_alu1_n23), .B1(oc8051_alu1_n24), .C0(
        oc8051_alu1_n25), .Y(desov) );
  AND2_X0P5M_A12TS oc8051_alu1_u49 ( .A(oc8051_alu1_des_acc_1[0]), .B(
        oc8051_alu1_n240), .Y(des_acc[0]) );
  AND2_X0P5M_A12TS oc8051_alu1_u48 ( .A(oc8051_alu1_des_acc_1[1]), .B(
        oc8051_alu1_n240), .Y(des_acc[1]) );
  AND2_X0P5M_A12TS oc8051_alu1_u47 ( .A(oc8051_alu1_des_acc_1[2]), .B(
        oc8051_alu1_n240), .Y(des_acc[2]) );
  AND2_X0P5M_A12TS oc8051_alu1_u46 ( .A(oc8051_alu1_des_acc_1[3]), .B(
        oc8051_alu1_n240), .Y(des_acc[3]) );
  AND2_X0P5M_A12TS oc8051_alu1_u45 ( .A(oc8051_alu1_des_acc_1[4]), .B(
        oc8051_alu1_n240), .Y(des_acc[4]) );
  AND2_X0P5M_A12TS oc8051_alu1_u44 ( .A(oc8051_alu1_des_acc_1[5]), .B(
        oc8051_alu1_n240), .Y(des_acc[5]) );
  AND2_X0P5M_A12TS oc8051_alu1_u43 ( .A(oc8051_alu1_des_acc_1[6]), .B(
        oc8051_alu1_n240), .Y(des_acc[6]) );
  AND2_X0P5M_A12TS oc8051_alu1_u42 ( .A(oc8051_alu1_des_acc_1[7]), .B(
        oc8051_alu1_n240), .Y(des_acc[7]) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u41 ( .A0(oc8051_alu1_n124), .A1(
        oc8051_alu1_n19), .B0(oc8051_alu1_n13), .C0(oc8051_alu1_n20), .Y(
        oc8051_alu1_n218) );
  OAI22_X0P5M_A12TS oc8051_alu1_u40 ( .A0(oc8051_alu1_n13), .A1(
        oc8051_alu1_n17), .B0(oc8051_alu1_n124), .B1(oc8051_alu1_n18), .Y(
        oc8051_alu1_n228) );
  OAI22_X0P5M_A12TS oc8051_alu1_u39 ( .A0(oc8051_alu1_n13), .A1(
        oc8051_alu1_n15), .B0(oc8051_alu1_n124), .B1(oc8051_alu1_n16), .Y(
        oc8051_alu1_n237) );
  OAI21_X0P5M_A12TS oc8051_alu1_u38 ( .A0(src2[3]), .A1(oc8051_alu1_n122), 
        .B0(oc8051_alu1_n12), .Y(oc8051_alu1_n245) );
  INV_X0P5B_A12TS oc8051_alu1_u37 ( .A(src1[3]), .Y(oc8051_alu1_n91) );
  INV_X0P5B_A12TS oc8051_alu1_u36 ( .A(src2[0]), .Y(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[0]) );
  INV_X0P5B_A12TS oc8051_alu1_u35 ( .A(src2[1]), .Y(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[1]) );
  INV_X0P5B_A12TS oc8051_alu1_u34 ( .A(src2[2]), .Y(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[2]) );
  INV_X0P5B_A12TS oc8051_alu1_u33 ( .A(src2[3]), .Y(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[3]) );
  TIEHI_X1M_A12TS oc8051_alu1_u32 ( .Y(oc8051_alu1_n14) );
  NAND2_X1M_A12TS oc8051_alu1_u31 ( .A(src3[6]), .B(oc8051_alu1_n9), .Y(
        oc8051_alu1_n11) );
  XNOR2_X1M_A12TS oc8051_alu1_u30 ( .A(src3[7]), .B(oc8051_alu1_n11), .Y(
        oc8051_alu1_n1410) );
  AND2_X1M_A12TS oc8051_alu1_u29 ( .A(src3[5]), .B(oc8051_alu1_n8), .Y(
        oc8051_alu1_n9) );
  AND2_X1M_A12TS oc8051_alu1_u28 ( .A(src3[4]), .B(oc8051_alu1_n7), .Y(
        oc8051_alu1_n8) );
  AND2_X1M_A12TS oc8051_alu1_u27 ( .A(src3[3]), .B(oc8051_alu1_n6), .Y(
        oc8051_alu1_n7) );
  AND2_X1M_A12TS oc8051_alu1_u26 ( .A(src3[2]), .B(oc8051_alu1_n5), .Y(
        oc8051_alu1_n6) );
  AND2_X1M_A12TS oc8051_alu1_u25 ( .A(src3[1]), .B(oc8051_alu1_n4), .Y(
        oc8051_alu1_n5) );
  AND2_X1M_A12TS oc8051_alu1_u24 ( .A(oc8051_alu1_addc_1_), .B(src3[0]), .Y(
        oc8051_alu1_n4) );
  XOR2_X1M_A12TS oc8051_alu1_u23 ( .A(src3[6]), .B(oc8051_alu1_n9), .Y(
        oc8051_alu1_n1400) );
  XOR2_X1M_A12TS oc8051_alu1_u22 ( .A(src3[5]), .B(oc8051_alu1_n8), .Y(
        oc8051_alu1_n1390) );
  XOR2_X1M_A12TS oc8051_alu1_u21 ( .A(src3[4]), .B(oc8051_alu1_n7), .Y(
        oc8051_alu1_n1380) );
  NAND2_X1M_A12TS oc8051_alu1_u20 ( .A(src1[7]), .B(oc8051_alu1_r450_carry_3_), 
        .Y(oc8051_alu1_n10) );
  XNOR2_X1M_A12TS oc8051_alu1_u19 ( .A(alu_cy), .B(oc8051_alu1_n10), .Y(
        oc8051_alu1_n1810) );
  AND2_X1M_A12TS oc8051_alu1_u18 ( .A(src1[3]), .B(oc8051_alu1_n2), .Y(
        oc8051_alu1_n3) );
  XOR2_X1M_A12TS oc8051_alu1_u17 ( .A(oc8051_alu1_addc_1_), .B(src3[0]), .Y(
        oc8051_alu1_n1340) );
  AND2_X1M_A12TS oc8051_alu1_u16 ( .A(src1[4]), .B(oc8051_alu1_u3_u2_z_0), .Y(
        oc8051_alu1_n1) );
  XOR2_X1M_A12TS oc8051_alu1_u15 ( .A(src1[4]), .B(oc8051_alu1_u3_u2_z_0), .Y(
        oc8051_alu1_n1770) );
  XOR2_X1M_A12TS oc8051_alu1_u14 ( .A(src1[7]), .B(oc8051_alu1_r450_carry_3_), 
        .Y(oc8051_alu1_n1800) );
  XOR2_X1M_A12TS oc8051_alu1_u13 ( .A(src3[1]), .B(oc8051_alu1_n4), .Y(
        oc8051_alu1_n1350) );
  XOR2_X0P5M_A12TS oc8051_alu1_u12 ( .A(src1[3]), .B(oc8051_alu1_n2), .Y(
        oc8051_alu1_n1520) );
  XOR2_X1M_A12TS oc8051_alu1_u11 ( .A(src3[2]), .B(oc8051_alu1_n5), .Y(
        oc8051_alu1_n1360) );
  XOR2_X1M_A12TS oc8051_alu1_u10 ( .A(src3[3]), .B(oc8051_alu1_n6), .Y(
        oc8051_alu1_n1370) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u9 ( .A(src1[2]), .B(src1[1]), .Y(
        oc8051_alu1_n1510) );
  OAI22_X1M_A12TS oc8051_alu1_u8 ( .A0(oc8051_alu1_n32), .A1(oc8051_alu1_n101), 
        .B0(oc8051_alu1_n95), .B1(oc8051_alu1_n102), .Y(wr_dat[4]) );
  NAND2_X1M_A12TS oc8051_alu1_u7 ( .A(oc8051_alu1_malicious1), .B(
        oc8051_alu1_n39), .Y(oc8051_alu1_n240) );
  OR2_X0P7M_A12TS oc8051_alu1_u6 ( .A(src1[1]), .B(src1[2]), .Y(oc8051_alu1_n2) );
  OAI22_X1M_A12TS oc8051_alu1_u5 ( .A0(oc8051_alu1_n32), .A1(oc8051_alu1_n98), 
        .B0(oc8051_alu1_n95), .B1(oc8051_alu1_n99), .Y(wr_dat[5]) );
  OAI22_X1M_A12TS oc8051_alu1_u4 ( .A0(oc8051_alu1_n32), .A1(oc8051_alu1_n96), 
        .B0(oc8051_alu1_n95), .B1(oc8051_alu1_n19), .Y(wr_dat[6]) );
  OAI22_X1M_A12TS oc8051_alu1_u3 ( .A0(oc8051_alu1_n32), .A1(oc8051_alu1_n94), 
        .B0(oc8051_alu1_n87), .B1(oc8051_alu1_n95), .Y(wr_dat[7]) );
  ADDFH_X1M_A12TS oc8051_alu1_sub_1_root_sub_189_2_u2_0 ( .A(src1[0]), .B(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[0]), .CI(
        oc8051_alu1_sub_1_root_sub_189_2_carry_0_), .CO(
        oc8051_alu1_sub_1_root_sub_189_2_carry_1_), .SUM(sub_result[0]) );
  ADDFH_X1M_A12TS oc8051_alu1_add_1_root_add_173_2_u1_0 ( .A(src1[0]), .B(
        src2[0]), .CI(alu_cy), .CO(oc8051_alu1_add_1_root_add_173_2_carry[1]), 
        .SUM(oc8051_alu1_add4_0_) );
  ADDFH_X1M_A12TS oc8051_alu1_sub_1_root_sub_189_2_u2_2 ( .A(src1[2]), .B(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[2]), .CI(
        oc8051_alu1_sub_1_root_sub_189_2_carry_2_), .CO(
        oc8051_alu1_sub_1_root_sub_189_2_carry_3_), .SUM(sub_result[2]) );
  ADDFH_X1M_A12TS oc8051_alu1_add_1_root_add_173_2_u1_2 ( .A(src1[2]), .B(
        src2[2]), .CI(oc8051_alu1_add_1_root_add_173_2_carry[2]), .CO(
        oc8051_alu1_add_1_root_add_173_2_carry[3]), .SUM(oc8051_alu1_add4_2_)
         );
  ADDF_X1M_A12TS oc8051_alu1_add_1_root_add_173_2_u1_3 ( .A(src1[3]), .B(
        src2[3]), .CI(oc8051_alu1_add_1_root_add_173_2_carry[3]), .CO(
        oc8051_alu1_add4_4_), .S(oc8051_alu1_add4_3_) );
  ADDF_X1M_A12TS oc8051_alu1_add_1_root_add_173_2_u1_1 ( .A(src1[1]), .B(
        src2[1]), .CI(oc8051_alu1_add_1_root_add_173_2_carry[1]), .CO(
        oc8051_alu1_add_1_root_add_173_2_carry[2]), .S(oc8051_alu1_add4_1_) );
  ADDF_X1M_A12TS oc8051_alu1_sub_1_root_sub_189_2_u2_3 ( .A(src1[3]), .B(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[3]), .CI(
        oc8051_alu1_sub_1_root_sub_189_2_carry_3_), .CO(oc8051_alu1_sub4_4_), 
        .S(sub_result[3]) );
  ADDF_X1M_A12TS oc8051_alu1_sub_1_root_sub_189_2_u2_1 ( .A(src1[1]), .B(
        oc8051_alu1_sub_1_root_sub_189_2_b_not[1]), .CI(
        oc8051_alu1_sub_1_root_sub_189_2_carry_1_), .CO(
        oc8051_alu1_sub_1_root_sub_189_2_carry_2_), .S(sub_result[1]) );
  ADDF_X1M_A12TS oc8051_alu1_r450_u1_2 ( .A(src1[6]), .B(oc8051_alu1_u3_u1_z_2), .CI(oc8051_alu1_r450_carry_2_), .CO(oc8051_alu1_r450_carry_3_), .S(
        oc8051_alu1_n1790) );
  ADDF_X1M_A12TS oc8051_alu1_r450_u1_1 ( .A(src1[5]), .B(oc8051_alu1_u3_u1_z_2), .CI(oc8051_alu1_n1), .CO(oc8051_alu1_r450_carry_2_), .S(oc8051_alu1_n1780)
         );
  AOI22_X3M_A12TS oc8051_alu1_u162 ( .A0(oc8051_alu1_dec[3]), .A1(
        oc8051_alu1_n138), .B0(oc8051_alu1_n224), .B1(oc8051_alu1_n91), .Y(
        oc8051_alu1_n243) );
  OAI221_X4M_A12TS oc8051_alu1_u160 ( .A0(src1[3]), .A1(oc8051_alu1_n122), 
        .B0(oc8051_alu1_n91), .B1(oc8051_alu1_n124), .C0(oc8051_alu1_n247), 
        .Y(oc8051_alu1_n246) );
  AOI222_X2M_A12TS oc8051_alu1_u159 ( .A0(oc8051_alu1_inc[3]), .A1(
        oc8051_alu1_n137), .B0(src1[3]), .B1(oc8051_alu1_n245), .C0(src2[3]), 
        .C1(oc8051_alu1_n246), .Y(oc8051_alu1_n244) );
  AOI221_X3M_A12TS oc8051_alu1_u147 ( .A0(oc8051_alu1_dec[4]), .A1(
        oc8051_alu1_n138), .B0(oc8051_alu1_inc[4]), .B1(oc8051_alu1_n137), 
        .C0(oc8051_alu1_n237), .Y(oc8051_alu1_n236) );
  AOI221_X3M_A12TS oc8051_alu1_u132 ( .A0(oc8051_alu1_dec[5]), .A1(
        oc8051_alu1_n138), .B0(oc8051_alu1_inc[5]), .B1(oc8051_alu1_n137), 
        .C0(oc8051_alu1_n228), .Y(oc8051_alu1_n227) );
  AOI221_X3M_A12TS oc8051_alu1_u118 ( .A0(oc8051_alu1_dec[6]), .A1(
        oc8051_alu1_n138), .B0(oc8051_alu1_inc[6]), .B1(oc8051_alu1_n137), 
        .C0(oc8051_alu1_n218), .Y(oc8051_alu1_n217) );
  NAND2_X2M_A12TS oc8051_alu1_u101 ( .A(oc8051_alu1_inc[7]), .B(
        oc8051_alu1_n137), .Y(oc8051_alu1_n202) );
  AOI22_X3M_A12TS oc8051_alu1_u100 ( .A0(oc8051_alu1_dec[7]), .A1(
        oc8051_alu1_n138), .B0(oc8051_alu1_n224), .B1(oc8051_alu1_n87), .Y(
        oc8051_alu1_n203) );
  AO21A1AI2_X3M_A12TS oc8051_alu1_u78 ( .A0(oc8051_alu1_n174), .A1(src1[3]), 
        .B0(oc8051_alu1_n176), .C0(oc8051_alu1_n240), .Y(oc8051_alu1_n175) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_0_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2130), .Q(oc8051_alu1_des_acc_1[0]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_1_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2140), .Q(oc8051_alu1_des_acc_1[1]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_2_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2150), .Q(oc8051_alu1_des_acc_1[2]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_3_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2160), .Q(oc8051_alu1_des_acc_1[3]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_4_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2170), .Q(oc8051_alu1_des_acc_1[4]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_5_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2180), .Q(oc8051_alu1_des_acc_1[5]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_6_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2190), .Q(oc8051_alu1_des_acc_1[6]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_7_ ( .G(oc8051_alu1_n240), .D(
        oc8051_alu1_n2200), .Q(oc8051_alu1_des_acc_1[7]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_alu_malicious_u12 ( .AN(oc8051_alu1_n223), .B(
        wb_rst_i), .Y(oc8051_alu1_alu_malicious_n5) );
  INV_X0P5B_A12TS oc8051_alu1_alu_malicious_u11 ( .A(
        oc8051_alu1_alu_malicious_state_0_), .Y(oc8051_alu1_alu_malicious_n2)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_alu_malicious_u10 ( .A(
        oc8051_alu1_alu_malicious_n5), .B(oc8051_alu1_alu_malicious_n2), .Y(
        oc8051_alu1_alu_malicious_n7) );
  INV_X0P5B_A12TS oc8051_alu1_alu_malicious_u9 ( .A(
        oc8051_alu1_alu_malicious_n7), .Y(oc8051_alu1_alu_malicious_n70) );
  NAND2_X0P5A_A12TS oc8051_alu1_alu_malicious_u8 ( .A(
        oc8051_alu1_alu_malicious_n5), .B(oc8051_alu1_alu_malicious_state_0_), 
        .Y(oc8051_alu1_alu_malicious_n6) );
  MXIT2_X0P5M_A12TS oc8051_alu1_alu_malicious_u7 ( .A(
        oc8051_alu1_alu_malicious_n6), .B(oc8051_alu1_alu_malicious_n7), .S0(
        oc8051_alu1_alu_malicious_state_1_), .Y(oc8051_alu1_alu_malicious_n8)
         );
  AOI2XB1_X0P5M_A12TS oc8051_alu1_alu_malicious_u6 ( .A1N(
        oc8051_alu1_alu_malicious_state_1_), .A0(oc8051_alu1_alu_malicious_n5), 
        .B0(oc8051_alu1_alu_malicious_n70), .Y(oc8051_alu1_alu_malicious_n3)
         );
  NAND3_X0P5A_A12TS oc8051_alu1_alu_malicious_u5 ( .A(
        oc8051_alu1_alu_malicious_n5), .B(oc8051_alu1_alu_malicious_state_0_), 
        .C(oc8051_alu1_alu_malicious_state_1_), .Y(
        oc8051_alu1_alu_malicious_n4) );
  MXIT2_X0P5M_A12TS oc8051_alu1_alu_malicious_u4 ( .A(
        oc8051_alu1_alu_malicious_n3), .B(oc8051_alu1_alu_malicious_n4), .S0(
        oc8051_alu1_alu_malicious_n1), .Y(oc8051_alu1_alu_malicious_n9) );
  NOR3_X0P5A_A12TS oc8051_alu1_alu_malicious_u3 ( .A(
        oc8051_alu1_alu_malicious_n2), .B(oc8051_alu1_alu_malicious_state_1_), 
        .C(oc8051_alu1_alu_malicious_n1), .Y(oc8051_alu1_malicious1) );
  DFFQN_X1M_A12TS oc8051_alu1_alu_malicious_state_reg_2_ ( .D(
        oc8051_alu1_alu_malicious_n9), .CK(wb_clk_i), .QN(
        oc8051_alu1_alu_malicious_n1) );
  DFFQ_X1M_A12TS oc8051_alu1_alu_malicious_state_reg_1_ ( .D(
        oc8051_alu1_alu_malicious_n8), .CK(wb_clk_i), .Q(
        oc8051_alu1_alu_malicious_state_1_) );
  DFFQ_X1M_A12TS oc8051_alu1_alu_malicious_state_reg_0_ ( .D(
        oc8051_alu1_alu_malicious_n70), .CK(wb_clk_i), .Q(
        oc8051_alu1_alu_malicious_state_0_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u47 ( .A(
        oc8051_alu1_oc8051_mul1_cycle_0_), .Y(oc8051_alu1_oc8051_mul1_n11) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u46 ( .A(
        oc8051_alu1_oc8051_mul1_cycle_1_), .B(oc8051_alu1_oc8051_mul1_n11), 
        .Y(oc8051_alu1_oc8051_mul1_n9) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u45 ( .A(oc8051_alu1_oc8051_mul1_n9), 
        .Y(oc8051_alu1_oc8051_mul1_n19) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u44 ( .A(
        oc8051_alu1_oc8051_mul1_cycle_0_), .B(oc8051_alu1_oc8051_mul1_cycle_1_), .Y(oc8051_alu1_oc8051_mul1_n7) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u43 ( .A0(src2[2]), .A1(
        oc8051_alu1_oc8051_mul1_n19), .B0(src2[6]), .B1(
        oc8051_alu1_oc8051_mul1_n7), .Y(oc8051_alu1_oc8051_mul1_n20) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u42 ( .A(
        oc8051_alu1_oc8051_mul1_n11), .B(oc8051_alu1_oc8051_mul1_cycle_1_), 
        .Y(oc8051_alu1_oc8051_mul1_n10) );
  AOI32_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u41 ( .A0(
        oc8051_alu1_oc8051_mul1_cycle_0_), .A1(
        oc8051_alu1_oc8051_mul1_cycle_1_), .A2(src2[0]), .B0(src2[4]), .B1(
        oc8051_alu1_oc8051_mul1_n10), .Y(oc8051_alu1_oc8051_mul1_n21) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u40 ( .A(
        oc8051_alu1_oc8051_mul1_n20), .B(oc8051_alu1_oc8051_mul1_n21), .Y(
        oc8051_alu1_oc8051_mul1_n70) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u39 ( .A0(src2[3]), .A1(
        oc8051_alu1_oc8051_mul1_n19), .B0(src2[7]), .B1(
        oc8051_alu1_oc8051_mul1_n7), .Y(oc8051_alu1_oc8051_mul1_n16) );
  AOI32_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u38 ( .A0(
        oc8051_alu1_oc8051_mul1_cycle_0_), .A1(
        oc8051_alu1_oc8051_mul1_cycle_1_), .A2(src2[1]), .B0(src2[5]), .B1(
        oc8051_alu1_oc8051_mul1_n10), .Y(oc8051_alu1_oc8051_mul1_n18) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u37 ( .A(
        oc8051_alu1_oc8051_mul1_n16), .B(oc8051_alu1_oc8051_mul1_n18), .Y(
        oc8051_alu1_oc8051_mul1_n80) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u36 ( .A(oc8051_alu1_mulsrc1[1]), 
        .B(oc8051_alu1_mulsrc1[0]), .Y(oc8051_alu1_oc8051_mul1_n12) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u35 ( .A(oc8051_alu1_mulsrc1[3]), 
        .B(oc8051_alu1_mulsrc1[2]), .Y(oc8051_alu1_oc8051_mul1_n13) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u34 ( .A(oc8051_alu1_mulsrc1[5]), 
        .B(oc8051_alu1_mulsrc1[4]), .Y(oc8051_alu1_oc8051_mul1_n14) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u33 ( .A(oc8051_alu1_mulsrc1[7]), 
        .B(oc8051_alu1_mulsrc1[6]), .Y(oc8051_alu1_oc8051_mul1_n15) );
  NAND4_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u32 ( .A(
        oc8051_alu1_oc8051_mul1_n12), .B(oc8051_alu1_oc8051_mul1_n13), .C(
        oc8051_alu1_oc8051_mul1_n14), .D(oc8051_alu1_oc8051_mul1_n15), .Y(
        oc8051_alu1_mulov) );
  XNOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u31 ( .A(oc8051_alu1_n225), .B(
        oc8051_alu1_oc8051_mul1_n11), .Y(oc8051_alu1_oc8051_mul1_n17) );
  MXIT2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u30 ( .A(
        oc8051_alu1_oc8051_mul1_cycle_1_), .B(oc8051_alu1_oc8051_mul1_n10), 
        .S0(oc8051_alu1_n225), .Y(oc8051_alu1_oc8051_mul1_n8) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u29 ( .A(
        oc8051_alu1_oc8051_mul1_n8), .B(oc8051_alu1_oc8051_mul1_n9), .Y(
        oc8051_alu1_oc8051_mul1_n22) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u28 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[8]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_10_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u27 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[9]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_11_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u26 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[10]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_12_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u25 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[11]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_13_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u24 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[12]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_14_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u23 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[13]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_15_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u22 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[0]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_2_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u21 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[1]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_3_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u20 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[2]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_4_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u19 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[3]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_5_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u18 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[4]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_6_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u17 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[5]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_7_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u16 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[6]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_8_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u15 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul[7]), .B(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_shifted_9_) );
  TIELO_X1M_A12TS oc8051_alu1_oc8051_mul1_u14 ( .Y(oc8051_alu1_oc8051_mul1_n5)
         );
  NAND2_X1M_A12TS oc8051_alu1_oc8051_mul1_u13 ( .A(oc8051_alu1_oc8051_mul1_n4), 
        .B(oc8051_alu1_oc8051_mul1_shifted_14_), .Y(oc8051_alu1_oc8051_mul1_n6) );
  XNOR2_X1M_A12TS oc8051_alu1_oc8051_mul1_u12 ( .A(
        oc8051_alu1_oc8051_mul1_shifted_15_), .B(oc8051_alu1_oc8051_mul1_n6), 
        .Y(oc8051_alu1_mulsrc1[7]) );
  AND2_X1M_A12TS oc8051_alu1_oc8051_mul1_u11 ( .A(oc8051_alu1_oc8051_mul1_n3), 
        .B(oc8051_alu1_oc8051_mul1_shifted_13_), .Y(oc8051_alu1_oc8051_mul1_n4) );
  AND2_X1M_A12TS oc8051_alu1_oc8051_mul1_u10 ( .A(oc8051_alu1_oc8051_mul1_n2), 
        .B(oc8051_alu1_oc8051_mul1_shifted_12_), .Y(oc8051_alu1_oc8051_mul1_n3) );
  AND2_X1M_A12TS oc8051_alu1_oc8051_mul1_u9 ( .A(oc8051_alu1_oc8051_mul1_n1), 
        .B(oc8051_alu1_oc8051_mul1_shifted_11_), .Y(oc8051_alu1_oc8051_mul1_n2) );
  AND2_X1M_A12TS oc8051_alu1_oc8051_mul1_u8 ( .A(
        oc8051_alu1_oc8051_mul1_add_96_carry_10_), .B(
        oc8051_alu1_oc8051_mul1_shifted_10_), .Y(oc8051_alu1_oc8051_mul1_n1)
         );
  XOR2_X1M_A12TS oc8051_alu1_oc8051_mul1_u7 ( .A(
        oc8051_alu1_oc8051_mul1_shifted_14_), .B(oc8051_alu1_oc8051_mul1_n4), 
        .Y(oc8051_alu1_mulsrc1[6]) );
  XOR2_X1M_A12TS oc8051_alu1_oc8051_mul1_u6 ( .A(
        oc8051_alu1_oc8051_mul1_shifted_12_), .B(oc8051_alu1_oc8051_mul1_n2), 
        .Y(oc8051_alu1_mulsrc1[4]) );
  XOR2_X1M_A12TS oc8051_alu1_oc8051_mul1_u5 ( .A(
        oc8051_alu1_oc8051_mul1_shifted_11_), .B(oc8051_alu1_oc8051_mul1_n1), 
        .Y(oc8051_alu1_mulsrc1[3]) );
  XOR2_X1M_A12TS oc8051_alu1_oc8051_mul1_u4 ( .A(
        oc8051_alu1_oc8051_mul1_shifted_13_), .B(oc8051_alu1_oc8051_mul1_n3), 
        .Y(oc8051_alu1_mulsrc1[5]) );
  XOR2_X1M_A12TS oc8051_alu1_oc8051_mul1_u3 ( .A(
        oc8051_alu1_oc8051_mul1_shifted_10_), .B(
        oc8051_alu1_oc8051_mul1_add_96_carry_10_), .Y(oc8051_alu1_mulsrc1[2])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_2 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[2]), .B(
        oc8051_alu1_oc8051_mul1_shifted_2_), .CI(oc8051_alu1_oc8051_mul1_n5), 
        .CO(oc8051_alu1_oc8051_mul1_add_96_carry_3_), .S(
        oc8051_alu1_mulsrc2[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_cycle_reg_1_ ( .D(
        oc8051_alu1_oc8051_mul1_n22), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_cycle_1_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_cycle_reg_0_ ( .D(
        oc8051_alu1_oc8051_mul1_n17), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_cycle_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_13_ ( .D(
        oc8051_alu1_mulsrc1[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[13]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_12_ ( .D(
        oc8051_alu1_mulsrc1[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[12]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_11_ ( .D(
        oc8051_alu1_mulsrc1[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[11]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_10_ ( .D(
        oc8051_alu1_mulsrc1[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[10]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_9_ ( .D(
        oc8051_alu1_mulsrc1[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[9]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_8_ ( .D(
        oc8051_alu1_mulsrc1[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[8]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_7_ ( .D(
        oc8051_alu1_mulsrc2[7]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_6_ ( .D(
        oc8051_alu1_mulsrc2[6]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_5_ ( .D(
        oc8051_alu1_mulsrc2[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_4_ ( .D(
        oc8051_alu1_mulsrc2[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_3_ ( .D(
        oc8051_alu1_mulsrc2[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_2_ ( .D(
        oc8051_alu1_mulsrc2[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_1_ ( .D(
        oc8051_alu1_mulsrc2[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_0_ ( .D(
        oc8051_alu1_mulsrc2[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul[0]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_9 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[9]), .B(
        oc8051_alu1_oc8051_mul1_shifted_9_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_9_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_10_), .S(oc8051_alu1_mulsrc1[1])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_8 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[8]), .B(
        oc8051_alu1_oc8051_mul1_shifted_8_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_8_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_9_), .S(oc8051_alu1_mulsrc1[0])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_7 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[7]), .B(
        oc8051_alu1_oc8051_mul1_shifted_7_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_7_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_8_), .S(oc8051_alu1_mulsrc2[7])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_6 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[6]), .B(
        oc8051_alu1_oc8051_mul1_shifted_6_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_6_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_7_), .S(oc8051_alu1_mulsrc2[6])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_5 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[5]), .B(
        oc8051_alu1_oc8051_mul1_shifted_5_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_5_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_6_), .S(oc8051_alu1_mulsrc2[5])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_4 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[4]), .B(
        oc8051_alu1_oc8051_mul1_shifted_4_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_4_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_5_), .S(oc8051_alu1_mulsrc2[4])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_add_96_u1_3 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1[3]), .B(
        oc8051_alu1_oc8051_mul1_shifted_3_), .CI(
        oc8051_alu1_oc8051_mul1_add_96_carry_3_), .CO(
        oc8051_alu1_oc8051_mul1_add_96_carry_4_), .S(oc8051_alu1_mulsrc2[3])
         );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u47 ( .A(
        oc8051_alu1_oc8051_mul1_n80), .Y(oc8051_alu1_oc8051_mul1_mult_90_n32)
         );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u46 ( .A(
        oc8051_alu1_oc8051_mul1_n70), .Y(oc8051_alu1_oc8051_mul1_mult_90_n33)
         );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u45 ( .A(src1[7]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n24) );
  INV_X0P8M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u44 ( .A(src1[6]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n25) );
  INV_X0P5M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u43 ( .A(src1[5]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n26) );
  INV_X0P6M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u42 ( .A(src1[4]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n27) );
  INV_X0P5M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u41 ( .A(src1[0]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n31) );
  INV_X0P5M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u40 ( .A(src1[1]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n30) );
  INV_X0P5M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u39 ( .A(src1[2]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n29) );
  INV_X0P5M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u38 ( .A(src1[3]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n28) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u25 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n31), .Y(oc8051_alu1_mulsrc2[0]) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u24 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n30), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n23) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u23 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n29), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n22) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u22 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n28), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n21) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u21 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n27), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n20) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u20 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n26), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n19) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u19 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n25), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n18) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u18 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n24), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n17) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u17 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n31), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n16) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u16 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n30), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n15) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u15 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n29), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n14) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u14 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n28), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n13) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u13 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n27), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n12) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u12 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n26), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n11) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u11 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n25), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n10) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u10 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n24), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n9) );
  ADDH_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u9 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n23), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n16), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n8), .S(oc8051_alu1_mulsrc2[1]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u8 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n22), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n15), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n8), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n7), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[2]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u7 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n21), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n14), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n7), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n6), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[3]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u6 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n20), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n13), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n6), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n5), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[4]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u5 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n19), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n12), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n5), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n4), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[5]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u4 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n18), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n11), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n4), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n3), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[6]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u3 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n17), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n10), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n3), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n2), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[7]) );
  ADDH_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u2 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n2), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n9), .CO(
        oc8051_alu1_oc8051_mul1_mul_result1[9]), .S(
        oc8051_alu1_oc8051_mul1_mul_result1[8]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u67 ( .A(src2[0]), .Y(
        oc8051_alu1_oc8051_div1_n7) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u66 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .B(oc8051_alu1_oc8051_div1_cycle_0_), .Y(oc8051_alu1_oc8051_div1_n18) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u65 ( .A(oc8051_alu1_oc8051_div1_n7), .B(oc8051_alu1_oc8051_div1_n18), .Y(oc8051_alu1_oc8051_div1_cmp1_1_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u64 ( .A(src2[1]), .Y(
        oc8051_alu1_oc8051_div1_n8) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u63 ( .A(
        oc8051_alu1_oc8051_div1_n18), .B(oc8051_alu1_oc8051_div1_n8), .Y(
        oc8051_alu1_oc8051_div1_cmp1_2_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u62 ( .A(src2[2]), .Y(
        oc8051_alu1_oc8051_div1_n9) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u61 ( .A(
        oc8051_alu1_oc8051_div1_cycle_0_), .Y(oc8051_alu1_oc8051_div1_n23) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u60 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .B(oc8051_alu1_oc8051_div1_n23), 
        .Y(oc8051_alu1_oc8051_div1_n3) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u59 ( .A0(
        oc8051_alu1_oc8051_div1_n9), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n3), .B1(oc8051_alu1_oc8051_div1_n7), .Y(
        oc8051_alu1_oc8051_div1_cmp1_3_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u58 ( .A(src2[3]), .Y(
        oc8051_alu1_oc8051_div1_n10) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u57 ( .A0(
        oc8051_alu1_oc8051_div1_n10), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n8), .B1(oc8051_alu1_oc8051_div1_n3), .Y(
        oc8051_alu1_oc8051_div1_cmp1_4_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u56 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .Y(oc8051_alu1_oc8051_div1_n24) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u55 ( .A(
        oc8051_alu1_oc8051_div1_cycle_0_), .B(oc8051_alu1_oc8051_div1_n24), 
        .Y(oc8051_alu1_oc8051_div1_n30) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u54 ( .A(src2[4]), .Y(
        oc8051_alu1_oc8051_div1_n11) );
  OAI222_X0P5M_A12TS oc8051_alu1_oc8051_div1_u53 ( .A0(
        oc8051_alu1_oc8051_div1_n9), .A1(oc8051_alu1_oc8051_div1_n3), .B0(
        oc8051_alu1_oc8051_div1_n30), .B1(oc8051_alu1_oc8051_div1_n7), .C0(
        oc8051_alu1_oc8051_div1_n11), .C1(oc8051_alu1_oc8051_div1_n18), .Y(
        oc8051_alu1_oc8051_div1_cmp1_5_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u52 ( .A(src2[5]), .Y(
        oc8051_alu1_oc8051_div1_n12) );
  OAI222_X0P5M_A12TS oc8051_alu1_oc8051_div1_u51 ( .A0(
        oc8051_alu1_oc8051_div1_n10), .A1(oc8051_alu1_oc8051_div1_n3), .B0(
        oc8051_alu1_oc8051_div1_n8), .B1(oc8051_alu1_oc8051_div1_n30), .C0(
        oc8051_alu1_oc8051_div1_n12), .C1(oc8051_alu1_oc8051_div1_n18), .Y(
        oc8051_alu1_oc8051_div1_cmp1_6_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u50 ( .A(src2[6]), .Y(
        oc8051_alu1_oc8051_div1_n13) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u49 ( .A(
        oc8051_alu1_oc8051_div1_n23), .B(oc8051_alu1_oc8051_div1_n24), .Y(
        oc8051_alu1_oc8051_div1_n15) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u48 ( .A(oc8051_alu1_oc8051_div1_n30), .Y(oc8051_alu1_oc8051_div1_n4) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u47 ( .A(oc8051_alu1_oc8051_div1_n3), 
        .Y(oc8051_alu1_oc8051_div1_n28) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u46 ( .A0(
        oc8051_alu1_oc8051_div1_n4), .A1(src2[2]), .B0(src2[4]), .B1(
        oc8051_alu1_oc8051_div1_n28), .Y(oc8051_alu1_oc8051_div1_n29) );
  OAI221_X0P5M_A12TS oc8051_alu1_oc8051_div1_u45 ( .A0(
        oc8051_alu1_oc8051_div1_n13), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n15), .B1(oc8051_alu1_oc8051_div1_n7), .C0(
        oc8051_alu1_oc8051_div1_n29), .Y(oc8051_alu1_oc8051_div1_cmp1_7_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u44 ( .A(src2[7]), .Y(
        oc8051_alu1_oc8051_div1_n14) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u43 ( .A0(
        oc8051_alu1_oc8051_div1_n4), .A1(src2[3]), .B0(
        oc8051_alu1_oc8051_div1_n28), .B1(src2[5]), .Y(
        oc8051_alu1_oc8051_div1_n27) );
  OAI221_X0P5M_A12TS oc8051_alu1_oc8051_div1_u42 ( .A0(
        oc8051_alu1_oc8051_div1_n14), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n15), .B1(oc8051_alu1_oc8051_div1_n8), .C0(
        oc8051_alu1_oc8051_div1_n27), .Y(oc8051_alu1_oc8051_div1_cmp0_7_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u41 ( .A(src1[0]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[0]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_sub1[0]) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u40 ( .A0(src2[5]), .A1(
        oc8051_alu1_oc8051_div1_n23), .B0(src2[3]), .B1(
        oc8051_alu1_oc8051_div1_n24), .Y(oc8051_alu1_oc8051_div1_n19) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u39 ( .A(oc8051_alu1_oc8051_div1_n15), .Y(oc8051_alu1_oc8051_div1_n21) );
  AOI21_X0P5M_A12TS oc8051_alu1_oc8051_div1_u38 ( .A0(
        oc8051_alu1_oc8051_div1_n11), .A1(oc8051_alu1_oc8051_div1_n12), .B0(
        oc8051_alu1_oc8051_div1_cycle_1_), .Y(oc8051_alu1_oc8051_div1_n22) );
  AOI221_X0P5M_A12TS oc8051_alu1_oc8051_div1_u37 ( .A0(
        oc8051_alu1_oc8051_div1_n18), .A1(src2[6]), .B0(
        oc8051_alu1_oc8051_div1_n21), .B1(src2[2]), .C0(
        oc8051_alu1_oc8051_div1_n22), .Y(oc8051_alu1_oc8051_div1_n16) );
  AOI211_X0P5M_A12TS oc8051_alu1_oc8051_div1_u36 ( .A0(src2[1]), .A1(
        oc8051_alu1_oc8051_div1_n21), .B0(oc8051_alu1_oc8051_div1_sub1[8]), 
        .C0(src2[7]), .Y(oc8051_alu1_oc8051_div1_n20) );
  AND3_X0P5M_A12TS oc8051_alu1_oc8051_div1_u35 ( .A(
        oc8051_alu1_oc8051_div1_n19), .B(oc8051_alu1_oc8051_div1_n16), .C(
        oc8051_alu1_oc8051_div1_n20), .Y(oc8051_alu1_divsrc2[1]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u34 ( .A(
        oc8051_alu1_oc8051_div1_sub1[0]), .B(oc8051_alu1_oc8051_div1_sub1[0]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_0_) );
  AOI21_X0P5M_A12TS oc8051_alu1_oc8051_div1_u33 ( .A0(src2[7]), .A1(
        oc8051_alu1_oc8051_div1_n18), .B0(oc8051_alu1_oc8051_div1_sub0[8]), 
        .Y(oc8051_alu1_oc8051_div1_n17) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u32 ( .A(
        oc8051_alu1_oc8051_div1_rem1_0_), .B(oc8051_alu1_oc8051_div1_sub0[0]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[0]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u31 ( .A(src1[1]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[1]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_1_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u30 ( .A(
        oc8051_alu1_oc8051_div1_rem2_1_), .B(oc8051_alu1_oc8051_div1_sub1[1]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_1_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u29 ( .A(
        oc8051_alu1_oc8051_div1_rem1_1_), .B(oc8051_alu1_oc8051_div1_sub0[1]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[1]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u28 ( .A(src1[2]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[2]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_2_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u27 ( .A(
        oc8051_alu1_oc8051_div1_rem2_2_), .B(oc8051_alu1_oc8051_div1_sub1[2]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_2_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u26 ( .A(
        oc8051_alu1_oc8051_div1_rem1_2_), .B(oc8051_alu1_oc8051_div1_sub0[2]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[2]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u25 ( .A(src1[3]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[3]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_3_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u24 ( .A(
        oc8051_alu1_oc8051_div1_rem2_3_), .B(oc8051_alu1_oc8051_div1_sub1[3]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_3_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u23 ( .A(
        oc8051_alu1_oc8051_div1_rem1_3_), .B(oc8051_alu1_oc8051_div1_sub0[3]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[3]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u22 ( .A(src1[4]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[4]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_4_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u21 ( .A(
        oc8051_alu1_oc8051_div1_rem2_4_), .B(oc8051_alu1_oc8051_div1_sub1[4]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_4_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u20 ( .A(
        oc8051_alu1_oc8051_div1_rem1_4_), .B(oc8051_alu1_oc8051_div1_sub0[4]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[4]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u19 ( .A(src1[5]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[5]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_5_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u18 ( .A(
        oc8051_alu1_oc8051_div1_rem2_5_), .B(oc8051_alu1_oc8051_div1_sub1[5]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_5_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u17 ( .A(
        oc8051_alu1_oc8051_div1_rem1_5_), .B(oc8051_alu1_oc8051_div1_sub0[5]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[5]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u16 ( .A(src1[6]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[6]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_6_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u15 ( .A(
        oc8051_alu1_oc8051_div1_rem2_6_), .B(oc8051_alu1_oc8051_div1_sub1[6]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_6_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u14 ( .A(
        oc8051_alu1_oc8051_div1_rem1_6_), .B(oc8051_alu1_oc8051_div1_sub0[6]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[6]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u13 ( .A(src1[7]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[7]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_7_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u12 ( .A(
        oc8051_alu1_oc8051_div1_rem2_7_), .B(oc8051_alu1_oc8051_div1_sub1[7]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_7_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u11 ( .A(
        oc8051_alu1_oc8051_div1_rem1_7_), .B(oc8051_alu1_oc8051_div1_sub0[7]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[7]) );
  NAND4_X0P5A_A12TS oc8051_alu1_oc8051_div1_u10 ( .A(
        oc8051_alu1_oc8051_div1_n11), .B(oc8051_alu1_oc8051_div1_n12), .C(
        oc8051_alu1_oc8051_div1_n13), .D(oc8051_alu1_oc8051_div1_n14), .Y(
        oc8051_alu1_oc8051_div1_n5) );
  NAND4_X0P5A_A12TS oc8051_alu1_oc8051_div1_u9 ( .A(oc8051_alu1_oc8051_div1_n7), .B(oc8051_alu1_oc8051_div1_n8), .C(oc8051_alu1_oc8051_div1_n9), .D(
        oc8051_alu1_oc8051_div1_n10), .Y(oc8051_alu1_oc8051_div1_n6) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u8 ( .A(oc8051_alu1_oc8051_div1_n5), 
        .B(oc8051_alu1_oc8051_div1_n6), .Y(oc8051_alu1_divov) );
  MXIT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u7 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .B(oc8051_alu1_oc8051_div1_n4), 
        .S0(oc8051_alu1_n222), .Y(oc8051_alu1_oc8051_div1_n2) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u6 ( .A(oc8051_alu1_oc8051_div1_n2), .B(oc8051_alu1_oc8051_div1_n3), .Y(oc8051_alu1_oc8051_div1_n25) );
  XOR2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u5 ( .A(oc8051_alu1_n222), .B(
        oc8051_alu1_oc8051_div1_cycle_0_), .Y(oc8051_alu1_oc8051_div1_n26) );
  TIELO_X1M_A12TS oc8051_alu1_oc8051_div1_u4 ( .Y(
        oc8051_alu1_oc8051_div1_cmp1_0_) );
  OA211_X1M_A12TS oc8051_alu1_oc8051_div1_u3 ( .A0(oc8051_alu1_oc8051_div1_n15), .A1(oc8051_alu1_oc8051_div1_n10), .B0(oc8051_alu1_oc8051_div1_n16), .C0(
        oc8051_alu1_oc8051_div1_n17), .Y(oc8051_alu1_divsrc2[0]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_cycle_reg_1_ ( .D(
        oc8051_alu1_oc8051_div1_n25), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_cycle_1_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_cycle_reg_0_ ( .D(
        oc8051_alu1_oc8051_div1_n26), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_cycle_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_3_ ( .D(
        oc8051_alu1_divsrc2[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_2_ ( .D(
        oc8051_alu1_divsrc2[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_1_ ( .D(
        oc8051_alu1_divsrc2[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_0_ ( .D(
        oc8051_alu1_divsrc2[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_5_ ( .D(
        oc8051_alu1_divsrc2[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_4_ ( .D(
        oc8051_alu1_divsrc2[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_2_ ( .D(
        oc8051_alu1_divsrc1[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_3_ ( .D(
        oc8051_alu1_divsrc1[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_4_ ( .D(
        oc8051_alu1_divsrc1[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_5_ ( .D(
        oc8051_alu1_divsrc1[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_6_ ( .D(
        oc8051_alu1_divsrc1[6]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_7_ ( .D(
        oc8051_alu1_divsrc1[7]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_1_ ( .D(
        oc8051_alu1_divsrc1[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_0_ ( .D(
        oc8051_alu1_divsrc1[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[0]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u11 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_1_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_0_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u10 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_2_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_1_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u9 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_3_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_2_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u8 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_4_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_3_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u7 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_5_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_4_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u6 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_6_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_5_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u5 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_7_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_6_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u4 ( .A(
        oc8051_alu1_oc8051_div1_cmp0_7_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_b_not_7_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_98_u3 ( .A(
        oc8051_alu1_oc8051_div1_sub_98_carry[8]), .Y(
        oc8051_alu1_oc8051_div1_sub0[8]) );
  OR2_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2 ( .A(
        oc8051_alu1_oc8051_div1_rem1_0_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_0_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_n1) );
  XNOR2_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u1 ( .A(
        oc8051_alu1_oc8051_div1_sub_98_b_not_0_), .B(
        oc8051_alu1_oc8051_div1_rem1_0_), .Y(oc8051_alu1_oc8051_div1_sub0[0])
         );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_1 ( .A(
        oc8051_alu1_oc8051_div1_rem1_1_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_1_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_n1), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[2]), .S(
        oc8051_alu1_oc8051_div1_sub0[1]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_2 ( .A(
        oc8051_alu1_oc8051_div1_rem1_2_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_2_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_carry[2]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[3]), .S(
        oc8051_alu1_oc8051_div1_sub0[2]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_3 ( .A(
        oc8051_alu1_oc8051_div1_rem1_3_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_3_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_carry[3]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[4]), .S(
        oc8051_alu1_oc8051_div1_sub0[3]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_4 ( .A(
        oc8051_alu1_oc8051_div1_rem1_4_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_4_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_carry[4]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[5]), .S(
        oc8051_alu1_oc8051_div1_sub0[4]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_5 ( .A(
        oc8051_alu1_oc8051_div1_rem1_5_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_5_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_carry[5]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[6]), .S(
        oc8051_alu1_oc8051_div1_sub0[5]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_6 ( .A(
        oc8051_alu1_oc8051_div1_rem1_6_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_6_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_carry[6]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[7]), .S(
        oc8051_alu1_oc8051_div1_sub0[6]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_7 ( .A(
        oc8051_alu1_oc8051_div1_rem1_7_), .B(
        oc8051_alu1_oc8051_div1_sub_98_b_not_7_), .CI(
        oc8051_alu1_oc8051_div1_sub_98_carry[7]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[8]), .S(
        oc8051_alu1_oc8051_div1_sub0[7]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u9 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_1_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[1]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u8 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_2_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[2]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u7 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_3_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[3]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u6 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_4_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[4]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u5 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_5_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[5]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u4 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_6_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[6]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u3 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_7_), .Y(
        oc8051_alu1_oc8051_div1_sub_94_b_not[7]) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_sub_94_u2 ( .A(
        oc8051_alu1_oc8051_div1_sub_94_carry[8]), .Y(
        oc8051_alu1_oc8051_div1_sub1[8]) );
  TIEHI_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u1 ( .Y(
        oc8051_alu1_oc8051_div1_sub_94_n1) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_1 ( .A(
        oc8051_alu1_oc8051_div1_rem2_1_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[1]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_n1), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[2]), .S(
        oc8051_alu1_oc8051_div1_sub1[1]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_2 ( .A(
        oc8051_alu1_oc8051_div1_rem2_2_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[2]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_carry[2]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[3]), .S(
        oc8051_alu1_oc8051_div1_sub1[2]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_3 ( .A(
        oc8051_alu1_oc8051_div1_rem2_3_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[3]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_carry[3]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[4]), .S(
        oc8051_alu1_oc8051_div1_sub1[3]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_4 ( .A(
        oc8051_alu1_oc8051_div1_rem2_4_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[4]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_carry[4]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[5]), .S(
        oc8051_alu1_oc8051_div1_sub1[4]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_5 ( .A(
        oc8051_alu1_oc8051_div1_rem2_5_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[5]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_carry[5]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[6]), .S(
        oc8051_alu1_oc8051_div1_sub1[5]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_6 ( .A(
        oc8051_alu1_oc8051_div1_rem2_6_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[6]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_carry[6]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[7]), .S(
        oc8051_alu1_oc8051_div1_sub1[6]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_7 ( .A(
        oc8051_alu1_oc8051_div1_rem2_7_), .B(
        oc8051_alu1_oc8051_div1_sub_94_b_not[7]), .CI(
        oc8051_alu1_oc8051_div1_sub_94_carry[7]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[8]), .S(
        oc8051_alu1_oc8051_div1_sub1[7]) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u30 ( .A(oc8051_alu1_sub_205_n8), .B(
        src2[3]), .Y(oc8051_alu1_sub_205_n13) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u29 ( .A(src2[3]), .B(
        oc8051_alu1_sub_205_n8), .Y(oc8051_alu1_dec[11]) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u28 ( .A(oc8051_alu1_sub_205_n13), .B(
        src2[4]), .Y(oc8051_alu1_sub_205_n12) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u27 ( .A(oc8051_alu1_sub_205_n12), .B(
        src2[5]), .Y(oc8051_alu1_sub_205_n11) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u26 ( .A(oc8051_alu1_sub_205_n7), .B(
        src2[0]), .Y(oc8051_alu1_sub_205_n10) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u25 ( .A(oc8051_alu1_sub_205_n10), .B(
        src2[1]), .Y(oc8051_alu1_sub_205_n9) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u24 ( .A(oc8051_alu1_sub_205_n9), .B(
        src2[2]), .Y(oc8051_alu1_sub_205_n8) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u23 ( .A(oc8051_alu1_sub_205_n6), .B(
        src1[7]), .Y(oc8051_alu1_sub_205_n7) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u22 ( .A(oc8051_alu1_sub_205_n5), .B(
        src1[6]), .Y(oc8051_alu1_sub_205_n6) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u21 ( .A(oc8051_alu1_sub_205_n4), .B(
        src1[5]), .Y(oc8051_alu1_sub_205_n5) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u20 ( .A(oc8051_alu1_sub_205_n1), .B(
        src1[4]), .Y(oc8051_alu1_sub_205_n4) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u19 ( .A(oc8051_alu1_sub_205_n3), .B(
        src1[3]), .Y(oc8051_alu1_sub_205_n1) );
  NOR2_X1A_A12TS oc8051_alu1_sub_205_u18 ( .A(oc8051_alu1_sub_205_n11), .B(
        src2[6]), .Y(oc8051_alu1_sub_205_n14) );
  XOR2_X1M_A12TS oc8051_alu1_sub_205_u17 ( .A(src2[7]), .B(
        oc8051_alu1_sub_205_n14), .Y(oc8051_alu1_dec[15]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u16 ( .A(src2[6]), .B(
        oc8051_alu1_sub_205_n11), .Y(oc8051_alu1_dec[14]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u15 ( .A(src2[4]), .B(
        oc8051_alu1_sub_205_n13), .Y(oc8051_alu1_dec[12]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u14 ( .A(src2[5]), .B(
        oc8051_alu1_sub_205_n12), .Y(oc8051_alu1_dec[13]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u13 ( .A(src2[0]), .B(
        oc8051_alu1_sub_205_n7), .Y(oc8051_alu1_dec[8]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u12 ( .A(src2[1]), .B(
        oc8051_alu1_sub_205_n10), .Y(oc8051_alu1_dec[9]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u11 ( .A(src2[2]), .B(
        oc8051_alu1_sub_205_n9), .Y(oc8051_alu1_dec[10]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u10 ( .A(src1[7]), .B(
        oc8051_alu1_sub_205_n6), .Y(oc8051_alu1_dec[7]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u9 ( .A(src1[6]), .B(
        oc8051_alu1_sub_205_n5), .Y(oc8051_alu1_dec[6]) );
  XNOR2_X0P7M_A12TS oc8051_alu1_sub_205_u8 ( .A(src1[5]), .B(
        oc8051_alu1_sub_205_n4), .Y(oc8051_alu1_dec[5]) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u7 ( .A(src1[2]), .B(
        oc8051_alu1_sub_205_n2), .Y(oc8051_alu1_dec[2]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u6 ( .A(src1[4]), .B(
        oc8051_alu1_sub_205_n1), .Y(oc8051_alu1_dec[4]) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u5 ( .A(src1[1]), .B(src1[0]), .Y(
        oc8051_alu1_dec[1]) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u4 ( .A(src1[3]), .B(
        oc8051_alu1_sub_205_n3), .Y(oc8051_alu1_dec[3]) );
  OR2_X0P7M_A12TS oc8051_alu1_sub_205_u3 ( .A(oc8051_alu1_sub_205_n2), .B(
        src1[2]), .Y(oc8051_alu1_sub_205_n3) );
  OR2_X0P7M_A12TS oc8051_alu1_sub_205_u2 ( .A(src1[0]), .B(src1[1]), .Y(
        oc8051_alu1_sub_205_n2) );
  INV_X0P5M_A12TS oc8051_alu1_sub_205_u1 ( .A(src1[0]), .Y(oc8051_alu1_dec[0])
         );
  XOR2_X0P5M_A12TS oc8051_alu1_add_204_u2 ( .A(oc8051_alu1_add_204_carry[15]), 
        .B(src2[7]), .Y(oc8051_alu1_inc[15]) );
  INV_X0P5M_A12TS oc8051_alu1_add_204_u1 ( .A(src1[0]), .Y(oc8051_alu1_inc[0])
         );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_3 ( .A(src1[3]), .B(
        oc8051_alu1_add_204_carry[3]), .CO(oc8051_alu1_add_204_carry[4]), .S(
        oc8051_alu1_inc[3]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_2 ( .A(src1[2]), .B(
        oc8051_alu1_add_204_carry[2]), .CO(oc8051_alu1_add_204_carry[3]), .S(
        oc8051_alu1_inc[2]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_1 ( .A(src1[1]), .B(src1[0]), .CO(
        oc8051_alu1_add_204_carry[2]), .S(oc8051_alu1_inc[1]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_4 ( .A(src1[4]), .B(
        oc8051_alu1_add_204_carry[4]), .CO(oc8051_alu1_add_204_carry[5]), .S(
        oc8051_alu1_inc[4]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_5 ( .A(src1[5]), .B(
        oc8051_alu1_add_204_carry[5]), .CO(oc8051_alu1_add_204_carry[6]), .S(
        oc8051_alu1_inc[5]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_6 ( .A(src1[6]), .B(
        oc8051_alu1_add_204_carry[6]), .CO(oc8051_alu1_add_204_carry[7]), .S(
        oc8051_alu1_inc[6]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_7 ( .A(src1[7]), .B(
        oc8051_alu1_add_204_carry[7]), .CO(oc8051_alu1_add_204_carry[8]), .S(
        oc8051_alu1_inc[7]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_10 ( .A(src2[2]), .B(
        oc8051_alu1_add_204_carry[10]), .CO(oc8051_alu1_add_204_carry[11]), 
        .S(oc8051_alu1_inc[10]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_9 ( .A(src2[1]), .B(
        oc8051_alu1_add_204_carry[9]), .CO(oc8051_alu1_add_204_carry[10]), .S(
        oc8051_alu1_inc[9]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_8 ( .A(src2[0]), .B(
        oc8051_alu1_add_204_carry[8]), .CO(oc8051_alu1_add_204_carry[9]), .S(
        oc8051_alu1_inc[8]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_13 ( .A(src2[5]), .B(
        oc8051_alu1_add_204_carry[13]), .CO(oc8051_alu1_add_204_carry[14]), 
        .S(oc8051_alu1_inc[13]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_12 ( .A(src2[4]), .B(
        oc8051_alu1_add_204_carry[12]), .CO(oc8051_alu1_add_204_carry[13]), 
        .S(oc8051_alu1_inc[12]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_14 ( .A(src2[6]), .B(
        oc8051_alu1_add_204_carry[14]), .CO(oc8051_alu1_add_204_carry[15]), 
        .S(oc8051_alu1_inc[14]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_11 ( .A(src2[3]), .B(
        oc8051_alu1_add_204_carry[11]), .CO(oc8051_alu1_add_204_carry[12]), 
        .S(oc8051_alu1_inc[11]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u106 ( .A(oc8051_ram_top1_bit_addr_r), .Y(
        oc8051_ram_top1_n19) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u105 ( .A(oc8051_ram_top1_n19), .B(
        wr_addr[7]), .Y(oc8051_ram_top1_n71) );
  INV_X0P5B_A12TS oc8051_ram_top1_u104 ( .A(bit_addr_o), .Y(
        oc8051_ram_top1_n72) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_u103 ( .A0(rd_addr[1]), .A1(
        oc8051_ram_top1_n72), .B0(oc8051_ram_top1_n70), .B1(rd_addr[4]), .Y(
        oc8051_ram_top1_n58) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_u102 ( .A(oc8051_ram_top1_n3), .B(
        oc8051_ram_top1_n58), .Y(oc8051_ram_top1_n74) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_u101 ( .A0(rd_addr[0]), .A1(
        oc8051_ram_top1_n72), .B0(rd_addr[3]), .B1(oc8051_ram_top1_n70), .Y(
        oc8051_ram_top1_n59) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_u100 ( .A(oc8051_ram_top1_n1), .B(
        oc8051_ram_top1_n59), .Y(oc8051_ram_top1_n75) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u99 ( .A(oc8051_ram_top1_n74), .B(n_0_net_), .C(oc8051_ram_top1_n75), .Y(oc8051_ram_top1_n60) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_u98 ( .A0(wr_addr[2]), .A1(
        oc8051_ram_top1_n19), .B0(wr_addr[5]), .B1(oc8051_ram_top1_n71), .Y(
        oc8051_ram_top1_n73) );
  INV_X0P5B_A12TS oc8051_ram_top1_u97 ( .A(oc8051_ram_top1_n73), .Y(
        oc8051_ram_top1_wr_addr_m_2_) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_u96 ( .A0(rd_addr[2]), .A1(
        oc8051_ram_top1_n72), .B0(rd_addr[5]), .B1(oc8051_ram_top1_n70), .Y(
        oc8051_ram_top1_n57) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_u95 ( .A(oc8051_ram_top1_wr_addr_m_2_), .B(
        oc8051_ram_top1_n57), .Y(oc8051_ram_top1_n61) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u94 ( .A(rd_addr[7]), .B(wr_addr[7]), .Y(
        oc8051_ram_top1_n62) );
  INV_X0P5B_A12TS oc8051_ram_top1_u93 ( .A(oc8051_ram_top1_n71), .Y(
        oc8051_ram_top1_n69) );
  AND2_X0P5M_A12TS oc8051_ram_top1_u92 ( .A(wr_addr[6]), .B(
        oc8051_ram_top1_n69), .Y(oc8051_ram_top1_wr_addr_m_6_) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_u91 ( .AN(rd_addr[6]), .B(
        oc8051_ram_top1_n70), .Y(oc8051_ram_top1_rd_addr_m_6_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u90 ( .A(oc8051_ram_top1_wr_addr_m_6_), 
        .B(oc8051_ram_top1_rd_addr_m_6_), .Y(oc8051_ram_top1_n64) );
  OR2_X0P5M_A12TS oc8051_ram_top1_u89 ( .A(wr_addr[5]), .B(oc8051_ram_top1_n71), .Y(oc8051_ram_top1_wr_addr_m_5_) );
  INV_X0P5B_A12TS oc8051_ram_top1_u88 ( .A(oc8051_ram_top1_n70), .Y(
        oc8051_ram_top1_n68) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u87 ( .A(oc8051_ram_top1_wr_addr_m_5_), 
        .B(oc8051_ram_top1_rd_addr_m_5_), .Y(oc8051_ram_top1_n65) );
  AND2_X0P5M_A12TS oc8051_ram_top1_u86 ( .A(wr_addr[4]), .B(
        oc8051_ram_top1_n69), .Y(oc8051_ram_top1_wr_addr_m_4_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u85 ( .A(oc8051_ram_top1_wr_addr_m_4_), 
        .B(oc8051_ram_top1_rd_addr_m_4_), .Y(oc8051_ram_top1_n66) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u84 ( .A(wr_addr[6]), .B(wr_addr[3]), .S0(
        oc8051_ram_top1_n69), .Y(oc8051_ram_top1_wr_addr_m_3_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u83 ( .A(oc8051_ram_top1_wr_addr_m_3_), 
        .B(oc8051_ram_top1_n2), .Y(oc8051_ram_top1_n67) );
  AND4_X0P5M_A12TS oc8051_ram_top1_u82 ( .A(oc8051_ram_top1_n64), .B(
        oc8051_ram_top1_n65), .C(oc8051_ram_top1_n66), .D(oc8051_ram_top1_n67), 
        .Y(oc8051_ram_top1_n63) );
  NAND4B_X0P5M_A12TS oc8051_ram_top1_u81 ( .AN(oc8051_ram_top1_n60), .B(
        oc8051_ram_top1_n61), .C(oc8051_ram_top1_n62), .D(oc8051_ram_top1_n63), 
        .Y(oc8051_ram_top1_n53) );
  INV_X0P5B_A12TS oc8051_ram_top1_u80 ( .A(oc8051_ram_top1_n53), .Y(
        oc8051_ram_top1_n8) );
  INV_X0P5B_A12TS oc8051_ram_top1_u79 ( .A(oc8051_ram_top1_n59), .Y(
        oc8051_ram_top1_rd_addr_m_0_) );
  INV_X0P5B_A12TS oc8051_ram_top1_u78 ( .A(oc8051_ram_top1_n58), .Y(
        oc8051_ram_top1_rd_addr_m_1_) );
  INV_X0P5B_A12TS oc8051_ram_top1_u77 ( .A(oc8051_ram_top1_n57), .Y(
        oc8051_ram_top1_rd_addr_m_2_) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u76 ( .A(oc8051_ram_top1_rd_data_m[0]), .B(
        oc8051_ram_top1_wr_data_r[0]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[0]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u75 ( .A(oc8051_ram_top1_rd_data_m[1]), .B(
        oc8051_ram_top1_wr_data_r[1]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[1]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u74 ( .A(oc8051_ram_top1_rd_data_m[2]), .B(
        oc8051_ram_top1_wr_data_r[2]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[2]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u73 ( .A(oc8051_ram_top1_rd_data_m[3]), .B(
        oc8051_ram_top1_wr_data_r[3]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[3]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u72 ( .A(oc8051_ram_top1_rd_data_m[4]), .B(
        oc8051_ram_top1_wr_data_r[4]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[4]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u71 ( .A(oc8051_ram_top1_rd_data_m[5]), .B(
        oc8051_ram_top1_wr_data_r[5]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[5]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u70 ( .A(oc8051_ram_top1_rd_data_m[6]), .B(
        oc8051_ram_top1_wr_data_r[6]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[6]) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u69 ( .A(oc8051_ram_top1_rd_data_m[7]), .B(
        oc8051_ram_top1_wr_data_r[7]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        ram_data[7]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u68 ( .A(descy), .Y(oc8051_ram_top1_n16) );
  INV_X0P5B_A12TS oc8051_ram_top1_u67 ( .A(oc8051_ram_top1_n260), .Y(
        oc8051_ram_top1_n54) );
  INV_X0P5B_A12TS oc8051_ram_top1_u66 ( .A(oc8051_ram_top1_n270), .Y(
        oc8051_ram_top1_n55) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u65 ( .A(oc8051_ram_top1_n19), .B(
        oc8051_ram_top1_n280), .Y(oc8051_ram_top1_n56) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u64 ( .A(oc8051_ram_top1_n54), .B(
        oc8051_ram_top1_n55), .C(oc8051_ram_top1_n56), .Y(oc8051_ram_top1_n46)
         );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u63 ( .A(oc8051_ram_top1_n270), .B(
        oc8051_ram_top1_n260), .C(oc8051_ram_top1_n56), .Y(oc8051_ram_top1_n38) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u62 ( .A(oc8051_ram_top1_n260), .B(
        oc8051_ram_top1_n55), .C(oc8051_ram_top1_n56), .Y(oc8051_ram_top1_n31)
         );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u61 ( .A(oc8051_ram_top1_n270), .B(
        oc8051_ram_top1_n54), .C(oc8051_ram_top1_n56), .Y(oc8051_ram_top1_n42)
         );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u60 ( .A(oc8051_ram_top1_n38), .B(
        oc8051_ram_top1_n31), .C(oc8051_ram_top1_n42), .Y(oc8051_ram_top1_n51)
         );
  AND2_X0P5M_A12TS oc8051_ram_top1_u59 ( .A(oc8051_ram_top1_n280), .B(
        oc8051_ram_top1_bit_addr_r), .Y(oc8051_ram_top1_n52) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u58 ( .A(oc8051_ram_top1_n54), .B(
        oc8051_ram_top1_n55), .C(oc8051_ram_top1_n52), .Y(oc8051_ram_top1_n32)
         );
  INV_X0P5B_A12TS oc8051_ram_top1_u57 ( .A(oc8051_ram_top1_n32), .Y(
        oc8051_ram_top1_n41) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u56 ( .A(oc8051_ram_top1_n52), .B(
        oc8051_ram_top1_n55), .C(oc8051_ram_top1_n260), .Y(oc8051_ram_top1_n27) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u55 ( .A(oc8051_ram_top1_n260), .B(
        oc8051_ram_top1_n52), .C(oc8051_ram_top1_n270), .Y(oc8051_ram_top1_n15) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u54 ( .A(oc8051_ram_top1_n52), .B(
        oc8051_ram_top1_n54), .C(oc8051_ram_top1_n270), .Y(oc8051_ram_top1_n23) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u53 ( .A(oc8051_ram_top1_n27), .B(
        oc8051_ram_top1_n15), .C(oc8051_ram_top1_n23), .Y(oc8051_ram_top1_n45)
         );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u52 ( .A0(oc8051_ram_top1_n51), .A1(
        oc8051_ram_top1_n41), .A2(oc8051_ram_top1_n45), .B0(ram_data[0]), .Y(
        oc8051_ram_top1_n49) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u51 ( .A(wr_dat[0]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n50) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u50 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n46), .B0(oc8051_ram_top1_n49), .C0(
        oc8051_ram_top1_n50), .Y(oc8051_ram_top1_wr_data_m[0]) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_u49 ( .A(oc8051_ram_top1_n32), .B(
        oc8051_ram_top1_n42), .C(oc8051_ram_top1_n38), .D(oc8051_ram_top1_n46), 
        .Y(oc8051_ram_top1_n30) );
  OAI21_X0P5M_A12TS oc8051_ram_top1_u48 ( .A0(oc8051_ram_top1_n30), .A1(
        oc8051_ram_top1_n45), .B0(ram_data[1]), .Y(oc8051_ram_top1_n47) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u47 ( .A(wr_dat[1]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n48) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u46 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n31), .B0(oc8051_ram_top1_n47), .C0(
        oc8051_ram_top1_n48), .Y(oc8051_ram_top1_wr_data_m[1]) );
  NAND3B_X0P5M_A12TS oc8051_ram_top1_u45 ( .AN(oc8051_ram_top1_n45), .B(
        oc8051_ram_top1_n46), .C(oc8051_ram_top1_n31), .Y(oc8051_ram_top1_n35)
         );
  INV_X0P5B_A12TS oc8051_ram_top1_u44 ( .A(oc8051_ram_top1_n38), .Y(
        oc8051_ram_top1_n36) );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u43 ( .A0(oc8051_ram_top1_n35), .A1(
        oc8051_ram_top1_n36), .A2(oc8051_ram_top1_n41), .B0(ram_data[2]), .Y(
        oc8051_ram_top1_n43) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u42 ( .A(wr_dat[2]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n44) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u41 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n42), .B0(oc8051_ram_top1_n43), .C0(
        oc8051_ram_top1_n44), .Y(oc8051_ram_top1_wr_data_m[2]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u40 ( .A(oc8051_ram_top1_n42), .Y(
        oc8051_ram_top1_n37) );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u39 ( .A0(oc8051_ram_top1_n35), .A1(
        oc8051_ram_top1_n37), .A2(oc8051_ram_top1_n41), .B0(ram_data[3]), .Y(
        oc8051_ram_top1_n39) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u38 ( .A(wr_dat[3]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n40) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u37 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n38), .B0(oc8051_ram_top1_n39), .C0(
        oc8051_ram_top1_n40), .Y(oc8051_ram_top1_wr_data_m[3]) );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u36 ( .A0(oc8051_ram_top1_n35), .A1(
        oc8051_ram_top1_n36), .A2(oc8051_ram_top1_n37), .B0(ram_data[4]), .Y(
        oc8051_ram_top1_n33) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u35 ( .A(wr_dat[4]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n34) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u34 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n32), .B0(oc8051_ram_top1_n33), .C0(
        oc8051_ram_top1_n34), .Y(oc8051_ram_top1_wr_data_m[4]) );
  NAND2B_X0P5M_A12TS oc8051_ram_top1_u33 ( .AN(oc8051_ram_top1_n30), .B(
        oc8051_ram_top1_n31), .Y(oc8051_ram_top1_n20) );
  INV_X0P5B_A12TS oc8051_ram_top1_u32 ( .A(oc8051_ram_top1_n15), .Y(
        oc8051_ram_top1_n26) );
  INV_X0P5B_A12TS oc8051_ram_top1_u31 ( .A(oc8051_ram_top1_n23), .Y(
        oc8051_ram_top1_n22) );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u30 ( .A0(oc8051_ram_top1_n20), .A1(
        oc8051_ram_top1_n26), .A2(oc8051_ram_top1_n22), .B0(ram_data[5]), .Y(
        oc8051_ram_top1_n28) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u29 ( .A(wr_dat[5]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n29) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u28 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n27), .B0(oc8051_ram_top1_n28), .C0(
        oc8051_ram_top1_n29), .Y(oc8051_ram_top1_wr_data_m[5]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u27 ( .A(oc8051_ram_top1_n27), .Y(
        oc8051_ram_top1_n21) );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u26 ( .A0(oc8051_ram_top1_n20), .A1(
        oc8051_ram_top1_n26), .A2(oc8051_ram_top1_n21), .B0(ram_data[6]), .Y(
        oc8051_ram_top1_n24) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u25 ( .A(wr_dat[6]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n25) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u24 ( .A0(oc8051_ram_top1_n16), .A1(
        oc8051_ram_top1_n23), .B0(oc8051_ram_top1_n24), .C0(
        oc8051_ram_top1_n25), .Y(oc8051_ram_top1_wr_data_m[6]) );
  OAI31_X0P5M_A12TS oc8051_ram_top1_u23 ( .A0(oc8051_ram_top1_n20), .A1(
        oc8051_ram_top1_n21), .A2(oc8051_ram_top1_n22), .B0(ram_data[7]), .Y(
        oc8051_ram_top1_n17) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u22 ( .A(wr_dat[7]), .B(
        oc8051_ram_top1_n19), .Y(oc8051_ram_top1_n18) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u21 ( .A0(oc8051_ram_top1_n15), .A1(
        oc8051_ram_top1_n16), .B0(oc8051_ram_top1_n17), .C0(
        oc8051_ram_top1_n18), .Y(oc8051_ram_top1_wr_data_m[7]) );
  TIEHI_X1M_A12TS oc8051_ram_top1_u20 ( .Y(oc8051_ram_top1__logic1_) );
  MXT4_X1M_A12TS oc8051_ram_top1_u19 ( .A(ram_data[4]), .B(ram_data[6]), .C(
        ram_data[5]), .D(ram_data[7]), .S0(oc8051_ram_top1_n270), .S1(
        oc8051_ram_top1_n260), .Y(oc8051_ram_top1_n5) );
  MXT4_X1M_A12TS oc8051_ram_top1_u18 ( .A(ram_data[0]), .B(ram_data[2]), .C(
        ram_data[1]), .D(ram_data[3]), .S0(oc8051_ram_top1_n270), .S1(
        oc8051_ram_top1_n260), .Y(oc8051_ram_top1_n4) );
  MXT2_X1M_A12TS oc8051_ram_top1_u17 ( .A(oc8051_ram_top1_n4), .B(
        oc8051_ram_top1_n5), .S0(oc8051_ram_top1_n280), .Y(bit_data) );
  BUFH_X1M_A12TS oc8051_ram_top1_u16 ( .A(oc8051_ram_top1_wr_data_m[0]), .Y(
        oc8051_ram_top1_n6) );
  BUFH_X1M_A12TS oc8051_ram_top1_u15 ( .A(oc8051_ram_top1_wr_data_m[1]), .Y(
        oc8051_ram_top1_n7) );
  BUFH_X1M_A12TS oc8051_ram_top1_u14 ( .A(oc8051_ram_top1_wr_data_m[2]), .Y(
        oc8051_ram_top1_n9) );
  BUFH_X1M_A12TS oc8051_ram_top1_u13 ( .A(oc8051_ram_top1_wr_data_m[3]), .Y(
        oc8051_ram_top1_n10) );
  BUFH_X1M_A12TS oc8051_ram_top1_u12 ( .A(oc8051_ram_top1_wr_data_m[6]), .Y(
        oc8051_ram_top1_n13) );
  BUFH_X1M_A12TS oc8051_ram_top1_u11 ( .A(oc8051_ram_top1_wr_data_m[5]), .Y(
        oc8051_ram_top1_n12) );
  BUFH_X1M_A12TS oc8051_ram_top1_u10 ( .A(oc8051_ram_top1_wr_data_m[4]), .Y(
        oc8051_ram_top1_n11) );
  BUFH_X1M_A12TS oc8051_ram_top1_u9 ( .A(oc8051_ram_top1_wr_data_m[7]), .Y(
        oc8051_ram_top1_n14) );
  NAND2B_X2M_A12TS oc8051_ram_top1_u8 ( .AN(rd_addr[5]), .B(
        oc8051_ram_top1_n68), .Y(oc8051_ram_top1_rd_addr_m_5_) );
  NOR2_X0P5M_A12TS oc8051_ram_top1_u7 ( .A(oc8051_ram_top1_n72), .B(rd_addr[7]), .Y(oc8051_ram_top1_n70) );
  NOR2B_X1M_A12TS oc8051_ram_top1_u6 ( .AN(rd_addr[4]), .B(oc8051_ram_top1_n70), .Y(oc8051_ram_top1_rd_addr_m_4_) );
  AO22_X1M_A12TS oc8051_ram_top1_u5 ( .A0(wr_addr[1]), .A1(oc8051_ram_top1_n19), .B0(oc8051_ram_top1_n71), .B1(wr_addr[4]), .Y(oc8051_ram_top1_n3) );
  MXT2_X1M_A12TS oc8051_ram_top1_u4 ( .A(rd_addr[6]), .B(rd_addr[3]), .S0(
        oc8051_ram_top1_n68), .Y(oc8051_ram_top1_n2) );
  AO22_X1M_A12TS oc8051_ram_top1_u3 ( .A0(wr_addr[0]), .A1(oc8051_ram_top1_n19), .B0(wr_addr[3]), .B1(oc8051_ram_top1_n71), .Y(oc8051_ram_top1_n1) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_rd_en_r_reg ( .D(oc8051_ram_top1_n8), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_rd_en_r) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_select_reg_1_ ( .D(rd_addr[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_n270) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_select_reg_0_ ( .D(rd_addr[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_n260) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_select_reg_2_ ( .D(rd_addr[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_n280) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_addr_r_reg ( .D(bit_addr_o), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_bit_addr_r) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_7_ ( .D(oc8051_ram_top1_n14), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_6_ ( .D(oc8051_ram_top1_n13), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_5_ ( .D(oc8051_ram_top1_n12), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_4_ ( .D(oc8051_ram_top1_n11), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_3_ ( .D(oc8051_ram_top1_n10), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_2_ ( .D(oc8051_ram_top1_n9), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_1_ ( .D(oc8051_ram_top1_n7), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_0_ ( .D(oc8051_ram_top1_n6), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[0]) );
  TIEHI_X1M_A12TS oc8051_ram_top1_oc8051_idata_u2 ( .Y(
        oc8051_ram_top1_oc8051_idata__logic1_) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3443 ( .A(
        n_0_net_), .B(oc8051_ram_top1__logic1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3324) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3442 ( .A(
        wr_addr[7]), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3416) );
  AND3_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3441 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3324), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3416), .C(
        oc8051_ram_top1_wr_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3183) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3440 ( .A(
        oc8051_ram_top1_wr_addr_m_5_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3417) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3439 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3417), .B(
        oc8051_ram_top1_wr_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3164) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3438 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3183), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3164), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3437 ( .A(
        oc8051_ram_top1_wr_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3428) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3436 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3428), .B(
        oc8051_ram_top1_wr_addr_m_3_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3430) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3435 ( .A(
        oc8051_ram_top1_n1), .B(oc8051_ram_top1_n3), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3415) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3434 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3430), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3415), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3433 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3432 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1000) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3431 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1001) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3430 ( .A(
        oc8051_ram_top1_n1), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3432) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3429 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3432), .B(oc8051_ram_top1_n3), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3413) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3428 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3413), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3430), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3427 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3426 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1002) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3425 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1003) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3424 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1004) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3423 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1005) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3422 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1006) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3421 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1007) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3420 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1008) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3419 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3434), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1009) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3418 ( .A(
        oc8051_ram_top1_n3), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3431) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3417 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3431), .B(oc8051_ram_top1_n1), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3411) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3416 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3411), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3430), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3415 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3414 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1010) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3413 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1011) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3412 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1012) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3411 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1013) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3410 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1014) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3409 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1015) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3408 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1016) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3407 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3433), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1017) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3406 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3431), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3432), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3409) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3405 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3409), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3430), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3404 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3403 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1018) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3402 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1019) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3401 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1020) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3400 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1021) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3399 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1022) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3398 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1023) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3397 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1024) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3396 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3429), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1025) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3395 ( .A(
        oc8051_ram_top1_wr_addr_m_3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3428), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3424) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3394 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3424), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3415), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3393 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3392 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1026) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3391 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1027) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3390 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1028) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3389 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1029) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3388 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1030) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3387 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1031) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3386 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1032) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3385 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3427), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1033) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3384 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3424), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3413), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3383 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3382 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1034) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3381 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1035) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3380 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1036) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3379 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1037) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3378 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1038) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3377 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1039) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3376 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1040) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3375 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3426), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1041) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3374 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3424), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3411), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3373 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3372 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1042) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3371 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1043) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3370 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1044) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3369 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1045) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3368 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1046) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3367 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1047) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3366 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1048) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3365 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3425), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1049) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3364 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3424), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3409), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3363 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3362 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1050) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3361 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1051) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3360 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1052) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3359 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1053) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3358 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1054) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3357 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1055) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3356 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1056) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3355 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3423), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1057) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3354 ( .A(
        oc8051_ram_top1_wr_addr_m_3_), .B(oc8051_ram_top1_wr_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3419) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3353 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3419), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3415), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3352 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3351 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1058) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3350 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1059) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3349 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1060) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3348 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1061) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3347 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1062) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3346 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1063) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3345 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1064) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3344 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3422), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1065) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3343 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3419), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3413), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3342 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3341 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1066) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3340 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1067) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3339 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1068) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3338 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1069) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3337 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1070) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3336 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1071) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3335 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1072) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3334 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3421), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1073) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3333 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3419), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3411), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3332 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3331 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1074) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3330 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1075) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3329 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1076) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3328 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1077) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3327 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1078) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3326 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1079) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3325 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1080) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3324 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3420), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1081) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3323 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3419), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3409), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3322 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3321 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1082) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3320 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1083) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3319 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1084) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3318 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1085) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3317 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1086) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3316 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1087) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3315 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1088) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3314 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3418), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1089) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3313 ( .A(
        oc8051_ram_top1_wr_addr_m_6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3417), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3255) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3312 ( .A(
        oc8051_ram_top1_wr_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3342) );
  AND3_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3311 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3342), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3416), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3324), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3163) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3310 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3255), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3163), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3309 ( .A(
        oc8051_ram_top1_wr_addr_m_2_), .B(oc8051_ram_top1_wr_addr_m_3_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3408) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3308 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3408), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3415), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3307 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3306 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1090) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3305 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1091) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3304 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1092) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3303 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1093) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3302 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1094) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3301 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1095) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3300 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1096) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3299 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3414), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1097) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3298 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3413), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3408), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3297 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3296 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1098) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3295 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1099) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3294 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1100) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3293 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1101) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3292 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1102) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3291 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1103) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3290 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1104) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3289 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3412), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1105) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3288 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3411), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3408), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3287 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3286 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1106) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3285 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1107) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3284 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1108) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3283 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1109) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3282 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1110) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3281 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1111) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3280 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1112) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3279 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3410), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1113) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3278 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3408), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3409), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3277 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3276 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1114) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3275 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1115) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3274 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1116) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3273 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1117) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3272 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1118) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3271 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1119) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3270 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1120) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3269 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3407), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1121) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3268 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3267 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1122) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3266 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1123) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3265 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1124) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3264 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1125) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3263 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1126) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3262 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1127) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3261 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1128) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3260 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3406), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1129) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3259 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3258 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1130) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3257 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1131) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3256 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1132) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3255 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1133) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3254 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1134) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3253 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1135) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3252 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1136) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3251 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3405), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1137) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3250 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3249 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1138) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3248 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1139) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3247 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1140) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3246 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1141) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3245 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1142) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3244 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1143) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3243 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1144) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3242 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3404), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1145) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3241 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3240 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1146) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3239 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1147) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3238 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1148) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3237 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1149) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3236 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1150) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3235 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1151) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3234 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1152) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3233 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3403), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1153) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3232 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3231 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1154) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3230 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1155) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3229 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1156) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3228 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1157) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3227 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1158) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3226 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1159) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3225 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1160) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3224 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3402), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1161) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3223 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3222 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1162) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3221 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1163) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3220 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1164) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3219 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1165) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3218 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1166) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3217 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1167) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3216 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1168) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3215 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3401), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1169) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3214 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3213 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1170) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3212 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1171) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3211 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1172) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3210 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1173) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3209 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1174) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3208 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1175) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3207 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1176) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3206 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3400), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1177) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3205 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3204 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1178) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3203 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1179) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3202 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1180) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3201 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1181) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3200 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1182) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3199 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1183) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3198 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1184) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3197 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3399), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1185) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3196 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3195 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1186) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3194 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1187) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3193 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1188) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3192 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1189) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3191 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1190) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3190 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1191) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3189 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1192) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3188 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3398), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1193) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3187 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3186 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1194) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3185 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1195) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3184 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1196) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3183 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1197) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3182 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1198) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3181 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1199) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3180 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1200) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3179 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3397), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1201) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3178 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3177 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1202) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3176 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1203) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3175 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1204) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3174 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1205) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3173 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1206) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3172 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1207) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3171 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1208) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3170 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3396), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1209) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3169 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3395), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3168 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1210) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3167 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1211) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3166 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1212) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3165 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1213) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3164 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1214) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3163 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1215) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3162 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1216) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3161 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3394), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1217) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3160 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3255), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3183), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3159 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3158 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1218) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3157 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1219) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3156 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1220) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3155 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1221) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3154 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1222) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3153 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1223) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3152 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1224) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3151 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3393), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1225) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3150 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3149 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1226) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3148 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1227) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3147 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1228) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3146 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1229) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3145 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1230) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3144 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1231) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3143 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1232) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3142 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3392), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1233) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3141 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3140 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1234) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3139 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1235) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3138 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1236) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3137 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1237) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3136 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1238) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3135 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1239) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3134 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1240) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3133 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3391), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1241) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3132 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3131 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1242) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3130 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1243) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3129 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1244) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3128 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1245) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3127 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1246) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3126 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1247) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3125 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1248) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3124 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3390), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1249) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3123 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3122 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1250) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3121 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1251) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3120 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1252) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3119 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1253) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3118 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1254) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3117 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1255) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3116 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1256) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3115 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3389), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1257) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3114 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3113 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1258) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3112 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1259) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3111 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1260) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3110 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1261) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3109 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1262) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3108 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1263) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3107 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1264) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3106 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3388), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1265) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3105 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3104 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1266) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3103 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1267) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3102 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1268) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3101 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1269) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3100 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1270) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3099 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1271) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3098 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1272) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3097 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3387), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1273) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3096 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3095 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1274) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3094 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1275) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3093 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1276) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3092 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1277) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3091 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1278) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3090 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1279) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3089 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1280) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3088 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3386), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1281) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3087 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3086 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1282) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3085 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1283) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3084 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1284) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3083 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1285) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3082 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1286) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3081 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1287) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3080 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1288) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3079 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3385), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1289) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3078 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3077 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1290) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3076 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1291) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3075 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1292) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3074 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1293) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3073 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1294) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3072 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1295) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3071 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1296) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3070 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1297) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3069 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3068 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1298) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3067 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1299) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3066 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1300) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3065 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1301) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3064 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1302) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3063 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1303) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3062 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1304) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3061 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1305) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3060 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3059 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1306) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3058 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1307) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3057 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1308) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3056 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1309) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3055 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1310) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3054 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1311) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3053 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1312) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3052 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1313) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3051 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3050 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1314) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3049 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1315) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3048 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1316) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3047 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1317) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3046 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1318) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3045 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1319) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3044 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1320) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3043 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1321) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3042 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3041 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1322) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3040 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1323) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3039 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1324) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3038 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1325) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3037 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1326) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3036 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1327) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3035 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1328) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3034 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1329) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3033 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3032 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1330) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3031 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1331) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3030 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1332) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3029 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1333) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3028 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1334) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3027 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1335) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3026 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1336) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3025 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1337) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3024 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3378), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3023 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1338) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3022 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1339) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3021 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1340) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3020 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1341) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3019 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1342) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3018 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1343) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3017 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1344) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3016 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1345) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3015 ( .A(
        oc8051_ram_top1_wr_addr_m_6_), .B(oc8051_ram_top1_wr_addr_m_5_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3219) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3014 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3219), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3163), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3013 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3012 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1346) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3011 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1347) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3010 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1348) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3009 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1349) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3008 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1350) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3007 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1351) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3006 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1352) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3005 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1353) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3004 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3003 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1354) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3002 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1355) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3001 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1356) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3000 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1357) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2999 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1358) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2998 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1359) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2997 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1360) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2996 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1361) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2995 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2994 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1362) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2993 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1363) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2992 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1364) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2991 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1365) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2990 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1366) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2989 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1367) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2988 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1368) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2987 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1369) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2986 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2985 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1370) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2984 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1371) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2983 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1372) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2982 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1373) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2981 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1374) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2980 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1375) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2979 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1376) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2978 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1377) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2977 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2976 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1378) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2975 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1379) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2974 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1380) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2973 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1381) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2972 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1382) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2971 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1383) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2970 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1384) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2969 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1385) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2968 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2967 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1386) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2966 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1387) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2965 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1388) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2964 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1389) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2963 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1390) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2962 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1391) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2961 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1392) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2960 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1393) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2959 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2958 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1394) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2957 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1395) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2956 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1396) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2955 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1397) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2954 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1398) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2953 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1399) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2952 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1400) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2951 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1401) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2950 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2949 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1402) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2948 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1403) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2947 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1404) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2946 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1405) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2945 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1406) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2944 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1407) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2943 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1408) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2942 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1409) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2941 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2940 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1410) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2939 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1411) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2938 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1412) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2937 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1413) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2936 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1414) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2935 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1415) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2934 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1416) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2933 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1417) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2932 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2931 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1418) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2930 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1419) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2929 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1420) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2928 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1421) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2927 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1422) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2926 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1423) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2925 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1424) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2924 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1425) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2923 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2922 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1426) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2921 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1427) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2920 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1428) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2919 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1429) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2918 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1430) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2917 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1431) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2916 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1432) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2915 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1433) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2914 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2913 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1434) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2912 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1435) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2911 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1436) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2910 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1437) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2909 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1438) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2908 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1439) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2907 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1440) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2906 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1441) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2905 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2904 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1442) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2903 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1443) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2902 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1444) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2901 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1445) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2900 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1446) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2899 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1447) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2898 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1448) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2897 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1449) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2896 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2895 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1450) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2894 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1451) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2893 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1452) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2892 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1453) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2891 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1454) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2890 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1455) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2889 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1456) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2888 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1457) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2887 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2886 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1458) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2885 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1459) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2884 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1460) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2883 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1461) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2882 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1462) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2881 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1463) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2880 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1464) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2879 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1465) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2878 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3361), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2877 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1466) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2876 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1467) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2875 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1468) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2874 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1469) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2873 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1470) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2872 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1471) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2871 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1472) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2870 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1473) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2869 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3219), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3183), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2868 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2867 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1474) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2866 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1475) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2865 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1476) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2864 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1477) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2863 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1478) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2862 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1479) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2861 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1480) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2860 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1481) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2859 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2858 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1482) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2857 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1483) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2856 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1484) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2855 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1485) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2854 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1486) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2853 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1487) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2852 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1488) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2851 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1489) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2850 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2849 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1490) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2848 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1491) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2847 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1492) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2846 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1493) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2845 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1494) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2844 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1495) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2843 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1496) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2842 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1497) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2841 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2840 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1498) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2839 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1499) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2838 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1500) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2837 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1501) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2836 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1502) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2835 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1503) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2834 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1504) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2833 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1505) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2832 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2831 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1506) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2830 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1507) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2829 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1508) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2828 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1509) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2827 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1510) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2826 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1511) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2825 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1512) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2824 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1513) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2823 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2822 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1514) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2821 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1515) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2820 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1516) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2819 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1517) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2818 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1518) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2817 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1519) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2816 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1520) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2815 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1521) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2814 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2813 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1522) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2812 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1523) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2811 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1524) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2810 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1525) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2809 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1526) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2808 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1527) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2807 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1528) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2806 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1529) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2805 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2804 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1530) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2803 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1531) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2802 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1532) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2801 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1533) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2800 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1534) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2799 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1535) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2798 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1536) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2797 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1537) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2796 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2795 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1538) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2794 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1539) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2793 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1540) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2792 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1541) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2791 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1542) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2790 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1543) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2789 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1544) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2788 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1545) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2787 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2786 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1546) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2785 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1547) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2784 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1548) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2783 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1549) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2782 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1550) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2781 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1551) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2780 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1552) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2779 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1553) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2778 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2777 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1554) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2776 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1555) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2775 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1556) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2774 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1557) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2773 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1558) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2772 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1559) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2771 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1560) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2770 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1561) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2769 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2768 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1562) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2767 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1563) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2766 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1564) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2765 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1565) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2764 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1566) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2763 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1567) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2762 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1568) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2761 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1569) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2760 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2759 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1570) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2758 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1571) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2757 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1572) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2756 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1573) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2755 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1574) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2754 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1575) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2753 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1576) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2752 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3347), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1577) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2751 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2750 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1578) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2749 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1579) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2748 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1580) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2747 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1581) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2746 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1582) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2745 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1583) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2744 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1584) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2743 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3346), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1585) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2742 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2741 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1586) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2740 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1587) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2739 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1588) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2738 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1589) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2737 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1590) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2736 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1591) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2735 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1592) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2734 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3345), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1593) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2733 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3344), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2732 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1594) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2731 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1595) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2730 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1596) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2729 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1597) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2728 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1598) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2727 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1599) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2726 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1600) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2725 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3343), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1601) );
  AND3_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2724 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3324), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3342), .C(wr_addr[7]), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3237) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2723 ( .A(
        oc8051_ram_top1_wr_addr_m_5_), .B(oc8051_ram_top1_wr_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3182) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2722 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3237), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3182), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2721 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2720 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1602) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2719 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1603) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2718 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1604) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2717 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1605) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2716 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1606) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2715 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1607) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2714 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1608) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2713 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3341), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1609) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2712 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2711 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1610) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2710 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1611) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2709 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1612) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2708 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1613) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2707 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1614) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2706 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1615) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2705 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1616) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2704 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3340), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1617) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2703 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2702 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1618) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2701 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1619) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2700 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1620) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2699 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1621) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2698 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1622) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2697 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1623) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2696 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1624) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2695 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3339), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1625) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2694 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2693 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1626) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2692 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1627) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2691 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1628) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2690 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1629) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2689 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1630) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2688 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1631) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2687 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1632) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2686 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3338), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1633) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2685 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2684 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1634) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2683 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1635) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2682 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1636) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2681 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1637) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2680 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1638) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2679 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1639) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2678 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1640) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2677 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3337), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1641) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2676 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2675 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1642) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2674 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1643) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2673 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1644) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2672 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1645) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2671 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1646) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2670 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1647) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2669 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1648) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2668 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3336), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1649) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2667 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2666 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1650) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2665 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1651) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2664 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1652) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2663 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1653) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2662 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1654) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2661 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1655) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2660 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1656) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2659 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3335), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1657) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2658 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2657 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1658) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2656 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1659) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2655 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1660) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2654 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1661) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2653 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1662) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2652 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1663) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2651 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1664) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2650 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3334), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1665) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2649 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2648 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1666) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2647 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1667) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2646 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1668) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2645 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1669) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2644 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1670) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2643 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1671) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2642 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1672) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2641 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3333), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1673) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2640 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2639 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1674) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2638 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1675) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2637 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1676) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2636 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1677) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2635 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1678) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2634 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1679) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2633 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1680) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2632 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3332), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1681) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2631 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2630 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1682) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2629 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1683) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2628 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1684) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2627 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1685) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2626 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1686) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2625 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1687) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2624 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1688) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2623 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3331), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1689) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2622 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2621 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1690) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2620 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1691) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2619 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1692) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2618 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1693) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2617 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1694) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2616 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1695) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2615 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1696) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2614 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3330), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1697) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2613 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2612 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1698) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2611 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1699) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2610 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1700) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2609 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1701) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2608 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1702) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2607 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1703) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2606 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1704) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2605 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3329), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1705) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2604 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2603 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1706) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2602 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1707) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2601 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1708) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2600 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1709) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2599 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1710) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2598 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1711) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2597 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1712) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2596 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3328), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1713) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2595 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2594 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1714) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2593 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1715) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2592 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1716) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2591 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1717) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2590 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1718) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2589 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1719) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2588 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1720) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2587 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3327), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1721) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2586 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3326), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2585 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1722) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2584 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1723) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2583 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1724) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2582 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1725) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2581 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1726) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2580 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1727) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2579 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1728) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2578 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3325), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1729) );
  AND3_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2577 ( .A(
        oc8051_ram_top1_wr_addr_m_4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3324), .C(wr_addr[7]), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3218) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2576 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3218), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3182), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2575 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2574 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1730) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2573 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1731) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2572 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1732) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2571 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1733) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2570 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1734) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2569 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1735) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2568 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1736) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2567 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3323), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1737) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2566 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2565 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1738) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2564 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1739) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2563 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1740) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2562 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1741) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2561 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1742) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2560 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1743) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2559 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1744) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2558 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3322), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1745) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2557 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2556 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1746) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2555 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1747) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2554 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1748) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2553 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1749) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2552 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1750) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2551 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1751) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2550 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1752) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2549 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3321), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1753) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2548 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2547 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1754) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2546 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1755) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2545 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1756) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2544 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1757) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2543 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1758) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2542 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1759) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2541 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1760) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2540 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3320), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1761) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2539 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2538 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1762) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2537 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1763) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2536 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1764) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2535 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1765) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2534 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1766) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2533 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1767) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2532 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1768) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2531 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3319), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1769) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2530 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2529 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1770) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2528 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1771) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2527 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1772) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2526 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1773) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2525 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1774) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2524 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1775) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2523 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1776) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2522 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3318), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1777) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2521 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2520 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1778) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2519 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1779) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2518 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1780) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2517 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1781) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2516 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1782) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2515 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1783) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2514 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1784) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2513 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3317), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1785) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2512 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2511 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1786) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2510 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1787) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2509 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1788) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2508 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1789) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2507 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1790) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2506 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1791) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2505 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1792) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2504 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3316), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1793) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2503 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2502 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1794) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2501 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1795) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2500 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1796) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2499 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1797) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2498 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1798) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2497 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1799) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2496 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1800) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2495 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3315), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1801) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2494 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2493 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1802) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2492 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1803) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2491 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1804) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2490 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1805) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2489 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1806) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2488 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1807) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2487 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1808) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2486 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3314), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1809) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2485 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2484 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1810) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2483 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1811) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2482 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1812) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2481 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1813) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2480 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1814) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2479 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1815) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2478 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1816) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2477 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3313), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1817) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2476 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2475 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1818) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2474 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1819) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2473 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1820) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2472 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1821) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2471 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1822) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2470 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1823) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2469 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1824) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2468 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3312), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1825) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2467 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2466 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1826) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2465 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1827) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2464 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1828) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2463 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1829) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2462 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1830) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2461 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1831) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2460 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1832) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2459 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3311), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1833) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2458 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2457 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1834) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2456 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1835) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2455 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1836) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2454 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1837) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2453 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1838) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2452 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1839) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2451 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1840) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2450 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3310), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1841) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2449 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2448 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1842) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2447 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1843) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2446 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1844) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2445 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1845) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2444 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1846) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2443 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1847) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2442 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1848) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2441 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3309), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1849) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2440 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3308), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2439 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1850) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2438 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1851) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2437 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1852) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2436 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1853) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2435 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1854) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2434 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1855) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2433 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1856) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2432 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1857) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2431 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3237), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3164), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2430 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2429 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1858) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2428 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1859) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2427 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1860) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2426 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1861) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2425 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1862) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2424 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1863) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2423 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1864) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2422 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1865) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2421 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2420 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1866) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2419 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1867) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2418 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1868) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2417 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1869) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2416 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1870) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2415 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1871) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2414 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1872) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2413 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1873) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2412 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2411 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1874) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2410 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1875) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2409 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1876) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2408 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1877) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2407 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1878) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2406 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1879) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2405 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1880) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2404 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1881) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2403 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2402 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1882) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2401 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1883) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2400 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1884) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2399 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1885) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2398 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1886) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2397 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1887) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2396 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1888) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2395 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1889) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2394 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2393 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1890) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2392 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1891) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2391 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1892) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2390 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1893) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2389 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1894) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2388 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1895) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2387 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1896) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2386 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1897) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2385 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2384 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1898) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2383 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1899) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2382 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1900) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2381 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1901) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2380 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1902) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2379 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1903) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2378 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1904) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2377 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1905) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2376 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2375 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1906) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2374 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1907) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2373 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1908) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2372 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1909) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2371 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1910) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2370 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1911) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2369 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1912) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2368 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1913) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2367 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2366 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1914) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2365 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1915) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2364 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1916) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2363 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1917) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2362 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1918) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2361 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1919) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2360 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1920) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2359 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1921) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2358 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2357 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1922) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2356 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1923) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2355 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1924) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2354 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1925) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2353 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1926) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2352 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1927) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2351 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1928) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2350 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1929) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2349 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2348 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1930) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2347 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1931) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2346 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1932) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2345 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1933) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2344 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1934) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2343 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1935) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2342 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1936) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2341 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1937) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2340 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2339 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1938) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2338 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1939) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2337 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1940) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2336 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1941) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2335 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1942) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2334 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1943) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2333 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1944) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2332 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1945) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2331 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2330 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1946) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2329 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1947) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2328 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1948) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2327 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1949) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2326 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1950) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2325 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1951) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2324 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1952) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2323 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1953) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2322 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2321 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1954) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2320 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1955) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2319 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1956) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2318 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1957) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2317 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1958) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2316 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1959) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2315 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1960) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2314 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1961) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2313 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2312 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1962) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2311 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1963) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2310 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1964) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2309 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1965) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2308 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1966) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2307 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1967) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2306 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1968) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2305 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1969) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2304 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2303 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1970) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2302 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1971) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2301 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1972) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2300 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1973) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2299 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1974) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2298 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1975) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2297 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1976) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2296 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1977) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2295 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3291), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2294 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1978) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2293 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1979) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2292 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1980) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2291 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1981) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2290 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1982) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2289 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1983) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2288 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1984) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2287 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1985) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2286 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3218), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3164), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2285 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2284 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1986) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2283 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1987) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2282 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1988) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2281 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1989) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2280 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1990) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2279 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1991) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2278 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1992) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2277 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1993) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2276 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2275 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1994) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2274 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1995) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2273 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1996) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2272 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1997) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2271 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1998) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2270 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1999) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2269 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2000) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2268 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2001) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2267 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2266 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2002) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2265 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2003) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2264 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2004) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2263 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2005) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2262 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2006) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2261 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2007) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2260 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2008) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2259 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2009) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2258 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2257 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2010) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2256 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2011) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2255 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2012) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2254 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2013) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2253 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2014) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2252 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2015) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2251 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2016) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2250 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2017) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2249 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2248 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2018) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2247 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2019) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2246 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2020) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2245 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2021) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2244 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2022) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2243 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2023) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2242 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2024) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2241 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2025) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2240 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2239 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2026) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2238 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2027) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2237 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2028) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2236 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2029) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2235 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2030) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2234 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2031) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2233 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2032) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2232 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2033) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2231 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2230 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2034) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2229 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2035) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2228 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2036) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2227 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2037) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2226 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2038) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2225 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2039) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2224 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2040) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2223 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2041) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2222 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2221 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2042) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2220 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2043) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2219 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2044) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2218 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2045) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2217 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2046) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2216 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2047) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2215 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2048) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2214 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2049) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2213 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2212 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2050) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2211 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2051) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2210 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2052) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2209 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2053) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2208 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2054) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2207 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2055) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2206 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2056) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2205 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2057) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2204 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2203 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2058) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2202 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2059) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2201 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2060) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2200 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2061) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2199 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2062) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2198 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2063) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2197 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2064) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2196 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2065) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2195 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2194 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2066) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2193 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2067) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2192 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2068) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2191 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2069) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2190 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2070) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2189 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2071) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2188 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2072) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2187 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2073) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2186 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2185 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2074) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2184 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2075) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2183 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2076) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2182 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2077) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2181 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2078) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2180 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2079) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2179 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2080) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2178 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2081) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2177 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2176 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2082) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2175 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2083) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2174 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2084) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2173 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2085) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2172 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2086) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2171 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2087) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2170 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2088) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2169 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2089) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2168 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2167 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2090) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2166 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2091) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2165 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2092) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2164 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2093) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2163 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2094) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2162 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2095) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2161 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2096) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2160 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2097) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2159 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2158 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2098) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2157 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2099) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2156 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2100) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2155 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2101) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2154 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2102) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2153 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2103) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2152 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2104) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2151 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2105) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2150 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3274), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2149 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2106) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2148 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2107) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2147 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2108) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2146 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2109) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2145 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2110) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2144 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2111) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2143 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2112) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2142 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2113) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2141 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3255), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3237), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2140 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2139 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2114) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2138 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2115) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2137 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2116) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2136 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2117) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2135 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2118) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2134 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2119) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2133 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2120) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2132 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2121) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2131 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2130 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2122) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2129 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2123) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2128 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2124) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2127 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2125) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2126 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2126) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2125 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2127) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2124 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2128) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2123 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2129) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2122 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2121 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2130) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2120 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2131) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2119 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2132) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2118 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2133) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2117 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2134) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2116 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2135) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2115 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2136) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2114 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2137) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2113 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2112 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2138) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2111 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2139) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2110 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2140) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2109 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2141) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2108 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2142) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2107 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2143) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2106 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2144) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2105 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2145) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2104 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2103 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2146) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2102 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2147) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2101 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2148) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2100 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2149) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2099 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2150) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2098 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2151) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2097 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2152) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2096 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2153) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2095 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2094 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2154) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2093 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2155) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2092 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2156) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2091 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2157) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2090 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2158) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2089 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2159) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2088 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2160) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2087 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2161) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2086 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2085 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2162) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2084 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2163) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2083 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2164) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2082 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2165) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2081 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2166) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2080 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2167) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2079 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2168) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2078 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2169) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2077 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2076 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2170) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2075 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2171) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2074 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2172) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2073 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2173) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2072 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2174) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2071 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2175) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2070 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2176) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2069 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2177) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2068 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2067 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2178) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2066 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2179) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2065 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2180) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2064 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2181) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2063 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2182) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2062 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2183) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2061 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2184) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2060 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2185) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2059 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2058 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2186) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2057 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2187) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2056 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2188) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2055 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2189) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2054 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2190) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2053 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2191) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2052 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2192) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2051 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2193) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2050 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2049 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2194) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2048 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2195) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2047 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2196) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2046 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2197) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2045 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2198) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2044 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2199) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2043 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2200) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2042 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2201) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2041 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2040 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2202) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2039 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2203) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2038 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2204) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2037 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2205) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2036 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2206) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2035 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2207) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2034 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2208) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2033 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2209) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2032 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2031 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2210) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2030 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2211) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2029 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2212) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2028 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2213) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2027 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2214) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2026 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2215) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2025 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2216) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2024 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2217) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2023 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2022 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2218) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2021 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2219) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2020 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2220) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2019 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2221) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2018 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2222) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2017 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2223) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2016 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2224) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2015 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2225) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2014 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2013 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2226) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2012 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2227) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2011 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2228) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2010 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2229) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2009 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2230) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2008 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2231) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2007 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2232) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2006 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2233) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2005 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3257), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2004 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2234) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2003 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2235) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2002 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2236) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2001 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2237) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2000 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2238) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1999 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2239) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1998 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2240) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1997 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2241) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1996 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3255), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3218), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1995 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1994 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2242) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1993 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2243) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1992 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2244) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1991 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2245) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1990 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2246) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1989 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2247) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1988 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2248) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1987 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2249) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1986 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1985 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2250) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1984 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2251) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1983 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2252) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1982 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2253) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1981 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2254) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1980 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2255) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1979 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2256) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1978 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2257) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1977 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1976 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2258) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1975 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2259) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1974 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2260) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1973 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2261) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1972 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2262) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1971 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2263) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1970 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2264) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1969 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2265) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1968 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1967 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2266) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1966 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2267) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1965 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2268) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1964 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2269) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1963 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2270) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1962 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2271) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1961 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2272) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1960 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2273) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1959 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1958 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2274) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1957 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2275) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1956 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2276) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1955 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2277) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1954 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2278) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1953 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2279) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1952 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2280) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1951 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2281) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1950 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1949 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2282) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1948 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2283) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1947 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2284) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1946 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2285) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1945 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2286) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1944 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2287) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1943 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2288) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1942 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2289) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1941 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1940 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2290) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1939 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2291) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1938 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2292) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1937 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2293) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1936 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2294) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1935 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2295) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1934 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2296) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1933 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2297) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1932 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1931 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2298) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1930 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2299) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1929 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2300) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1928 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2301) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1927 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2302) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1926 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2303) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1925 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2304) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1924 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2305) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1923 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1922 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2306) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1921 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2307) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1920 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2308) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1919 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2309) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1918 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2310) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1917 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2311) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1916 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2312) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1915 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2313) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1914 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1913 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2314) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1912 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2315) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1911 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2316) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1910 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2317) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1909 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2318) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1908 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2319) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1907 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2320) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1906 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2321) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1905 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1904 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2322) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1903 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2323) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1902 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2324) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1901 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2325) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1900 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2326) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1899 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2327) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1898 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2328) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1897 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2329) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1896 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1895 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2330) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1894 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2331) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1893 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2332) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1892 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2333) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1891 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2334) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1890 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2335) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1889 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2336) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1888 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2337) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1887 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1886 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2338) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1885 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2339) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1884 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2340) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1883 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2341) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1882 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2342) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1881 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2343) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1880 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2344) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1879 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2345) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1878 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1877 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2346) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1876 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2347) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1875 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2348) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1874 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2349) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1873 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2350) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1872 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2351) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1871 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2352) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1870 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2353) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1869 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1868 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2354) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1867 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2355) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1866 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2356) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1865 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2357) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1864 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2358) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1863 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2359) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1862 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2360) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1861 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2361) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1860 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3239), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1859 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2362) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1858 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2363) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1857 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2364) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1856 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2365) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1855 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2366) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1854 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2367) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1853 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2368) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1852 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2369) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1851 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3237), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3219), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1850 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1849 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2370) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1848 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2371) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1847 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2372) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1846 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2373) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1845 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2374) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1844 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2375) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1843 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2376) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1842 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2377) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1841 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1840 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2378) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1839 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2379) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1838 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2380) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1837 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2381) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1836 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2382) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1835 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2383) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1834 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2384) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1833 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2385) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1832 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1831 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2386) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1830 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2387) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1829 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2388) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1828 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2389) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1827 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2390) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1826 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2391) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1825 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2392) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1824 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2393) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1823 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1822 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2394) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1821 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2395) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1820 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2396) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1819 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2397) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1818 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2398) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1817 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2399) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1816 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2400) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1815 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2401) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1814 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1813 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2402) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1812 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2403) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1811 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2404) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1810 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2405) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1809 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2406) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1808 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2407) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1807 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2408) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1806 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2409) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1805 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1804 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2410) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1803 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2411) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1802 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2412) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1801 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2413) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1800 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2414) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1799 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2415) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1798 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2416) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1797 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2417) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1796 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1795 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2418) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1794 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2419) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1793 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2420) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1792 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2421) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1791 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2422) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1790 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2423) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1789 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2424) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1788 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3230), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2425) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1787 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1786 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2426) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1785 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2427) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1784 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2428) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1783 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2429) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1782 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2430) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1781 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2431) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1780 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2432) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1779 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3229), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2433) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1778 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1777 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2434) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1776 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2435) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1775 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2436) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1774 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2437) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1773 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2438) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1772 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2439) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1771 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2440) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1770 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3228), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2441) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1769 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1768 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2442) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1767 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2443) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1766 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2444) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1765 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2445) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1764 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2446) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1763 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2447) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1762 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2448) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1761 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3227), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2449) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1760 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1759 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2450) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1758 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2451) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1757 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2452) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1756 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2453) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1755 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2454) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1754 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2455) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1753 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2456) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1752 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3226), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2457) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1751 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1750 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2458) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1749 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2459) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1748 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2460) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1747 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2461) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1746 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2462) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1745 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2463) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1744 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2464) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1743 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3225), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2465) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1742 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1741 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2466) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1740 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2467) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1739 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2468) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1738 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2469) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1737 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2470) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1736 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2471) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1735 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2472) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1734 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3224), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2473) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1733 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1732 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2474) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1731 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2475) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1730 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2476) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1729 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2477) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1728 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2478) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1727 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2479) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1726 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2480) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1725 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3223), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2481) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1724 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1723 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2482) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1722 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2483) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1721 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2484) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1720 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2485) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1719 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2486) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1718 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2487) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1717 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2488) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1716 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3222), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2489) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1715 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3221), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1714 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2490) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1713 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2491) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1712 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2492) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1711 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2493) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1710 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2494) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1709 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2495) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1708 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2496) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1707 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3220), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2497) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1706 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3218), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3219), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1705 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1704 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2498) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1703 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2499) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1702 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2500) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1701 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2501) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1700 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2502) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1699 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2503) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1698 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2504) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1697 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3217), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2505) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1696 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1695 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2506) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1694 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2507) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1693 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2508) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1692 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2509) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1691 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2510) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1690 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2511) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1689 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2512) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1688 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3216), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2513) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1687 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1686 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2514) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1685 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2515) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1684 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2516) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1683 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2517) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1682 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2518) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1681 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2519) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1680 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2520) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1679 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3215), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2521) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1678 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1677 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2522) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1676 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2523) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1675 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2524) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1674 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2525) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1673 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2526) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1672 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2527) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1671 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2528) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1670 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3214), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2529) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1669 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1668 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2530) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1667 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2531) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1666 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2532) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1665 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2533) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1664 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2534) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1663 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2535) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1662 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2536) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1661 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3213), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2537) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1660 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1659 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2538) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1658 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2539) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1657 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2540) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1656 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2541) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1655 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2542) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1654 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2543) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1653 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2544) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1652 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3212), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2545) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1651 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1650 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2546) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1649 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2547) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1648 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2548) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1647 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2549) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1646 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2550) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1645 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2551) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1644 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2552) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1643 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3211), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2553) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1642 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1641 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2554) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1640 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2555) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1639 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2556) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1638 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2557) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1637 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2558) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1636 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2559) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1635 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2560) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1634 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2561) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1633 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1632 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2562) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1631 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2563) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1630 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2564) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1629 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2565) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1628 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2566) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1627 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2567) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1626 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2568) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1625 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2569) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1624 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1623 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2570) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1622 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2571) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1621 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2572) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1620 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2573) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1619 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2574) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1618 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2575) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1617 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2576) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1616 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2577) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1615 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1614 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2578) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1613 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2579) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1612 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2580) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1611 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2581) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1610 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2582) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1609 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2583) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1608 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2584) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1607 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2585) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1606 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1605 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2586) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1604 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2587) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1603 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2588) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1602 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2589) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1601 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2590) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1600 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2591) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1599 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2592) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1598 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2593) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1597 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1596 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2594) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1595 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2595) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1594 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2596) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1593 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2597) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1592 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2598) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1591 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2599) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1590 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2600) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1589 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2601) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1588 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1587 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2602) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1586 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2603) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1585 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2604) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1584 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2605) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1583 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2606) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1582 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2607) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1581 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2608) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1580 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2609) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1579 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1578 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2610) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1577 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2611) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1576 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2612) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1575 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2613) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1574 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2614) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1573 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2615) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1572 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2616) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1571 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2617) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1570 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3202), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1569 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2618) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1568 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2619) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1567 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2620) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1566 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2621) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1565 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2622) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1564 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2623) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1563 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2624) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1562 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2625) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1561 ( .A(
        oc8051_ram_top1_oc8051_idata__logic1_), .B(oc8051_ram_top1_n53), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1560 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4110), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n570) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1559 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4010), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n571) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1558 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3910), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n572) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1557 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3810), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n573) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1556 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3710), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n574) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1555 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3610), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n575) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1554 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3510), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n576) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1553 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3435), .S0(
        oc8051_ram_top1_n53), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n577) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1552 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3182), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3163), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1551 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1550 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n578) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1549 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n579) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1548 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n580) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1547 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n581) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1546 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n582) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1545 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n583) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1544 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n584) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1543 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3200), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n585) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1542 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1541 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n586) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1540 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n587) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1539 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n588) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1538 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n589) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1537 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n590) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1536 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n591) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1535 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n592) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1534 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3199), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n593) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1533 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1532 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n594) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1531 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n595) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1530 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n596) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1529 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n597) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1528 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n598) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1527 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n599) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1526 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n600) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1525 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3198), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n601) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1524 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1523 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n602) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1522 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n603) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1521 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n604) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1520 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n605) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1519 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n606) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1518 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n607) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1517 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n608) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1516 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3197), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n609) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1515 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1514 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n610) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1513 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n611) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1512 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n612) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1511 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n613) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1510 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n614) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1509 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n615) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1508 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n616) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1507 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3196), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n617) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1506 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1505 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n618) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1504 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n619) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1503 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n620) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1502 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n621) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1501 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n622) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1500 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n623) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1499 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n624) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1498 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3195), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n625) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1497 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1496 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n626) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1495 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n627) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1494 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n628) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1493 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n629) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1492 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n630) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1491 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n631) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1490 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n632) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1489 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3194), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n633) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1488 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1487 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n634) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1486 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n635) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1485 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n636) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1484 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n637) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1483 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n638) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1482 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n639) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1481 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n640) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1480 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3193), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n641) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1479 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1478 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n642) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1477 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n643) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1476 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n644) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1475 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n645) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1474 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n646) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1473 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n647) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1472 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n648) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1471 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3192), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n649) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1470 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1469 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n650) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1468 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n651) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1467 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n652) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1466 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n653) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1465 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n654) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1464 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n655) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1463 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n656) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1462 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3191), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n657) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1461 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1460 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n658) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1459 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n659) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1458 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n660) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1457 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n661) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1456 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n662) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1455 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n663) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1454 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n664) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1453 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3190), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n665) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1452 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1451 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n666) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1450 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n667) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1449 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n668) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1448 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n669) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1447 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n670) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1446 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n671) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1445 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n672) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1444 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3189), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n673) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1443 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1442 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n674) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1441 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n675) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1440 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n676) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1439 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n677) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1438 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n678) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1437 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n679) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1436 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n680) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1435 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3188), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n681) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1434 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1433 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n682) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1432 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n683) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1431 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n684) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1430 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n685) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1429 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n686) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1428 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n687) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1427 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n688) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1426 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3187), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n689) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1425 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1424 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n690) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1423 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n691) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1422 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n692) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1421 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n693) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1420 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n694) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1419 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n695) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1418 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n696) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1417 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3186), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n697) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1416 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3185), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1415 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n698) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1414 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n699) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1413 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n700) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1412 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n701) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1411 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n702) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1410 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n703) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1409 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n704) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1408 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3184), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n705) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1407 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3182), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3183), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1406 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1405 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n706) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1404 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n707) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1403 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n708) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1402 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n709) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1401 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n710) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1400 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n711) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1399 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n712) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1398 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3181), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n713) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1397 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1396 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n714) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1395 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n715) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1394 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n716) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1393 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n717) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1392 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n718) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1391 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n719) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1390 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n720) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1389 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n721) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1388 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1387 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n722) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1386 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n723) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1385 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n724) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1384 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n725) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1383 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n726) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1382 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n727) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1381 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n728) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1380 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n729) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1379 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1378 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n730) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1377 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n731) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1376 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n732) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1375 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n733) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1374 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n734) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1373 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n735) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1372 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n736) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1371 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n737) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1370 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1369 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n738) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1368 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n739) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1367 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n740) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1366 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n741) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1365 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n742) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1364 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n743) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1363 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n744) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1362 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n745) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1361 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1360 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n746) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1359 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n747) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1358 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n748) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1357 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n749) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1356 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n750) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1355 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n751) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1354 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n752) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1353 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n753) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1352 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1351 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n754) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1350 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n755) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1349 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n756) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1348 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n757) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1347 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n758) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1346 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n759) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1345 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n760) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1344 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n761) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1343 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1342 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n762) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1341 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n763) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1340 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n764) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1339 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n765) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1338 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n766) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1337 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n767) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1336 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n768) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1335 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n769) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1334 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1333 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n770) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1332 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n771) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1331 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n772) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1330 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n773) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1329 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n774) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1328 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n775) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1327 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n776) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1326 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n777) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1325 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1324 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n778) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1323 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n779) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1322 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n780) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1321 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n781) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1320 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n782) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1319 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n783) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1318 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n784) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1317 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n785) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1316 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1315 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n786) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1314 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n787) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1313 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n788) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1312 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n789) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1311 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n790) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1310 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n791) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1309 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n792) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1308 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n793) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1307 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1306 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n794) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1305 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n795) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1304 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n796) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1303 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n797) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1302 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n798) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1301 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n799) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1300 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n800) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1299 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3170), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n801) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1298 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1297 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n802) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1296 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n803) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1295 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n804) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1294 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n805) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1293 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n806) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1292 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n807) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1291 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n808) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1290 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3169), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n809) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1289 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1288 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n810) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1287 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n811) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1286 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n812) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1285 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n813) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1284 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n814) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1283 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n815) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1282 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n816) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1281 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3168), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n817) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1280 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1279 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n818) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1278 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n819) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1277 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n820) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1276 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n821) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1275 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n822) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1274 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n823) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1273 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n824) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1272 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3167), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n825) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1271 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3166), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1270 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n826) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1269 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n827) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1268 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n828) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1267 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n829) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1266 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n830) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1265 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n831) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1264 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n832) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1263 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3165), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n833) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1262 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3163), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3164), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1261 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1260 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n834) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1259 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n835) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1258 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n836) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1257 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n837) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1256 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n838) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1255 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n839) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1254 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n840) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1253 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3162), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n841) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1252 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1251 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n842) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1250 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n843) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1249 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n844) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1248 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n845) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1247 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n846) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1246 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n847) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1245 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n848) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1244 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3161), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n849) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1243 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1242 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n850) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1241 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n851) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1240 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n852) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1239 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n853) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1238 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n854) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1237 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n855) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1236 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n856) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1235 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3160), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n857) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1234 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1233 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n858) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1232 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n859) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1231 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n860) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1230 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n861) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1229 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n862) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1228 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n863) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1227 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n864) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1226 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3159), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n865) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1225 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3158), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1224 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n866) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1223 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n867) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1222 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n868) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1221 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n869) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1220 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n870) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1219 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n871) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1218 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n872) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1217 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3157), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n873) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1216 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3156), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1215 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n874) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1214 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n875) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1213 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n876) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1212 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n877) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1211 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n878) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1210 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n879) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1209 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n880) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1208 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3155), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n881) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1207 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3154), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1206 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n882) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1205 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n883) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1204 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n884) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1203 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n885) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1202 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n886) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1201 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n887) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1200 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n888) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1199 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3153), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n889) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1198 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3152), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1197 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n890) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1196 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n891) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1195 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n892) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1194 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n893) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1193 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n894) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1192 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n895) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1191 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n896) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1190 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3151), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n897) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1189 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3150), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1188 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n898) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1187 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n899) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1186 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n900) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1185 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n901) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1184 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n902) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1183 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n903) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1182 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n904) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1181 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n905) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1180 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3148), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1179 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n906) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1178 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n907) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1177 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n908) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1176 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n909) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1175 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n910) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1174 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n911) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1173 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n912) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1172 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n913) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1171 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3146), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1170 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n914) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1169 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n915) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1168 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n916) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1167 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n917) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1166 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n918) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1165 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n919) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1164 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n920) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1163 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n921) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1162 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3144), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1161 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n922) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1160 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n923) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1159 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n924) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1158 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n925) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1157 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n926) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1156 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n927) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1155 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n928) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1154 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n929) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1153 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3142), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1152 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n930) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1151 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n931) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1150 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n932) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1149 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n933) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1148 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n934) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1147 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n935) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1146 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n936) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1145 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n937) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1144 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3140), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1143 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n938) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1142 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n939) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1141 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n940) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1140 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n941) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1139 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n942) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1138 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n943) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1137 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n944) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1136 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3139), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n945) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1135 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3138), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1134 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n946) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1133 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n947) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1132 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n948) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1131 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n949) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1130 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n950) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1129 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n951) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1128 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n952) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1127 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3137), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n953) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1126 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3135), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3136), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1125 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n954) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1124 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n955) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1123 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n956) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1122 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n957) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1121 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n958) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1120 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n959) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1119 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n960) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1118 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3134), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n961) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1117 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3133), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1116 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n962) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1115 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n963) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1114 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n964) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1113 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n965) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1112 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n966) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1111 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n967) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1110 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n968) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1109 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3132), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n969) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1108 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3131), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1107 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n970) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1106 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n971) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1105 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n972) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1104 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n973) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1103 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n974) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1102 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n975) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1101 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n976) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1100 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3130), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n977) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1099 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3129), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1098 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n978) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1097 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n979) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1096 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n980) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1095 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n981) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1094 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n982) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1093 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n983) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1092 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n984) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1091 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3128), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n985) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1090 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3126), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3127), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1089 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n986) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1088 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n987) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1087 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n988) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1086 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n989) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1085 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n990) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1084 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n991) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1083 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n992) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1082 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3125), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n993) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1081 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n994) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1080 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n995) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1079 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n996) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1078 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n997) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1077 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n998) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1076 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3124), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n999) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1075 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3041) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1074 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3043) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1073 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3044) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1072 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3041), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3042), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3043), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3044), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3040) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1071 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3081) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1070 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3083) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1069 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3084) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1068 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3081), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3082), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3083), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3084), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3080) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1067 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2957) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1066 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2959) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1065 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2960) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1064 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2957), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2958), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2959), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2960), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2956) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1063 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2997) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1062 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2999) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1061 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3000) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1060 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2997), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2998), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2999), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3000), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2996) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1059 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2873) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1058 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2875) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1057 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2876) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1056 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2873), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2874), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2875), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2876), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2872) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1055 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2913) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1054 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2915) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1053 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2916) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1052 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2913), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2914), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2915), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2916), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2912) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1051 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2789) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1050 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2791) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1049 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2792) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1048 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2789), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2790), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2791), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2792), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2788) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1047 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2829) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1046 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2831) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1045 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2832) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1044 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2829), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2830), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2831), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2832), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2828) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1043 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2705) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1042 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2707) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1041 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2708) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1040 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2705), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2706), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2707), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2708), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2704) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1039 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2745) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1038 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2747) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1037 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2748) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1036 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2745), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2746), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2747), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2748), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2744) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1035 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n564) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1034 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n566) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1033 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n567) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1032 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n564), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n565), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n566), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n567), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n563) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1031 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2661) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1030 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2663) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1029 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2664) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1028 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2661), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2662), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2663), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2664), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2660) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1027 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n480) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1026 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n482) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1025 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n483) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1024 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n480), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n481), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n482), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n483), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n479) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1023 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n520) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1022 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n522) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1021 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n523) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1020 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n520), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n521), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n522), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n523), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n519) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1019 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n396) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1018 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n398) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1017 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n399) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1016 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n396), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n397), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n398), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n399), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n395) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1015 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n436) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1014 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n438) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1013 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n439) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1012 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n436), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n437), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n438), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n439), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n435) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1011 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3104) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1010 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3114) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1009 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3119) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1008 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3064) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1007 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3074) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1006 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3079) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1005 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3020) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1004 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3030) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1003 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3035) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1002 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2980) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1001 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2990) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u1000 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2995) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u999 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2936) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u998 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2946) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u997 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2951) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u996 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2896) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u995 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2906) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u994 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2911) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u993 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2852) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u992 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2862) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u991 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2867) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u990 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2812) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u989 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2822) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u988 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2827) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u987 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2768) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u986 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2778) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u985 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2783) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u984 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2728) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u983 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2738) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u982 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2743) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u981 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2684) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u980 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2694) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u979 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2699) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u978 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2644) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u977 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2654) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u976 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2659) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u975 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n543) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u974 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n553) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u973 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n558) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u972 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n503) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u971 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n513) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u970 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n518) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u969 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n459) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u968 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n469) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u967 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n474) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u966 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n419) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u965 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n429) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u964 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n434) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u963 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3051) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u962 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3053) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u961 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3054) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u960 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3051), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3052), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3053), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3054), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3050) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u959 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3091) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u958 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3093) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u957 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3094) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u956 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3091), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3092), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3093), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3094), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3090) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u955 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2967) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u954 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2969) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u953 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2970) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u952 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2967), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2968), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2969), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2970), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2966) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u951 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3007) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u950 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3009) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u949 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3010) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u948 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3007), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3008), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3009), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3010), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3006) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u947 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2883) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u946 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2885) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u945 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2886) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u944 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2883), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2884), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2885), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2886), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2882) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u943 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2923) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u942 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2925) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u941 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2926) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u940 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2923), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2924), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2925), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2926), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2922) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u939 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2799) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u938 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2801) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u937 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2802) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u936 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2799), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2800), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2801), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2802), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2798) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u935 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2839) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u934 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2841) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u933 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2842) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u932 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2839), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2840), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2841), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2842), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2838) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u931 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2715) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u930 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2717) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u929 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2718) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u928 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2715), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2716), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2717), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2718), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2714) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u927 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2755) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u926 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2757) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u925 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2758) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u924 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2755), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2756), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2757), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2758), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2754) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u923 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2631) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u922 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2633) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u921 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2634) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u920 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2631), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2632), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2633), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2634), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2630) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u919 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2671) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u918 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2673) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u917 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2674) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u916 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2671), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2672), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2673), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2674), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2670) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u915 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n490) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u914 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n492) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u913 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n493) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u912 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n490), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n491), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n492), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n493), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n489) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u911 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n530) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u910 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n532) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u909 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n533) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u908 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n530), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n531), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n532), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n533), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n529) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u907 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n406) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u906 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n408) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u905 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n409) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u904 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n406), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n407), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n408), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n409), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n405) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u903 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n446) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u902 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n448) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u901 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n449) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u900 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n446), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n447), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n448), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n449), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n445) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u899 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3103) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u898 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3113) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u897 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3118) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u896 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3063) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u895 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3073) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u894 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3078) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u893 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3019) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u892 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3029) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u891 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3034) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u890 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2979) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u889 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2989) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u888 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2994) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u887 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2935) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u886 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2945) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u885 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2950) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u884 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2895) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u883 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2905) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u882 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2910) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u881 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2851) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u880 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2861) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u879 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2866) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u878 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2811) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u877 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2821) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u876 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2826) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u875 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2767) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u874 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2777) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u873 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2782) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u872 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2727) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u871 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2737) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u870 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2742) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u869 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2683) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u868 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2693) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u867 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2698) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u866 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2643) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u865 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2653) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u864 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2658) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u863 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n542) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u862 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n552) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u861 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n557) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u860 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n502) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u859 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n512) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u858 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n517) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u857 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n458) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u856 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n468) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u855 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n473) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u854 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n418) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u853 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n428) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u852 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n433) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u851 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3056) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u850 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3058) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u849 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3059) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u848 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3056), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3057), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3058), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3059), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3055) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u847 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3096) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u846 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3098) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u845 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3099) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u844 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3096), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3097), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3098), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3099), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3095) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u843 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2972) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u842 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2974) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u841 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2975) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u840 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2972), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2973), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2974), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2975), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2971) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u839 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3012) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u838 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3014) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u837 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3015) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u836 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3012), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3013), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3014), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3015), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3011) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u835 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2888) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u834 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2890) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u833 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2891) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u832 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2888), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2889), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2890), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2891), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2887) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u831 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2928) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u830 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2930) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u829 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2931) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u828 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2928), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2929), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2930), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2931), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2927) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u827 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2804) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u826 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2806) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u825 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2807) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u824 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2804), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2805), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2806), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2807), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2803) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u823 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2844) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u822 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2846) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u821 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2847) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u820 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2844), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2845), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2846), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2847), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2843) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u819 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2720) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u818 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2722) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u817 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2723) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u816 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2720), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2721), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2722), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2723), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2719) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u815 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2760) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u814 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2762) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u813 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2763) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u812 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2760), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2761), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2762), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2763), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2759) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u811 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2636) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u810 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2638) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u809 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2639) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u808 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2636), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2637), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2638), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2639), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2635) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u807 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2676) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u806 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2678) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u805 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2679) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u804 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2676), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2677), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2678), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2679), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2675) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u803 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n495) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u802 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n497) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u801 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n498) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u800 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n495), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n496), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n497), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n498), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n494) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u799 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n535) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u798 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n537) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u797 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n538) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u796 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n535), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n536), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n537), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n538), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n534) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u795 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n411) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u794 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n413) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u793 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n414) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u792 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n411), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n412), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n413), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n414), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n410) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u791 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n451) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u790 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n453) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u789 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n454) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u788 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n451), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n452), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n453), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n454), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n450) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u787 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3101) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u786 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3111) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u785 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3116) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u784 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3061) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u783 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3071) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u782 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3076) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u781 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3017) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u780 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3027) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u779 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3032) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u778 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2977) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u777 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2987) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u776 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2992) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u775 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2933) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u774 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2943) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u773 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2948) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u772 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2893) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u771 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2903) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u770 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2908) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u769 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2849) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u768 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2859) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u767 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2864) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u766 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2809) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u765 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2819) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u764 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2824) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u763 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2765) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u762 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2775) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u761 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2780) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u760 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2725) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u759 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2735) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u758 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2740) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u757 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2681) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u756 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2691) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u755 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2696) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u754 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2641) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u753 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2651) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u752 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2656) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u751 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n540) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u750 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n550) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u749 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n555) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u748 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n500) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u747 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n510) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u746 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n515) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u745 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n456) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u744 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n466) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u743 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n471) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u742 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n416) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u741 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n426) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u740 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n431) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u739 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3046) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u738 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3048) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u737 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3049) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u736 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3046), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3047), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3048), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3049), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3045) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u735 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3086) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u734 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3088) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u733 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3089) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u732 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3086), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3087), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3088), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3089), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3085) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u731 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3106) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u730 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3108) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u729 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3109) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u728 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3106), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3107), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3108), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3109), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3105) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u727 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3066) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u726 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3068) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u725 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3069) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u724 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3066), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3067), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3068), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3069), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3065) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u723 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2962) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u722 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2964) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u721 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2965) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u720 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2962), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2963), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2964), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2965), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2961) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u719 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3002) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u718 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3004) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u717 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3005) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u716 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3002), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3003), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3004), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3005), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3001) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u715 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3022) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u714 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3024) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u713 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3025) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u712 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3022), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3023), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3024), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3025), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3021) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u711 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2982) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u710 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2984) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u709 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2985) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u708 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2982), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2983), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2984), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2985), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2981) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u707 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2878) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u706 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2880) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u705 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2881) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u704 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2878), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2879), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2880), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2881), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2877) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u703 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2918) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u702 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2920) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u701 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2921) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u700 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2918), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2919), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2920), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2921), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2917) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u699 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2938) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u698 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2940) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u697 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2941) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u696 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2938), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2939), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2940), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2941), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2937) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u695 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2898) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u694 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2900) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u693 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2901) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u692 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2898), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2899), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2900), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2901), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2897) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u691 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2794) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u690 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2796) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u689 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2797) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u688 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2794), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2795), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2796), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2797), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2793) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u687 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2834) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u686 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2836) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u685 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2837) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u684 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2834), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2835), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2836), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2837), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2833) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u683 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2854) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u682 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2856) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u681 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2857) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u680 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2854), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2855), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2856), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2857), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2853) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u679 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2814) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u678 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2816) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u677 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2817) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u676 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2814), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2815), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2816), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2817), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2813) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u675 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2710) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u674 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2712) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u673 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2713) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u672 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2710), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2711), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2712), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2713), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2709) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u671 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2750) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u670 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2752) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u669 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2753) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u668 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2750), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2751), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2752), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2753), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2749) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u667 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2770) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u666 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2772) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u665 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2773) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u664 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2770), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2771), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2772), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2773), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2769) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u663 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2730) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u662 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2732) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u661 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2733) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u660 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2730), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2731), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2732), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2733), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2729) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u659 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2626) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u658 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2628) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u657 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2629) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u656 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2626), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2627), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2628), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2629), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n568) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u655 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2666) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u654 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2668) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u653 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2669) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u652 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2666), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2667), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2668), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2669), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2665) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u651 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2686) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u650 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2688) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u649 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2689) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u648 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2686), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2687), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2688), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2689), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2685) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u647 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2646) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u646 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2648) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u645 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2649) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u644 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2646), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2647), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2648), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2649), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2645) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u643 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n485) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u642 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n487) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u641 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n488) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u640 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n485), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n486), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n487), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n488), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n484) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u639 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n525) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u638 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n527) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u637 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n528) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u636 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n525), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n526), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n527), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n528), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n524) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u635 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n545) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u634 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n547) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u633 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n548) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u632 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n545), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n546), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n547), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n548), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n544) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u631 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n505) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u630 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n507) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u629 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n508) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u628 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n505), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n506), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n507), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n508), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n504) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u627 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n401) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u626 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n403) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u625 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n404) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u624 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n401), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n402), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n403), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n404), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n400) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u623 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n441) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u622 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n443) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u621 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n444) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u620 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n441), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n442), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n443), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n444), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n440) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u619 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n461) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u618 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n463) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u617 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n464) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u616 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n461), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n462), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n463), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n464), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n460) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u615 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n421) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u614 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n423) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u613 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n424) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u612 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n421), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n422), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n423), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n424), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n420) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u611 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3042) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u610 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3052) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u609 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3057) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u608 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3047) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u607 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3082) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u606 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3092) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u605 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3097) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u604 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3087) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u603 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3102) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u602 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3112) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u601 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3117) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u600 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3107) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u599 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3062) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u598 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3072) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u597 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3077) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u596 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__7_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__7_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__7_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__7_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3067) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u595 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2958) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u594 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2968) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u593 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2973) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u592 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2963) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u591 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2998) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u590 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3008) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u589 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3013) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u588 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3003) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u587 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3018) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u586 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3028) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u585 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3033) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u584 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3023) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u583 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2978) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u582 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2988) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u581 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2993) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u580 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__6_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__6_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__6_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__6_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2983) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u579 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2874) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u578 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2884) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u577 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2889) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u576 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2879) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u575 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2914) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u574 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2924) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u573 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2929) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u572 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2919) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u571 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2934) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u570 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2944) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u569 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2949) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u568 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2939) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u567 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2894) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u566 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2904) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u565 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2909) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u564 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__5_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__5_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__5_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__5_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2899) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u563 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2790) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u562 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2800) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u561 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2805) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u560 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2795) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u559 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2830) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u558 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2840) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u557 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2845) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u556 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2835) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u555 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2850) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u554 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2860) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u553 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2865) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u552 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2855) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u551 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2810) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u550 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2820) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u549 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2825) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u548 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__4_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__4_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__4_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__4_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2815) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u547 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2706) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u546 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2716) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u545 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2721) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u544 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2711) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u543 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2746) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u542 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2756) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u541 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2761) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u540 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2751) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u539 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2766) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u538 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2776) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u537 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2781) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u536 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2771) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u535 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2726) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u534 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2736) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u533 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2741) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u532 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__3_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__3_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__3_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__3_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2731) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u531 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n565) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u530 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2632) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u529 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2637) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u528 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2627) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u527 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2662) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u526 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2672) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u525 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2677) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u524 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2667) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u523 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2682) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u522 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2692) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u521 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2697) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u520 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2687) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u519 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2642) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u518 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2652) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u517 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2657) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u516 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__2_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__2_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__2_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__2_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2647) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u515 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n481) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u514 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n491) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u513 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n496) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u512 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n486) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u511 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n521) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u510 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n531) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u509 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n536) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u508 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n526) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u507 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n541) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u506 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n551) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u505 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n556) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u504 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n546) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u503 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n501) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u502 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n511) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u501 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n516) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u500 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__1_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__1_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__1_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__1_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n506) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u499 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n397) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u498 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n407) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u497 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n412) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u496 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n402) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u495 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n437) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u494 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n447) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u493 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n452) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u492 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n442) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u491 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n457) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u490 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n467) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u489 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n472) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u488 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n462) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u487 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n417) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u486 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n427) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u485 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n432) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u484 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__0_), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__0_), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__0_), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__0_), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n422) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u483 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3095), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3085), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3090), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3080), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3122) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u482 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3055), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3045), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3050), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3040), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3123) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u481 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3120), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3121), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3122), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3123), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3435) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u480 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3011), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3001), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3006), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2996), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3038) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u479 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2971), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2961), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2966), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2956), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3039) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u478 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3036), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3037), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3038), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3039), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3510) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u477 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2927), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2917), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2922), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2912), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2954) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u476 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2887), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2877), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2882), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2872), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2955) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u475 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2952), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2953), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2954), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2955), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3610) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u474 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2843), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2833), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2838), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2828), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2870) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u473 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2803), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2793), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2798), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2788), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2871) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u472 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2868), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2869), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2870), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2871), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3710) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u471 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2759), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2749), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2754), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2744), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2786) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u470 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2719), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2709), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2714), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2704), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2787) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u469 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2784), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2785), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2786), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2787), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3810) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u468 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2675), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2665), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2670), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2660), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2702) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u467 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2635), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n568), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2630), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n563), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2703) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u466 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2700), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2701), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2702), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2703), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3910) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u465 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n534), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n524), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n529), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n519), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n561) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u464 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n494), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n484), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n489), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n479), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n562) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u463 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n559), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n560), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n561), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n562), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4010) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u462 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n450), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n440), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n445), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n435), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n477) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u461 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n410), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n400), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n405), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n395), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n478) );
  MXIT4_X0P7M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u460 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n475), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n476), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n477), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n478), .S0(rd_addr[7]), .S1(
        oc8051_ram_top1_rd_addr_m_6_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4110) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u459 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3116), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3117), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3118), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3119), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3115) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u458 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3111), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3112), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3113), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3114), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3110) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u457 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3101), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3102), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3103), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3104), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3100) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u456 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3115), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3105), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3110), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3100), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3120) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u455 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3032), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3033), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3034), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3035), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3031) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u454 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3027), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3028), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3029), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3030), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3026) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u453 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3017), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3018), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3019), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3020), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3016) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u452 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3031), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3021), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3026), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3016), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3036) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u451 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2948), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2949), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2950), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2951), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2947) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u450 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2943), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2944), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2945), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2946), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2942) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u449 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2933), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2934), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2935), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2936), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2932) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u448 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2947), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2937), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2942), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2932), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2952) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u447 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2864), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2865), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2866), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2867), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2863) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u446 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2859), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2860), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2861), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2862), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2858) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u445 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2849), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2850), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2851), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2852), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2848) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u444 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2863), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2853), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2858), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2848), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2868) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u443 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2780), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2781), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2782), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2783), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2779) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u442 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2775), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2776), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2777), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2778), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2774) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u441 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2765), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2766), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2767), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2768), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2764) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u440 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2779), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2769), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2774), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2764), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2784) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u439 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2696), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2697), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2698), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2699), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2695) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u438 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2691), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2692), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2693), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2694), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2690) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u437 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2681), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2682), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2683), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2684), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2680) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u436 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2695), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2685), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2690), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2680), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2700) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u435 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n555), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n556), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n557), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n558), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n554) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u434 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n550), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n551), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n552), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n553), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n549) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u433 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n540), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n541), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n542), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n543), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n539) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u432 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n554), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n544), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n549), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n539), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n559) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u431 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n471), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n472), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n473), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n474), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n470) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u430 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n466), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n467), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n468), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n469), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n465) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u429 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n456), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n457), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n458), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n459), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n455) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u428 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n470), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n460), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n465), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n455), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n475) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u427 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3076), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3077), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3078), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3079), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3075) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u426 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3071), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3072), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3073), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3074), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3070) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u425 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3061), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3062), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3063), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3064), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3060) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u424 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3075), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3065), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3070), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3060), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3121) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u423 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2992), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2993), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2994), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2995), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2991) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u422 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2987), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2988), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2989), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2990), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2986) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u421 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2977), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2978), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2979), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2980), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2976) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u420 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2991), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2981), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2986), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2976), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3037) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u419 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2908), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2909), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2910), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2911), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2907) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u418 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2903), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2904), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2905), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2906), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2902) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u417 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2893), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2894), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2895), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2896), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2892) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u416 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2907), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2897), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2902), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2892), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2953) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u415 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2824), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2825), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2826), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2827), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2823) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u414 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2819), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2820), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2821), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2822), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2818) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u413 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2809), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2810), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2811), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2812), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2808) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u412 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2823), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2813), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2818), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2808), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2869) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u411 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2740), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2741), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2742), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2743), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2739) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u410 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2735), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2736), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2737), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2738), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2734) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u409 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2725), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2726), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2727), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2728), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2724) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u408 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2739), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2729), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2734), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2724), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2785) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u407 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2656), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2657), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2658), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2659), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2655) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u406 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2651), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2652), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2653), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2654), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2650) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u405 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2641), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2642), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2643), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2644), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2640) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u404 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2655), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2645), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2650), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2640), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2701) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u403 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n515), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n516), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n517), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n518), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n514) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u402 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n510), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n511), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n512), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n513), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n509) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u401 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n500), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n501), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n502), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n503), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n499) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u400 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n514), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n504), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n509), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n499), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n560) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u399 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n431), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n432), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n433), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n434), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n430) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u398 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n426), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n427), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n428), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n429), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n425) );
  MXIT4_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u397 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n416), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n417), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n418), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n419), .S0(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385), .S1(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n415) );
  MXIT4_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u396 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n430), .B(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n420), .C(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n425), .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n415), .S0(
        oc8051_ram_top1_rd_addr_m_5_), .S1(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n476) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u395 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n118) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u394 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n88)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u393 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n58)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u392 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n28)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u391 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n117) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u390 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n87)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u389 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n57)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u388 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n27)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u387 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n116) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u386 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n86)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u385 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n56)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u384 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n26)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u383 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n115) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u382 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n85)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u381 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n55)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u380 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n25)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u379 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n114) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u378 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n84)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u377 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n54)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u376 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n24)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u375 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n113) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u374 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n83)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u373 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n53)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u372 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n23)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u371 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n112) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u370 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n82)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u369 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n52)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u368 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n22)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u367 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n111) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u366 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n81)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u365 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n51)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u364 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n21)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u363 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n120) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u362 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n90)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u361 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n60)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u360 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n30)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u359 ( .A(
        oc8051_ram_top1_n10), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n119) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u358 ( .A(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n89)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u357 ( .A(
        oc8051_ram_top1_n7), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n59)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u356 ( .A(
        oc8051_ram_top1_n6), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n29)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u355 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n208) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u354 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n178) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u353 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n148) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u352 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n177) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u351 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n147) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u350 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n207) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u349 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n176) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u348 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n146) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u347 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n206) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u346 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n175) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u345 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n145) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u344 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n205) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u343 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n174) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u342 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n144) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u341 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n204) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u340 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n173) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u339 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n143) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u338 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n203) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u337 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n172) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u336 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n142) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u335 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n202) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u334 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n171) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u333 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n141) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u332 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n201) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u331 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n180) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u330 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n150) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u329 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n210) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u328 ( .A(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n179) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u327 ( .A(
        oc8051_ram_top1_n11), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n149) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u326 ( .A(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n209) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u325 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n238) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u324 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n237) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u323 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n236) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u322 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n235) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u321 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n234) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u320 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n233) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u319 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n232) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u318 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n231) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u317 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n240) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u316 ( .A(
        oc8051_ram_top1_n14), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n239) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u315 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n170) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u314 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n140) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u313 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n111), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n110) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u312 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n81), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n80) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u311 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n51), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n50) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u310 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n21), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n20) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u309 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n230) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u308 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n200) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u307 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n215) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u306 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n185) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u305 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n155) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u304 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n125) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u303 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n118), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n95) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u302 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n88), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n65) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u301 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n58), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n35) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u300 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n28), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n5) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u299 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n178), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n156) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u298 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n148), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n126) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u297 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n118), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n96) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u296 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n88), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n66) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u295 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n58), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n36) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u294 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n28), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n6) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u293 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n238), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n216) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u292 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n208), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n186) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u291 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n157) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u290 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n127) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u289 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n117), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n97) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u288 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n87), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n67) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u287 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n57), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n37) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u286 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n27), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n7) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u285 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n237), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n217) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u284 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n187) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u283 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n177), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n158) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u282 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n147), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n128) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u281 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n117), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n98) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u280 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n87), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n68) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u279 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n57), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n38) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u278 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n27), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n8) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u277 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n237), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n218) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u276 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n207), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n188) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u275 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n159) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u274 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n129) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u273 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n116), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n99) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u272 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n86), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n69) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u271 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n56), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n39) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u270 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n26), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n9) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u269 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n219) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u268 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n189) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u267 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n176), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n160) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u266 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n146), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n130) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u265 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n116), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n100) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u264 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n86), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n70) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u263 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n56), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n40) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u262 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n26), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n10) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u261 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n236), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n220) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u260 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n206), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n190) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u259 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n161) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u258 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n131) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u257 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n115), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n101) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u256 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n85), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n71) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u255 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n55), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n41) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u254 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n25), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n11) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u253 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n221) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u252 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n191) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u251 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n175), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n162) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u250 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n145), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n132) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u249 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n115), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n102) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u248 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n85), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n72) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u247 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n55), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n42) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u246 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n25), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n12) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u245 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n235), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n222) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u244 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n205), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n192) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u243 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n163) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u242 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n133) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u241 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n114), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n103) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u240 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n84), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n73) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u239 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n54), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n43) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u238 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n24), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n13) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u237 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n223) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u236 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n193) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u235 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n174), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n164) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u234 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n144), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n134) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u233 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n114), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n104) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u232 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n84), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n74) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u231 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n54), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n44) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u230 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n24), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n14) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u229 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n234), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n224) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u228 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n204), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n194) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u227 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n165) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u226 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n135) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u225 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n113), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n105) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u224 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n83), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n75) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u223 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n53), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n45) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u222 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n23), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n15) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u221 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n225) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u220 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n195) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u219 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n173), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n166) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u218 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n143), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n136) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u217 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n113), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n106) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u216 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n83), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n76) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u215 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n53), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n46) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u214 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n23), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n16) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u213 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n233), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n226) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u212 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n203), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n196) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u211 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n167) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u210 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n137) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u209 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n112), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n107) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u208 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n82), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n77) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u207 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n52), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n47) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u206 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n22), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n17) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u205 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n227) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u204 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n202), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n197) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u203 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n172), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n168) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u202 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n142), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n138) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u201 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n112), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n108) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u200 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n82), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n78) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u199 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n52), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n48) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u198 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n22), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n18) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u197 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n232), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n228) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u196 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n202), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n198) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u195 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n171), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n169) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u194 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n141), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n139) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u193 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n111), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n109) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u192 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n81), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n79) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u191 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n51), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n49) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u190 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n21), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n19) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u189 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n231), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n229) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u188 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n201), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n199) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u187 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n151) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u186 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n121) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u185 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n120), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n91) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u184 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n90), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n61) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u183 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n60), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n31) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u182 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n30), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u181 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n211) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u180 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n181) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u179 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n180), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n152) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u178 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n150), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n122) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u177 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n120), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n92) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u176 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n90), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n62) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u175 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n60), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n32) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u174 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n30), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u173 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n240), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n212) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u172 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n210), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n182) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u171 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n153) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u170 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n123) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u169 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n119), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n93) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u168 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n89), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n63) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u167 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n59), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n33) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u166 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n29), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n3) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u165 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n239), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n213) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u164 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n183) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u163 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n179), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n154) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u162 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n149), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n124) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u161 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n119), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n94) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u160 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n89), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n64) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u159 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n59), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n34) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u158 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n29), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n4) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u157 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n239), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n214) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u156 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n209), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n184) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u155 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n394)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u154 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n393)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u153 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n392)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u152 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n391)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u151 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n389)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u150 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n390)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u149 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n388)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u148 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n387)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u147 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n386)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u146 ( .A(
        oc8051_ram_top1_n2), .Y(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n385)
         );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u145 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n384) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u144 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n383) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u143 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n382) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u142 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n381) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u141 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n379) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u140 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n380) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u139 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n378) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u138 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n377) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u137 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n376) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u136 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n375) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u135 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n374) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u134 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n307) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u133 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n373) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u132 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n372) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u131 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n371) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u130 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n370) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u129 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n369) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u128 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n368) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u127 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n306) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u126 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n305) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u125 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n304) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u124 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n303) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u123 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n302) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u122 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n301) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u121 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n349) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u120 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n374), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n348) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u119 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n282) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u118 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n307), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n281) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u117 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n350) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u116 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n353) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u115 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n352) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u114 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n373), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n351) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u113 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n355) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u112 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n372), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n354) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u111 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n358) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u110 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n357) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u109 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n371), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n356) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u108 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n360) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u107 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n359) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u106 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n363) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u105 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n362) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u104 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n370), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n361) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u103 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n365) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u102 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n369), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n364) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u101 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n367) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u100 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n368), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n366) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u99 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n283) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u98 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n286) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u97 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n285) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u96 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n306), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n284) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u95 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n288) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u94 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n305), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n287) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u93 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n291) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u92 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n290) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u91 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n304), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n289) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u90 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n293) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u89 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n292) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u88 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n296) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u87 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n295) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u86 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n303), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n294) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u85 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n298) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u84 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n302), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n297) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u83 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n300) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u82 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n301), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n299) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u81 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n280) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u80 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n347) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u79 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n277) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u78 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n282), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n278) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u77 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n281), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n279) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u76 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n275) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u75 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n283), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n276) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u74 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n270) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u73 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n271) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u72 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n273) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u71 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n284), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n274) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u70 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n285), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n272) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u69 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n265) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u68 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n288), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n266) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u67 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n268) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u66 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n286), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n269) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u65 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n287), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n267) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u64 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n291), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n260) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u63 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n261) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u62 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n263) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u61 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n289), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n264) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u60 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n290), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n262) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u59 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n255) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u58 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n293), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n256) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u57 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n258) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u56 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n291), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n259) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u55 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n292), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n257) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u54 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n250) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u53 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n251) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u52 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n295), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n252) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u51 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n253) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u50 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n294), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n254) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u49 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n245) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u48 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n298), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n246) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u47 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n247) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u46 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n297), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n248) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u45 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n296), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n249) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u44 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n241) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u43 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n300), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n242) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u42 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n243) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u41 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n299), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n244) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u40 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n344) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u39 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n349), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n345) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u38 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n348), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n346) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u37 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n342) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u36 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n350), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n343) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u35 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n337) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u34 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n338) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u33 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n340) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u32 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n351), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n341) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u31 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n352), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n339) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u30 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n332) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u29 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n355), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n333) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u28 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n335) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u27 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n353), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n336) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u26 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n354), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n334) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u25 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n327) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u24 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n328) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u23 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n330) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u22 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n356), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n331) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u21 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n357), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n329) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u20 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n322) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u19 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n360), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n323) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u18 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n325) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u17 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n358), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n326) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u16 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n359), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n324) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u15 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n317) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u14 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n318) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u13 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n362), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n319) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u12 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n361), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n320) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u11 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n361), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n321) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u10 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n312) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u9 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n365), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n313) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u8 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n314) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u7 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n364), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n315) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u6 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n363), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n316) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u5 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n308) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u4 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n367), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n309) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u3 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n310) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_u2 ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n366), .Y(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n311) );
  BUFZ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_3_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_3_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[3]) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n570), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n571), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n572), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n573), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n574), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n575), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n576), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_reg_7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n577), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n594), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n595), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n596), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n597), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n598), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n599), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n600), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_2__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n601), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_2__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n626), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n627), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n628), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n629), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n630), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n631), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n632), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_6__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n633), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_6__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n658), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n659), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n660), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n661), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n662), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n663), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n664), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_10__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n665), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_10__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n690), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n691), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n692), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n693), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n694), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n695), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n696), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_14__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n697), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_14__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n722), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n723), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n724), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n725), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n726), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n727), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n728), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_18__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n729), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_18__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n754), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n755), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n756), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n757), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n758), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n759), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n760), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_22__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n761), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_22__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n786), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n787), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n788), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n789), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n790), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n791), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n792), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_26__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n793), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_26__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n818), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n819), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n820), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n821), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n822), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n823), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n824), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_30__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n825), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_30__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n850), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n851), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n852), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n853), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n854), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n855), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n856), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_34__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n857), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_34__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n882), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n883), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n884), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n885), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n886), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n887), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n888), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_38__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n889), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_38__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n914), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n915), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n916), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n917), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n918), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n919), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n920), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_42__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n921), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_42__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n946), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n947), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n948), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n949), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n950), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n951), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n952), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_46__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n953), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_46__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n978), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n979), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n980), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n981), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n982), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n983), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n984), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_50__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n985), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_50__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1010), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1011), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1012), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1013), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1014), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1015), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1016), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_54__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1017), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_54__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1042), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1043), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1044), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1045), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1046), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1047), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1048), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_58__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1049), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_58__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1074), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1075), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1076), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1077), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1078), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1079), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1080), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_62__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1081), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_62__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1106), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1107), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1108), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1109), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1110), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1111), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1112), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_66__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1113), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_66__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1138), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1139), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1140), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1141), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1142), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1143), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1144), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_70__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1145), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_70__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1170), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1171), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1172), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1173), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1174), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1175), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1176), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_74__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1177), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_74__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1202), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1203), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1204), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1205), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1206), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1207), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1208), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_78__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1209), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_78__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1234), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1235), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1236), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1237), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1238), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1239), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1240), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_82__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1241), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_82__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1266), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1267), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1268), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1269), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1270), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1271), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1272), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_86__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1273), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_86__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1298), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1299), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1300), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1301), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1302), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1303), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1304), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_90__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1305), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_90__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1330), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1331), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1332), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1333), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1334), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1335), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1336), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_94__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1337), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_94__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1362), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1363), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1364), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1365), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1366), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1367), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1368), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_98__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1369), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_98__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1394), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1395), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1396), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1397), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1398), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1399), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1400), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_102__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1401), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_102__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1426), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1427), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1428), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1429), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1430), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1431), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1432), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_106__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1433), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_106__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1458), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1459), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1460), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1461), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1462), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1463), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1464), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_110__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1465), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_110__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1490), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1491), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1492), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1493), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1494), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1495), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1496), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_114__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1497), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_114__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1522), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1523), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1524), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1525), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1526), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1527), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1528), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_118__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1529), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_118__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1554), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1555), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1556), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1557), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1558), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1559), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1560), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_122__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1561), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_122__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1586), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1587), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1588), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1589), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1590), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1591), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1592), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_126__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1593), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_126__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1618), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1619), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1620), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1621), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1622), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1623), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1624), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_130__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1625), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_130__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1650), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1651), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1652), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1653), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1654), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1655), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1656), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_134__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1657), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_134__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1682), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1683), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1684), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1685), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1686), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1687), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1688), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_138__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1689), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_138__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1714), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1715), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1716), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1717), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1718), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1719), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1720), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_142__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1721), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_142__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1746), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1747), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1748), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1749), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1750), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1751), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1752), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_146__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1753), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_146__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1778), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1779), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1780), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1781), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1782), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1783), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1784), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_150__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1785), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_150__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1810), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1811), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1812), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1813), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1814), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1815), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1816), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_154__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1817), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_154__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1842), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1843), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1844), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1845), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1846), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1847), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1848), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_158__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1849), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_158__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1874), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1875), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1876), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1877), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1878), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1879), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1880), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_162__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1881), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_162__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1906), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1907), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1908), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1909), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1910), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1911), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1912), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_166__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1913), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_166__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1938), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1939), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1940), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1941), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1942), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1943), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1944), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_170__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1945), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_170__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1970), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1971), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1972), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1973), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1974), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1975), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1976), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_174__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1977), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_174__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2002), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2003), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2004), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2005), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2006), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2007), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2008), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_178__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2009), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_178__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2034), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2035), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2036), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2037), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2038), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2039), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2040), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_182__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2041), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_182__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2066), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2067), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2068), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2069), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2070), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2071), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2072), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_186__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2073), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_186__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2098), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2099), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2100), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2101), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2102), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2103), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2104), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_190__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2105), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_190__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2130), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2131), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2132), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2133), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2134), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2135), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2136), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_194__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2137), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_194__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2162), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2163), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2164), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2165), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2166), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2167), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2168), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_198__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2169), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_198__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2194), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2195), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2196), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2197), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2198), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2199), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2200), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_202__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2201), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_202__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2226), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2227), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2228), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2229), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2230), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2231), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2232), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_206__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2233), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_206__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2258), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2259), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2260), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2261), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2262), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2263), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2264), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_210__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2265), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_210__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2290), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2291), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2292), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2293), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2294), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2295), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2296), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_214__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2297), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_214__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2322), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2323), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2324), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2325), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2326), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2327), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2328), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_218__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2329), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_218__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2354), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2355), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2356), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2357), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2358), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2359), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2360), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_222__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2361), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_222__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2386), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2387), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2388), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2389), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2390), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2391), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2392), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_226__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2393), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_226__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2418), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2419), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2420), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2421), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2422), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2423), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2424), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_230__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2425), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_230__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2450), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2451), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2452), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2453), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2454), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2455), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2456), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_234__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2457), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_234__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2482), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2483), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2484), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2485), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2486), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2487), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2488), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_238__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2489), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_238__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2514), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2515), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2516), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2517), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2518), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2519), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2520), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_242__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2521), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_242__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2546), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2547), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2548), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2549), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2550), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2551), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2552), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_246__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2553), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_246__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2578), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2579), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2580), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2581), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2582), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2583), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2584), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_250__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2585), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_250__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2610), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2611), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2612), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2613), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2614), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2615), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2616), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_254__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2617), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_254__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n578), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n579), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n580), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n581), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n582), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n583), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n584), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_0__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n585), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_0__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n610), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n611), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n612), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n613), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n614), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n615), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n616), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_4__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n617), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_4__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n642), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n643), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n644), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n645), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n646), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n647), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n648), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_8__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n649), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_8__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n674), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n675), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n676), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n677), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n678), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n679), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n680), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_12__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n681), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_12__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n706), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n707), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n708), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n709), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n710), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n711), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n712), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_16__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n713), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_16__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n738), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n739), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n740), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n741), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n742), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n743), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n744), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_20__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n745), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_20__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n770), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n771), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n772), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n773), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n774), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n775), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n776), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_24__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n777), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_24__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n802), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n803), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n804), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n805), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n806), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n807), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n808), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_28__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n809), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_28__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n834), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n835), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n836), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n837), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n838), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n839), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n840), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_32__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n841), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_32__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n866), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n867), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n868), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n869), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n870), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n871), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n872), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_36__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n873), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_36__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n898), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n899), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n900), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n901), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n902), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n903), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n904), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_40__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n905), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_40__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n930), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n931), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n932), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n933), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n934), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n935), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n936), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_44__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n937), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_44__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n962), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n963), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n964), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n965), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n966), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n967), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n968), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_48__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n969), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_48__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n994), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n995), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n996), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n997), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n998), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n999), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1000), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_52__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1001), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_52__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1026), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1027), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1028), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1029), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1030), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1031), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1032), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_56__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1033), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_56__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1058), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1059), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1060), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1061), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1062), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1063), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1064), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_60__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1065), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_60__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1090), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1091), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1092), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1093), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1094), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1095), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1096), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_64__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1097), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_64__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1122), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1123), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1124), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1125), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1126), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1127), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1128), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_68__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1129), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_68__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1154), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1155), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1156), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1157), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1158), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1159), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1160), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_72__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1161), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_72__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1186), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1187), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1188), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1189), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1190), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1191), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1192), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_76__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1193), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_76__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1218), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1219), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1220), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1221), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1222), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1223), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1224), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_80__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1225), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_80__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1250), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1251), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1252), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1253), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1254), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1255), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1256), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_84__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1257), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_84__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1282), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1283), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1284), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1285), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1286), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1287), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1288), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_88__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1289), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_88__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1314), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1315), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1316), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1317), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1318), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1319), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1320), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_92__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1321), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_92__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1346), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1347), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1348), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1349), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1350), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1351), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1352), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_96__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1353), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_96__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1378), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1379), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1380), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1381), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1382), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1383), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1384), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_100__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1385), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_100__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1410), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1411), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1412), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1413), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1414), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1415), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1416), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_104__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1417), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_104__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1442), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1443), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1444), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1445), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1446), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1447), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1448), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_108__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1449), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_108__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1474), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1475), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1476), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1477), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1478), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1479), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1480), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_112__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1481), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_112__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1506), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1507), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1508), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1509), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1510), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1511), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1512), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_116__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1513), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_116__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1538), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1539), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1540), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1541), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1542), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1543), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1544), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_120__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1545), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_120__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1570), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1571), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1572), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1573), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1574), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1575), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1576), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_124__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1577), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_124__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1602), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1603), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1604), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1605), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1606), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1607), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1608), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_128__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1609), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_128__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1634), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1635), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1636), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1637), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1638), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1639), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1640), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_132__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1641), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_132__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1666), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1667), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1668), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1669), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1670), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1671), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1672), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_136__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1673), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_136__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1698), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1699), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1700), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1701), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1702), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1703), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1704), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_140__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1705), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_140__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1730), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1731), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1732), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1733), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1734), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1735), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1736), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_144__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1737), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_144__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1762), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1763), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1764), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1765), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1766), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1767), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1768), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_148__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1769), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_148__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1794), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1795), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1796), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1797), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1798), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1799), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1800), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_152__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1801), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_152__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1826), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1827), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1828), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1829), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1830), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1831), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1832), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_156__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1833), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_156__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1858), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1859), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1860), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1861), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1862), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1863), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1864), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_160__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1865), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_160__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1890), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1891), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1892), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1893), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1894), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1895), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1896), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_164__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1897), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_164__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1922), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1923), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1924), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1925), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1926), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1927), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1928), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_168__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1929), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_168__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1954), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1955), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1956), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1957), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1958), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1959), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1960), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_172__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1961), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_172__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1986), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1987), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1988), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1989), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1990), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1991), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1992), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_176__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1993), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_176__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2018), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2019), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2020), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2021), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2022), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2023), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2024), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_180__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2025), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_180__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2050), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2051), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2052), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2053), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2054), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2055), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2056), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_184__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2057), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_184__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2082), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2083), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2084), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2085), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2086), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2087), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2088), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_188__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2089), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_188__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2114), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2115), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2116), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2117), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2118), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2119), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2120), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_192__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2121), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_192__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2146), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2147), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2148), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2149), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2150), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2151), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2152), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_196__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2153), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_196__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2178), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2179), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2180), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2181), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2182), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2183), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2184), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_200__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2185), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_200__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2210), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2211), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2212), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2213), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2214), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2215), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2216), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_204__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2217), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_204__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2242), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2243), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2244), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2245), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2246), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2247), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2248), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_208__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2249), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_208__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2274), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2275), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2276), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2277), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2278), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2279), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2280), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_212__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2281), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_212__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2306), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2307), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2308), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2309), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2310), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2311), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2312), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_216__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2313), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_216__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2338), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2339), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2340), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2341), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2342), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2343), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2344), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_220__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2345), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_220__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2370), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2371), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2372), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2373), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2374), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2375), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2376), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_224__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2377), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_224__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2402), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2403), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2404), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2405), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2406), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2407), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2408), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_228__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2409), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_228__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2434), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2435), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2436), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2437), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2438), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2439), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2440), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_232__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2441), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_232__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2466), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2467), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2468), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2469), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2470), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2471), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2472), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_236__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2473), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_236__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2498), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2499), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2500), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2501), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2502), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2503), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2504), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_240__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2505), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_240__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2530), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2531), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2532), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2533), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2534), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2535), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2536), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_244__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2537), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_244__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2562), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2563), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2564), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2565), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2566), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2567), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2568), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_248__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2569), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_248__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2594), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2595), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2596), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2597), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2598), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2599), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2600), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_252__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2601), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_252__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n586), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n587), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n588), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n589), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n590), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n591), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n592), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_1__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n593), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_1__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n618), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n619), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n620), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n621), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n622), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n623), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n624), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_5__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n625), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_5__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n650), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n651), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n652), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n653), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n654), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n655), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n656), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_9__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n657), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_9__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n682), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n683), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n684), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n685), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n686), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n687), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n688), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_13__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n689), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_13__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n714), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n715), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n716), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n717), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n718), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n719), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n720), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_17__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n721), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_17__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n746), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n747), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n748), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n749), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n750), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n751), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n752), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_21__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n753), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_21__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n778), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n779), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n780), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n781), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n782), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n783), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n784), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_25__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n785), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_25__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n810), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n811), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n812), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n813), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n814), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n815), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n816), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_29__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n817), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_29__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n842), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n843), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n844), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n845), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n846), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n847), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n848), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_33__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n849), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_33__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n874), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n875), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n876), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n877), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n878), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n879), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n880), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_37__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n881), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_37__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n906), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n907), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n908), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n909), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n910), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n911), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n912), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_41__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n913), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_41__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n938), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n939), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n940), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n941), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n942), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n943), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n944), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_45__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n945), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_45__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n970), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n971), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n972), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n973), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n974), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n975), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n976), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_49__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n977), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_49__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1002), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1003), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1004), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1005), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1006), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1007), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1008), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_53__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1009), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_53__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1034), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1035), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1036), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1037), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1038), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1039), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1040), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_57__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1041), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_57__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1066), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1067), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1068), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1069), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1070), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1071), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1072), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_61__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1073), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_61__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1098), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1099), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1100), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1101), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1102), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1103), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1104), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_65__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1105), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_65__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1130), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1131), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1132), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1133), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1134), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1135), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1136), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_69__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1137), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_69__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1162), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1163), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1164), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1165), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1166), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1167), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1168), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_73__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1169), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_73__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1194), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1195), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1196), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1197), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1198), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1199), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1200), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_77__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1201), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_77__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1226), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1227), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1228), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1229), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1230), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1231), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1232), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_81__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1233), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_81__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1258), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1259), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1260), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1261), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1262), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1263), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1264), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_85__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1265), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_85__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1290), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1291), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1292), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1293), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1294), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1295), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1296), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_89__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1297), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_89__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1322), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1323), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1324), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1325), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1326), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1327), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1328), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_93__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1329), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_93__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1354), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1355), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1356), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1357), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1358), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1359), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1360), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_97__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1361), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_97__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1386), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1387), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1388), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1389), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1390), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1391), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1392), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_101__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1393), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_101__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1418), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1419), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1420), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1421), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1422), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1423), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1424), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_105__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1425), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_105__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1450), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1451), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1452), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1453), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1454), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1455), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1456), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_109__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1457), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_109__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1482), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1483), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1484), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1485), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1486), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1487), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1488), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_113__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1489), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_113__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1514), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1515), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1516), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1517), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1518), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1519), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1520), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_117__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1521), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_117__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1546), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1547), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1548), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1549), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1550), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1551), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1552), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_121__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1553), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_121__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1578), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1579), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1580), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1581), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1582), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1583), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1584), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_125__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1585), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_125__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1610), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1611), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1612), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1613), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1614), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1615), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1616), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_129__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1617), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_129__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1642), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1643), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1644), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1645), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1646), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1647), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1648), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_133__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1649), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_133__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1674), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1675), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1676), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1677), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1678), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1679), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1680), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_137__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1681), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_137__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1706), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1707), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1708), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1709), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1710), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1711), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1712), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_141__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1713), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_141__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1738), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1739), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1740), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1741), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1742), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1743), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1744), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_145__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1745), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_145__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1770), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1771), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1772), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1773), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1774), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1775), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1776), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_149__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1777), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_149__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1802), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1803), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1804), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1805), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1806), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1807), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1808), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_153__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1809), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_153__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1834), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1835), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1836), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1837), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1838), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1839), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1840), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_157__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1841), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_157__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1866), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1867), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1868), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1869), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1870), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1871), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1872), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_161__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1873), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_161__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1898), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1899), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1900), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1901), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1902), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1903), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1904), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_165__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1905), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_165__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1930), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1931), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1932), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1933), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1934), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1935), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1936), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_169__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1937), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_169__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1962), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1963), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1964), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1965), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1966), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1967), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1968), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_173__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1969), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_173__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1994), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1995), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1996), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1997), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1998), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1999), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2000), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_177__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2001), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_177__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2026), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2027), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2028), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2029), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2030), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2031), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2032), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_181__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2033), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_181__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2058), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2059), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2060), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2061), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2062), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2063), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2064), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_185__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2065), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_185__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2090), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2091), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2092), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2093), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2094), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2095), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2096), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_189__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2097), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_189__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2122), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2123), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2124), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2125), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2126), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2127), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2128), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_193__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2129), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_193__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2154), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2155), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2156), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2157), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2158), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2159), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2160), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_197__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2161), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_197__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2186), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2187), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2188), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2189), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2190), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2191), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2192), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_201__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2193), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_201__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2218), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2219), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2220), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2221), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2222), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2223), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2224), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_205__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2225), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_205__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2250), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2251), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2252), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2253), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2254), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2255), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2256), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_209__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2257), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_209__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2282), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2283), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2284), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2285), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2286), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2287), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2288), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_213__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2289), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_213__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2314), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2315), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2316), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2317), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2318), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2319), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2320), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_217__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2321), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_217__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2346), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2347), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2348), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2349), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2350), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2351), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2352), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_221__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2353), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_221__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2378), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2379), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2380), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2381), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2382), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2383), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2384), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_225__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2385), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_225__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2410), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2411), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2412), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2413), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2414), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2415), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2416), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_229__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2417), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_229__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2442), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2443), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2444), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2445), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2446), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2447), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2448), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_233__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2449), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_233__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2474), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2475), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2476), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2477), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2478), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2479), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2480), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_237__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2481), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_237__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2506), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2507), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2508), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2509), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2510), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2511), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2512), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_241__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2513), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_241__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2538), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2539), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2540), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2541), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2542), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2543), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2544), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_245__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2545), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_245__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2570), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2571), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2572), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2573), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2574), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2575), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2576), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_249__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2577), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_249__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2602), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2603), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2604), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2605), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2606), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2607), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2608), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_253__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2609), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_253__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n602), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n603), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n604), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n605), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n606), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n607), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n608), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_3__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n609), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_3__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n634), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n635), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n636), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n637), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n638), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n639), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n640), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_7__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n641), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_7__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n666), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n667), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n668), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n669), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n670), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n671), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n672), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_11__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n673), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_11__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n698), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n699), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n700), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n701), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n702), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n703), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n704), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_15__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n705), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_15__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n730), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n731), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n732), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n733), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n734), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n735), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n736), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_19__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n737), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_19__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n762), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n763), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n764), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n765), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n766), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n767), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n768), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_23__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n769), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_23__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n794), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n795), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n796), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n797), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n798), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n799), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n800), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_27__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n801), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_27__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n826), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n827), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n828), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n829), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n830), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n831), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n832), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_31__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n833), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_31__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n858), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n859), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n860), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n861), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n862), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n863), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n864), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_35__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n865), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_35__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n890), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n891), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n892), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n893), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n894), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n895), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n896), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_39__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n897), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_39__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n922), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n923), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n924), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n925), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n926), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n927), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n928), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_43__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n929), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_43__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n954), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n955), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n956), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n957), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n958), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n959), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n960), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_47__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n961), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_47__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n986), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n987), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n988), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n989), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n990), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n991), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n992), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_51__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n993), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_51__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1018), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1019), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1020), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1021), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1022), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1023), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1024), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_55__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1025), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_55__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1050), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1051), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1052), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1053), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1054), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1055), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1056), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_59__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1057), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_59__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1082), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1083), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1084), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1085), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1086), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1087), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1088), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_63__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1089), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_63__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1114), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1115), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1116), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1117), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1118), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1119), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1120), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_67__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1121), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_67__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1146), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1147), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1148), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1149), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1150), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1151), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1152), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_71__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1153), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_71__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1178), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1179), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1180), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1181), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1182), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1183), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1184), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_75__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1185), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_75__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1210), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1211), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1212), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1213), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1214), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1215), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1216), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_79__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1217), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_79__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1242), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1243), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1244), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1245), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1246), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1247), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1248), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_83__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1249), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_83__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1274), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1275), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1276), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1277), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1278), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1279), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1280), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_87__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1281), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_87__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1306), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1307), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1308), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1309), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1310), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1311), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1312), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_91__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1313), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_91__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1338), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1339), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1340), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1341), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1342), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1343), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1344), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_95__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1345), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_95__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1370), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1371), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1372), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1373), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1374), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1375), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1376), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_99__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1377), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_99__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1402), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1403), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1404), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1405), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1406), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1407), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1408), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_103__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1409), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_103__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1434), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1435), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1436), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1437), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1438), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1439), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1440), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_107__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1441), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_107__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1466), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1467), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1468), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1469), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1470), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1471), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1472), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_111__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1473), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_111__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1498), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1499), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1500), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1501), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1502), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1503), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1504), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_115__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1505), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_115__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1530), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1531), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1532), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1533), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1534), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1535), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1536), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_119__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1537), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_119__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1562), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1563), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1564), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1565), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1566), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1567), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1568), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_123__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1569), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_123__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1594), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1595), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1596), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1597), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1598), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1599), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1600), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_127__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1601), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_127__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1626), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1627), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1628), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1629), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1630), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1631), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1632), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_131__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1633), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_131__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1658), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1659), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1660), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1661), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1662), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1663), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1664), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_135__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1665), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_135__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1690), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1691), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1692), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1693), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1694), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1695), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1696), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_139__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1697), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_139__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1722), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1723), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1724), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1725), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1726), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1727), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1728), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_143__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1729), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_143__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1754), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1755), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1756), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1757), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1758), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1759), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1760), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_147__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1761), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_147__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1786), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1787), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1788), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1789), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1790), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1791), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1792), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_151__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1793), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_151__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1818), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1819), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1820), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1821), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1822), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1823), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1824), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_155__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1825), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_155__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1850), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1851), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1852), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1853), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1854), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1855), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1856), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_159__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1857), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_159__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1882), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1883), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1884), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1885), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1886), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1887), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1888), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_163__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1889), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_163__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1914), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1915), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1916), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1917), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1918), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1919), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1920), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_167__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1921), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_167__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1946), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1947), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1948), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1949), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1950), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1951), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1952), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_171__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1953), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_171__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1978), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1979), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1980), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1981), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1982), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1983), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1984), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_175__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n1985), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_175__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2010), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2011), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2012), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2013), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2014), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2015), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2016), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_179__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2017), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_179__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2042), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2043), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2044), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2045), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2046), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2047), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2048), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_183__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2049), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_183__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2074), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2075), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2076), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2077), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2078), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2079), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2080), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_187__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2081), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_187__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2106), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2107), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2108), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2109), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2110), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2111), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2112), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_191__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2113), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_191__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2138), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2139), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2140), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2141), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2142), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2143), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2144), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_195__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2145), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_195__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2170), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2171), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2172), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2173), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2174), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2175), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2176), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_199__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2177), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_199__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2202), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2203), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2204), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2205), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2206), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2207), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2208), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_203__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2209), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_203__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2234), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2235), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2236), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2237), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2238), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2239), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2240), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_207__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2241), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_207__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2266), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2267), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2268), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2269), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2270), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2271), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2272), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_211__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2273), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_211__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2298), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2299), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2300), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2301), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2302), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2303), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2304), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_215__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2305), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_215__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2330), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2331), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2332), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2333), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2334), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2335), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2336), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_219__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2337), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_219__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2362), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2363), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2364), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2365), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2366), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2367), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2368), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_223__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2369), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_223__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2394), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2395), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2396), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2397), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2398), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2399), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2400), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_227__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2401), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_227__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2426), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2427), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2428), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2429), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2430), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2431), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2432), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_231__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2433), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_231__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2458), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2459), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2460), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2461), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2462), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2463), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2464), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_235__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2465), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_235__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2490), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2491), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2492), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2493), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2494), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2495), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2496), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_239__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2497), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_239__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2522), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2523), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2524), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2525), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2526), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2527), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2528), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_243__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2529), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_243__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2554), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2555), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2556), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2557), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2558), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2559), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2560), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_247__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2561), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_247__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2586), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2587), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2588), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2589), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2590), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2591), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2592), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_251__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2593), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_251__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__0_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2618), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__1_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2619), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__2_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2620), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__3_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2621), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__4_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2622), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__5_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2623), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__6_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2624), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_reg_255__7_ ( 
        .D(oc8051_ram_top1_oc8051_idata_oc8051_ram1_n2625), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_mem_255__7_) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_7_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_7_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[7]) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_6_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_6_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[6]) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_5_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_5_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[5]) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_4_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_4_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[4]) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_2_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_2_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[2]) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_1_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_1_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[1]) );
  BUFZ_X6M_A12TS oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_tri_0_ ( .A(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_do_reg_0_), .OE(
        oc8051_ram_top1_oc8051_idata_oc8051_ram1_n569), .Y(
        oc8051_ram_top1_rd_data_m[0]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u87 ( .A(ram_out[3]), .Y(
        oc8051_alu_src_sel1_n25) );
  OR2_X0P5M_A12TS oc8051_alu_src_sel1_u86 ( .A(src_sel2[0]), .B(src_sel2[1]), 
        .Y(oc8051_alu_src_sel1_n29) );
  NAND2_X0P5A_A12TS oc8051_alu_src_sel1_u85 ( .A(src_sel2[1]), .B(src_sel2[0]), 
        .Y(oc8051_alu_src_sel1_n30) );
  NAND2B_X0P5M_A12TS oc8051_alu_src_sel1_u84 ( .AN(src_sel2[1]), .B(
        src_sel2[0]), .Y(oc8051_alu_src_sel1_n31) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u83 ( .A(oc8051_alu_src_sel1_op2_r_3_), 
        .Y(oc8051_alu_src_sel1_n61) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u82 ( .A(acc[3]), .Y(
        oc8051_alu_src_sel1_n60) );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u81 ( .A(src_sel1[1]), .B(src_sel1[2]), 
        .C(src_sel1[0]), .Y(oc8051_alu_src_sel1_n34) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u80 ( .A(src_sel1[2]), .Y(
        oc8051_alu_src_sel1_n58) );
  NOR2_X0P5A_A12TS oc8051_alu_src_sel1_u79 ( .A(oc8051_alu_src_sel1_n58), .B(
        src_sel1[0]), .Y(oc8051_alu_src_sel1_n35) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u78 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[0]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[8]), .Y(
        oc8051_alu_src_sel1_n54) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u77 ( .A(src_sel1[0]), .Y(
        oc8051_alu_src_sel1_n57) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u76 ( .A(src_sel1[1]), .Y(
        oc8051_alu_src_sel1_n59) );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u75 ( .A(oc8051_alu_src_sel1_n57), .B(
        src_sel1[2]), .C(oc8051_alu_src_sel1_n59), .Y(oc8051_alu_src_sel1_n32)
         );
  NOR2_X0P5A_A12TS oc8051_alu_src_sel1_u74 ( .A(oc8051_alu_src_sel1_n58), .B(
        oc8051_alu_src_sel1_n59), .Y(oc8051_alu_src_sel1_n33) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u73 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[0]), .B0(oc8051_alu_src_sel1_op1_r[0]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n55) );
  NOR2_X0P5A_A12TS oc8051_alu_src_sel1_u72 ( .A(oc8051_alu_src_sel1_n59), .B(
        src_sel1[0]), .Y(oc8051_alu_src_sel1_n26) );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u71 ( .A(oc8051_alu_src_sel1_n57), .B(
        src_sel1[1]), .C(oc8051_alu_src_sel1_n58), .Y(oc8051_alu_src_sel1_n27)
         );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u70 ( .A(src_sel1[1]), .B(src_sel1[2]), 
        .C(oc8051_alu_src_sel1_n57), .Y(oc8051_alu_src_sel1_n28) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u69 ( .A0(
        oc8051_alu_src_sel1_op3_r[0]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[0]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_0_), .Y(oc8051_alu_src_sel1_n56) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u68 ( .A(oc8051_alu_src_sel1_n54), .B(
        oc8051_alu_src_sel1_n55), .C(oc8051_alu_src_sel1_n56), .Y(src1[0]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u67 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[1]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[9]), .Y(
        oc8051_alu_src_sel1_n51) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u66 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[1]), .B0(oc8051_alu_src_sel1_op1_r[1]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n52) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u65 ( .A0(
        oc8051_alu_src_sel1_op3_r[1]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[1]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_1_), .Y(oc8051_alu_src_sel1_n53) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u64 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[2]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[10]), .Y(
        oc8051_alu_src_sel1_n48) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u63 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[2]), .B0(oc8051_alu_src_sel1_op1_r[2]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n49) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u62 ( .A0(
        oc8051_alu_src_sel1_op3_r[2]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[2]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_2_), .Y(oc8051_alu_src_sel1_n50) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u61 ( .A(oc8051_alu_src_sel1_n48), .B(
        oc8051_alu_src_sel1_n49), .C(oc8051_alu_src_sel1_n50), .Y(src1[2]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u60 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[3]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[11]), .Y(
        oc8051_alu_src_sel1_n45) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u59 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[3]), .B0(oc8051_alu_src_sel1_op1_r[3]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n46) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u58 ( .A0(
        oc8051_alu_src_sel1_op3_r[3]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[3]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_3_), .Y(oc8051_alu_src_sel1_n47) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u57 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[4]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[12]), .Y(
        oc8051_alu_src_sel1_n42) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u56 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[4]), .B0(oc8051_alu_src_sel1_op1_r[4]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n43) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u55 ( .A0(
        oc8051_alu_src_sel1_op3_r[4]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[4]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_4_), .Y(oc8051_alu_src_sel1_n44) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u54 ( .A(oc8051_alu_src_sel1_n42), .B(
        oc8051_alu_src_sel1_n43), .C(oc8051_alu_src_sel1_n44), .Y(src1[4]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u53 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[5]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[13]), .Y(
        oc8051_alu_src_sel1_n39) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u52 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[5]), .B0(oc8051_alu_src_sel1_op1_r[5]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n40) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u51 ( .A0(
        oc8051_alu_src_sel1_op3_r[5]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[5]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_5_), .Y(oc8051_alu_src_sel1_n41) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u50 ( .A(oc8051_alu_src_sel1_n39), .B(
        oc8051_alu_src_sel1_n40), .C(oc8051_alu_src_sel1_n41), .Y(src1[5]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u49 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[6]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[14]), .Y(
        oc8051_alu_src_sel1_n36) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u48 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[6]), .B0(oc8051_alu_src_sel1_op1_r[6]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n37) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u47 ( .A0(
        oc8051_alu_src_sel1_op3_r[6]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[6]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_6_), .Y(oc8051_alu_src_sel1_n38) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u46 ( .A(oc8051_alu_src_sel1_n36), .B(
        oc8051_alu_src_sel1_n37), .C(oc8051_alu_src_sel1_n38), .Y(src1[6]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u45 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(ram_out[7]), .B0(oc8051_alu_src_sel1_n35), .B1(pc[15]), .Y(
        oc8051_alu_src_sel1_n22) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u44 ( .A0(oc8051_alu_src_sel1_n32), 
        .A1(acc[7]), .B0(oc8051_alu_src_sel1_op1_r[7]), .B1(
        oc8051_alu_src_sel1_n33), .Y(oc8051_alu_src_sel1_n23) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u43 ( .A0(
        oc8051_alu_src_sel1_op3_r[7]), .A1(oc8051_alu_src_sel1_n26), .B0(pc[7]), .B1(oc8051_alu_src_sel1_n27), .C0(oc8051_alu_src_sel1_n28), .C1(
        oc8051_alu_src_sel1_op2_r_7_), .Y(oc8051_alu_src_sel1_n24) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u42 ( .A(oc8051_alu_src_sel1_n22), .B(
        oc8051_alu_src_sel1_n23), .C(oc8051_alu_src_sel1_n24), .Y(src1[7]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u41 ( .A(oc8051_alu_src_sel1_op2_r_0_), 
        .Y(oc8051_alu_src_sel1_n19) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u40 ( .A(ram_out[0]), .Y(
        oc8051_alu_src_sel1_n20) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u39 ( .A(acc[0]), .Y(
        oc8051_alu_src_sel1_n21) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u38 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n19), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n20), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n21), .Y(src2[0]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u37 ( .A(oc8051_alu_src_sel1_op2_r_1_), 
        .Y(oc8051_alu_src_sel1_n16) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u36 ( .A(ram_out[1]), .Y(
        oc8051_alu_src_sel1_n17) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u35 ( .A(acc[1]), .Y(
        oc8051_alu_src_sel1_n18) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u34 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n16), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n17), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n18), .Y(src2[1]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u33 ( .A(oc8051_alu_src_sel1_op2_r_2_), 
        .Y(oc8051_alu_src_sel1_n13) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u32 ( .A(ram_out[2]), .Y(
        oc8051_alu_src_sel1_n14) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u31 ( .A(acc[2]), .Y(
        oc8051_alu_src_sel1_n15) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u30 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n13), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n14), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n15), .Y(src2[2]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u29 ( .A(oc8051_alu_src_sel1_op2_r_4_), 
        .Y(oc8051_alu_src_sel1_n10) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u28 ( .A(ram_out[4]), .Y(
        oc8051_alu_src_sel1_n11) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u27 ( .A(acc[4]), .Y(
        oc8051_alu_src_sel1_n12) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u26 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n10), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n11), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n12), .Y(src2[4]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u25 ( .A(oc8051_alu_src_sel1_op2_r_5_), 
        .Y(oc8051_alu_src_sel1_n7) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u24 ( .A(ram_out[5]), .Y(
        oc8051_alu_src_sel1_n8) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u23 ( .A(acc[5]), .Y(
        oc8051_alu_src_sel1_n9) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u22 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n7), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n8), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n9), .Y(src2[5]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u21 ( .A(oc8051_alu_src_sel1_op2_r_6_), 
        .Y(oc8051_alu_src_sel1_n4) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u20 ( .A(ram_out[6]), .Y(
        oc8051_alu_src_sel1_n5) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u19 ( .A(acc[6]), .Y(
        oc8051_alu_src_sel1_n6) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u18 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n4), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n5), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n6), .Y(src2[6]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u17 ( .A(oc8051_alu_src_sel1_op2_r_7_), 
        .Y(oc8051_alu_src_sel1_n1) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u16 ( .A(ram_out[7]), .Y(
        oc8051_alu_src_sel1_n2) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u14 ( .A(acc[7]), .Y(
        oc8051_alu_src_sel1_n3) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u13 ( .A0(oc8051_alu_src_sel1_n30), 
        .A1(oc8051_alu_src_sel1_n1), .B0(oc8051_alu_src_sel1_n29), .B1(
        oc8051_alu_src_sel1_n2), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n3), .Y(src2[7]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u12 ( .A(dptr_hi[0]), .B(pc[8]), .S0(
        src_sel3), .Y(src3[0]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u11 ( .A(dptr_hi[1]), .B(pc[9]), .S0(
        src_sel3), .Y(src3[1]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u10 ( .A(dptr_hi[2]), .B(pc[10]), .S0(
        src_sel3), .Y(src3[2]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u9 ( .A(dptr_hi[3]), .B(pc[11]), .S0(
        src_sel3), .Y(src3[3]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u8 ( .A(dptr_hi[4]), .B(pc[12]), .S0(
        src_sel3), .Y(src3[4]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u7 ( .A(dptr_hi[5]), .B(pc[13]), .S0(
        src_sel3), .Y(src3[5]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u6 ( .A(dptr_hi[6]), .B(pc[14]), .S0(
        src_sel3), .Y(src3[6]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u5 ( .A(dptr_hi[7]), .B(pc[15]), .S0(
        src_sel3), .Y(src3[7]) );
  NAND3_X1M_A12TS oc8051_alu_src_sel1_u4 ( .A(oc8051_alu_src_sel1_n45), .B(
        oc8051_alu_src_sel1_n46), .C(oc8051_alu_src_sel1_n47), .Y(src1[3]) );
  NAND3_X1M_A12TS oc8051_alu_src_sel1_u3 ( .A(oc8051_alu_src_sel1_n51), .B(
        oc8051_alu_src_sel1_n52), .C(oc8051_alu_src_sel1_n53), .Y(src1[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_0_ ( .D(op2_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_1_ ( .D(op2_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_1_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_2_ ( .D(op2_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_2_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_3_ ( .D(op2_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_3_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_4_ ( .D(op2_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_4_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_5_ ( .D(op2_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_5_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_6_ ( .D(op2_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_6_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_7_ ( .D(op2_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_7_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_0_ ( .D(op1_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_1_ ( .D(op1_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_2_ ( .D(op1_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_3_ ( .D(op1_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_4_ ( .D(op1_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_5_ ( .D(op1_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_6_ ( .D(op1_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_7_ ( .D(op1_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_0_ ( .D(op3_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_1_ ( .D(op3_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_2_ ( .D(op3_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_3_ ( .D(op3_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_4_ ( .D(op3_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_5_ ( .D(op3_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_6_ ( .D(op3_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_7_ ( .D(op3_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[7]) );
  OAI222_X4M_A12TS oc8051_alu_src_sel1_u15 ( .A0(oc8051_alu_src_sel1_n29), 
        .A1(oc8051_alu_src_sel1_n25), .B0(oc8051_alu_src_sel1_n30), .B1(
        oc8051_alu_src_sel1_n61), .C0(oc8051_alu_src_sel1_n31), .C1(
        oc8051_alu_src_sel1_n60), .Y(src2[3]) );
  NOR2_X0P5A_A12TS oc8051_comp1_u11 ( .A(acc[1]), .B(acc[0]), .Y(
        oc8051_comp1_n7) );
  NOR2_X0P5A_A12TS oc8051_comp1_u10 ( .A(acc[3]), .B(acc[2]), .Y(
        oc8051_comp1_n8) );
  NOR2_X0P5A_A12TS oc8051_comp1_u9 ( .A(acc[5]), .B(acc[4]), .Y(
        oc8051_comp1_n9) );
  NOR2_X0P5A_A12TS oc8051_comp1_u8 ( .A(acc[7]), .B(acc[6]), .Y(
        oc8051_comp1_n10) );
  AND4_X0P5M_A12TS oc8051_comp1_u7 ( .A(oc8051_comp1_n7), .B(oc8051_comp1_n8), 
        .C(oc8051_comp1_n9), .D(oc8051_comp1_n10), .Y(oc8051_comp1_n1) );
  NOR2_X0P5A_A12TS oc8051_comp1_u6 ( .A(sub_result[1]), .B(sub_result[0]), .Y(
        oc8051_comp1_n3) );
  NOR2_X0P5A_A12TS oc8051_comp1_u5 ( .A(sub_result[3]), .B(sub_result[2]), .Y(
        oc8051_comp1_n4) );
  NOR2_X0P5A_A12TS oc8051_comp1_u4 ( .A(sub_result[5]), .B(sub_result[4]), .Y(
        oc8051_comp1_n5) );
  NOR2_X0P5A_A12TS oc8051_comp1_u3 ( .A(sub_result[7]), .B(sub_result[6]), .Y(
        oc8051_comp1_n6) );
  AND4_X0P5M_A12TS oc8051_comp1_u2 ( .A(oc8051_comp1_n3), .B(oc8051_comp1_n4), 
        .C(oc8051_comp1_n5), .D(oc8051_comp1_n6), .Y(oc8051_comp1_n2) );
  MXT4_X0P5M_A12TS oc8051_comp1_u1 ( .A(oc8051_comp1_n1), .B(cy), .C(
        oc8051_comp1_n2), .D(bit_out), .S0(comp_sel[1]), .S1(comp_sel[0]), .Y(
        eq) );
  OAI21_X0P5M_A12TS oc8051_cy_select1_u4 ( .A0(cy_sel[0]), .A1(bit_out), .B0(
        cy_sel[1]), .Y(oc8051_cy_select1_n1) );
  AO1B2_X0P5M_A12TS oc8051_cy_select1_u3 ( .B0(cy_sel[0]), .B1(cy), .A0N(
        oc8051_cy_select1_n1), .Y(alu_cy) );
  INV_X0P5B_A12TS oc8051_indi_addr1_u116 ( .A(wr_addr[0]), .Y(
        oc8051_indi_addr1_n26) );
  INV_X0P5B_A12TS oc8051_indi_addr1_u115 ( .A(wr_addr[3]), .Y(
        oc8051_indi_addr1_n92) );
  NOR2B_X0P5M_A12TS oc8051_indi_addr1_u114 ( .AN(wr_o), .B(
        oc8051_indi_addr1_wr_bit_r), .Y(oc8051_indi_addr1_n22) );
  NOR2B_X0P5M_A12TS oc8051_indi_addr1_u113 ( .AN(oc8051_indi_addr1_n22), .B(
        wr_addr[4]), .Y(oc8051_indi_addr1_n95) );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u112 ( .A(oc8051_indi_addr1_n26), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n95), .Y(
        oc8051_indi_addr1_n98) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u111 ( .A(oc8051_indi_addr1_buff_0__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n28)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u110 ( .A(oc8051_indi_addr1_buff_0__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n29)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u109 ( .A(oc8051_indi_addr1_buff_0__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n30)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u108 ( .A(oc8051_indi_addr1_buff_0__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n31)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u107 ( .A(oc8051_indi_addr1_buff_0__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n32)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u106 ( .A(oc8051_indi_addr1_buff_0__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n33)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u105 ( .A(oc8051_indi_addr1_buff_0__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n34)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u104 ( .A(oc8051_indi_addr1_buff_0__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n35)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u103 ( .A(wr_addr[0]), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n95), .Y(
        oc8051_indi_addr1_n97) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u102 ( .A(oc8051_indi_addr1_buff_1__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n36)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u101 ( .A(oc8051_indi_addr1_buff_1__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n37)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u100 ( .A(oc8051_indi_addr1_buff_1__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n38)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u99 ( .A(oc8051_indi_addr1_buff_1__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n39)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u98 ( .A(oc8051_indi_addr1_buff_1__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n40)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u97 ( .A(oc8051_indi_addr1_buff_1__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n41)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u96 ( .A(oc8051_indi_addr1_buff_1__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n42)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u95 ( .A(oc8051_indi_addr1_buff_1__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n43)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u94 ( .A(wr_addr[3]), .B(
        oc8051_indi_addr1_n26), .C(oc8051_indi_addr1_n95), .Y(
        oc8051_indi_addr1_n96) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u93 ( .A(oc8051_indi_addr1_buff_2__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n44)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u92 ( .A(oc8051_indi_addr1_buff_2__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n45)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u91 ( .A(oc8051_indi_addr1_buff_2__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n46)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u90 ( .A(oc8051_indi_addr1_buff_2__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n47)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u89 ( .A(oc8051_indi_addr1_buff_2__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n48)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u88 ( .A(oc8051_indi_addr1_buff_2__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n49)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u87 ( .A(oc8051_indi_addr1_buff_2__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n50)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u86 ( .A(oc8051_indi_addr1_buff_2__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n51)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u85 ( .A(wr_addr[3]), .B(wr_addr[0]), .C(
        oc8051_indi_addr1_n95), .Y(oc8051_indi_addr1_n94) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u84 ( .A(oc8051_indi_addr1_buff_3__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n52)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u83 ( .A(oc8051_indi_addr1_buff_3__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n53)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u82 ( .A(oc8051_indi_addr1_buff_3__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n54)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u81 ( .A(oc8051_indi_addr1_buff_3__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n55)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u80 ( .A(oc8051_indi_addr1_buff_3__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n56)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u79 ( .A(oc8051_indi_addr1_buff_3__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n57)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u78 ( .A(oc8051_indi_addr1_buff_3__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n58)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u77 ( .A(oc8051_indi_addr1_buff_3__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n59)
         );
  AND2_X0P5M_A12TS oc8051_indi_addr1_u76 ( .A(oc8051_indi_addr1_n22), .B(
        wr_addr[4]), .Y(oc8051_indi_addr1_n24) );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u75 ( .A(oc8051_indi_addr1_n26), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n24), .Y(
        oc8051_indi_addr1_n93) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u74 ( .A(oc8051_indi_addr1_buff_4__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n60)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u73 ( .A(oc8051_indi_addr1_buff_4__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n61)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u72 ( .A(oc8051_indi_addr1_buff_4__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n62)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u71 ( .A(oc8051_indi_addr1_buff_4__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n63)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u70 ( .A(oc8051_indi_addr1_buff_4__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n64)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u69 ( .A(oc8051_indi_addr1_buff_4__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n65)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u68 ( .A(oc8051_indi_addr1_buff_4__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n66)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u67 ( .A(oc8051_indi_addr1_buff_4__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n67)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u66 ( .A(wr_addr[0]), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n24), .Y(
        oc8051_indi_addr1_n27) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u65 ( .A(oc8051_indi_addr1_buff_5__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n68)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u64 ( .A(oc8051_indi_addr1_buff_5__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n69)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u63 ( .A(oc8051_indi_addr1_buff_5__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n70)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u62 ( .A(oc8051_indi_addr1_buff_5__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n71)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u61 ( .A(oc8051_indi_addr1_buff_5__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n72)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u60 ( .A(oc8051_indi_addr1_buff_5__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n73)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u59 ( .A(oc8051_indi_addr1_buff_5__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n74)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u58 ( .A(oc8051_indi_addr1_buff_5__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n75)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u57 ( .A(wr_addr[3]), .B(
        oc8051_indi_addr1_n26), .C(oc8051_indi_addr1_n24), .Y(
        oc8051_indi_addr1_n25) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u56 ( .A(oc8051_indi_addr1_buff_6__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n76)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u55 ( .A(oc8051_indi_addr1_buff_6__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n77)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u54 ( .A(oc8051_indi_addr1_buff_6__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n78)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u53 ( .A(oc8051_indi_addr1_buff_6__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n79)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u52 ( .A(oc8051_indi_addr1_buff_6__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n80)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u51 ( .A(oc8051_indi_addr1_buff_6__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n81)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u50 ( .A(oc8051_indi_addr1_buff_6__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n82)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u49 ( .A(oc8051_indi_addr1_buff_6__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n83)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u48 ( .A(wr_addr[3]), .B(wr_addr[0]), .C(
        oc8051_indi_addr1_n24), .Y(oc8051_indi_addr1_n23) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u47 ( .A(oc8051_indi_addr1_buff_7__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n84)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u46 ( .A(oc8051_indi_addr1_buff_7__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n85)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u45 ( .A(oc8051_indi_addr1_buff_7__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n86)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u44 ( .A(oc8051_indi_addr1_buff_7__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n87)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u43 ( .A(oc8051_indi_addr1_buff_7__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n88)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u42 ( .A(oc8051_indi_addr1_buff_7__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n89)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u41 ( .A(oc8051_indi_addr1_buff_7__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n90)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u40 ( .A(oc8051_indi_addr1_buff_7__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n91)
         );
  XNOR2_X0P5M_A12TS oc8051_indi_addr1_u39 ( .A(wr_addr[4]), .B(bank_sel[1]), 
        .Y(oc8051_indi_addr1_n19) );
  XNOR2_X0P5M_A12TS oc8051_indi_addr1_u38 ( .A(wr_addr[3]), .B(bank_sel[0]), 
        .Y(oc8051_indi_addr1_n20) );
  XNOR2_X0P5M_A12TS oc8051_indi_addr1_u37 ( .A(wr_addr[0]), .B(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n21) );
  NAND4_X0P5A_A12TS oc8051_indi_addr1_u36 ( .A(oc8051_indi_addr1_n19), .B(
        oc8051_indi_addr1_n20), .C(oc8051_indi_addr1_n21), .D(
        oc8051_indi_addr1_n22), .Y(oc8051_indi_addr1_n18) );
  OR6_X0P5M_A12TS oc8051_indi_addr1_u35 ( .A(wr_addr[7]), .B(wr_addr[6]), .C(
        wr_addr[5]), .D(wr_addr[2]), .E(wr_addr[1]), .F(oc8051_indi_addr1_n18), 
        .Y(oc8051_indi_addr1_n17) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u34 ( .A(wr_dat[0]), .B(
        oc8051_indi_addr1_n106), .S0(oc8051_indi_addr1_n17), .Y(ri[0]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u33 ( .A(wr_dat[1]), .B(
        oc8051_indi_addr1_n105), .S0(oc8051_indi_addr1_n17), .Y(ri[1]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u32 ( .A(wr_dat[2]), .B(
        oc8051_indi_addr1_n104), .S0(oc8051_indi_addr1_n17), .Y(ri[2]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u31 ( .A(wr_dat[3]), .B(
        oc8051_indi_addr1_n103), .S0(oc8051_indi_addr1_n17), .Y(ri[3]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u30 ( .A(wr_dat[4]), .B(
        oc8051_indi_addr1_n102), .S0(oc8051_indi_addr1_n17), .Y(ri[4]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u29 ( .A(wr_dat[5]), .B(
        oc8051_indi_addr1_n101), .S0(oc8051_indi_addr1_n17), .Y(ri[5]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u28 ( .A(wr_dat[6]), .B(
        oc8051_indi_addr1_n100), .S0(oc8051_indi_addr1_n17), .Y(ri[6]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u27 ( .A(wr_dat[7]), .B(
        oc8051_indi_addr1_n99), .S0(oc8051_indi_addr1_n17), .Y(ri[7]) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u26 ( .A(oc8051_indi_addr1_buff_4__1_), .B(
        oc8051_indi_addr1_buff_6__1_), .C(oc8051_indi_addr1_buff_5__1_), .D(
        oc8051_indi_addr1_buff_7__1_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n16) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u25 ( .A(oc8051_indi_addr1_buff_0__1_), .B(
        oc8051_indi_addr1_buff_2__1_), .C(oc8051_indi_addr1_buff_1__1_), .D(
        oc8051_indi_addr1_buff_3__1_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n15) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u24 ( .A(oc8051_indi_addr1_n15), .B(
        oc8051_indi_addr1_n16), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n105)
         );
  MXT4_X1M_A12TS oc8051_indi_addr1_u23 ( .A(oc8051_indi_addr1_buff_4__0_), .B(
        oc8051_indi_addr1_buff_6__0_), .C(oc8051_indi_addr1_buff_5__0_), .D(
        oc8051_indi_addr1_buff_7__0_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n14) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u22 ( .A(oc8051_indi_addr1_buff_0__0_), .B(
        oc8051_indi_addr1_buff_2__0_), .C(oc8051_indi_addr1_buff_1__0_), .D(
        oc8051_indi_addr1_buff_3__0_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n13) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u21 ( .A(oc8051_indi_addr1_n13), .B(
        oc8051_indi_addr1_n14), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n106)
         );
  MXT4_X1M_A12TS oc8051_indi_addr1_u20 ( .A(oc8051_indi_addr1_buff_4__2_), .B(
        oc8051_indi_addr1_buff_6__2_), .C(oc8051_indi_addr1_buff_5__2_), .D(
        oc8051_indi_addr1_buff_7__2_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n12) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u19 ( .A(oc8051_indi_addr1_buff_0__2_), .B(
        oc8051_indi_addr1_buff_2__2_), .C(oc8051_indi_addr1_buff_1__2_), .D(
        oc8051_indi_addr1_buff_3__2_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n11) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u18 ( .A(oc8051_indi_addr1_n11), .B(
        oc8051_indi_addr1_n12), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n104)
         );
  MXT4_X1M_A12TS oc8051_indi_addr1_u17 ( .A(oc8051_indi_addr1_buff_4__3_), .B(
        oc8051_indi_addr1_buff_6__3_), .C(oc8051_indi_addr1_buff_5__3_), .D(
        oc8051_indi_addr1_buff_7__3_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n10) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u16 ( .A(oc8051_indi_addr1_buff_0__3_), .B(
        oc8051_indi_addr1_buff_2__3_), .C(oc8051_indi_addr1_buff_1__3_), .D(
        oc8051_indi_addr1_buff_3__3_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n9) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u15 ( .A(oc8051_indi_addr1_n9), .B(
        oc8051_indi_addr1_n10), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n103)
         );
  MXT4_X1M_A12TS oc8051_indi_addr1_u14 ( .A(oc8051_indi_addr1_buff_4__6_), .B(
        oc8051_indi_addr1_buff_6__6_), .C(oc8051_indi_addr1_buff_5__6_), .D(
        oc8051_indi_addr1_buff_7__6_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n8) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u13 ( .A(oc8051_indi_addr1_buff_0__6_), .B(
        oc8051_indi_addr1_buff_2__6_), .C(oc8051_indi_addr1_buff_1__6_), .D(
        oc8051_indi_addr1_buff_3__6_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n7) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u12 ( .A(oc8051_indi_addr1_n7), .B(
        oc8051_indi_addr1_n8), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n100) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u11 ( .A(oc8051_indi_addr1_buff_4__7_), .B(
        oc8051_indi_addr1_buff_6__7_), .C(oc8051_indi_addr1_buff_5__7_), .D(
        oc8051_indi_addr1_buff_7__7_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n6) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u10 ( .A(oc8051_indi_addr1_buff_0__7_), .B(
        oc8051_indi_addr1_buff_2__7_), .C(oc8051_indi_addr1_buff_1__7_), .D(
        oc8051_indi_addr1_buff_3__7_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n5) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u9 ( .A(oc8051_indi_addr1_n5), .B(
        oc8051_indi_addr1_n6), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n99) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u8 ( .A(oc8051_indi_addr1_buff_4__5_), .B(
        oc8051_indi_addr1_buff_6__5_), .C(oc8051_indi_addr1_buff_5__5_), .D(
        oc8051_indi_addr1_buff_7__5_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n4) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u7 ( .A(oc8051_indi_addr1_buff_0__5_), .B(
        oc8051_indi_addr1_buff_2__5_), .C(oc8051_indi_addr1_buff_1__5_), .D(
        oc8051_indi_addr1_buff_3__5_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n3) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u6 ( .A(oc8051_indi_addr1_n3), .B(
        oc8051_indi_addr1_n4), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n101) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u5 ( .A(oc8051_indi_addr1_buff_4__4_), .B(
        oc8051_indi_addr1_buff_6__4_), .C(oc8051_indi_addr1_buff_5__4_), .D(
        oc8051_indi_addr1_buff_7__4_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n2) );
  MXT4_X1M_A12TS oc8051_indi_addr1_u4 ( .A(oc8051_indi_addr1_buff_0__4_), .B(
        oc8051_indi_addr1_buff_2__4_), .C(oc8051_indi_addr1_buff_1__4_), .D(
        oc8051_indi_addr1_buff_3__4_), .S0(bank_sel[0]), .S1(op1_cur[0]), .Y(
        oc8051_indi_addr1_n1) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u3 ( .A(oc8051_indi_addr1_n1), .B(
        oc8051_indi_addr1_n2), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n102) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__0_ ( .D(oc8051_indi_addr1_n83), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__1_ ( .D(oc8051_indi_addr1_n82), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__2_ ( .D(oc8051_indi_addr1_n81), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__3_ ( .D(oc8051_indi_addr1_n80), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__4_ ( .D(oc8051_indi_addr1_n79), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__5_ ( .D(oc8051_indi_addr1_n78), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__6_ ( .D(oc8051_indi_addr1_n77), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__7_ ( .D(oc8051_indi_addr1_n76), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__0_ ( .D(oc8051_indi_addr1_n51), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__1_ ( .D(oc8051_indi_addr1_n50), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__2_ ( .D(oc8051_indi_addr1_n49), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__3_ ( .D(oc8051_indi_addr1_n48), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__4_ ( .D(oc8051_indi_addr1_n47), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__5_ ( .D(oc8051_indi_addr1_n46), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__6_ ( .D(oc8051_indi_addr1_n45), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__7_ ( .D(oc8051_indi_addr1_n44), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__0_ ( .D(oc8051_indi_addr1_n67), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__1_ ( .D(oc8051_indi_addr1_n66), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__2_ ( .D(oc8051_indi_addr1_n65), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__3_ ( .D(oc8051_indi_addr1_n64), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__4_ ( .D(oc8051_indi_addr1_n63), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__5_ ( .D(oc8051_indi_addr1_n62), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__6_ ( .D(oc8051_indi_addr1_n61), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__7_ ( .D(oc8051_indi_addr1_n60), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__0_ ( .D(oc8051_indi_addr1_n35), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__1_ ( .D(oc8051_indi_addr1_n34), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__2_ ( .D(oc8051_indi_addr1_n33), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__3_ ( .D(oc8051_indi_addr1_n32), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__4_ ( .D(oc8051_indi_addr1_n31), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__5_ ( .D(oc8051_indi_addr1_n30), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__6_ ( .D(oc8051_indi_addr1_n29), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__7_ ( .D(oc8051_indi_addr1_n28), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__0_ ( .D(oc8051_indi_addr1_n75), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__1_ ( .D(oc8051_indi_addr1_n74), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__2_ ( .D(oc8051_indi_addr1_n73), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__3_ ( .D(oc8051_indi_addr1_n72), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__4_ ( .D(oc8051_indi_addr1_n71), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__5_ ( .D(oc8051_indi_addr1_n70), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__6_ ( .D(oc8051_indi_addr1_n69), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__7_ ( .D(oc8051_indi_addr1_n68), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__0_ ( .D(oc8051_indi_addr1_n43), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__1_ ( .D(oc8051_indi_addr1_n42), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__2_ ( .D(oc8051_indi_addr1_n41), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__3_ ( .D(oc8051_indi_addr1_n40), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__4_ ( .D(oc8051_indi_addr1_n39), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__5_ ( .D(oc8051_indi_addr1_n38), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__6_ ( .D(oc8051_indi_addr1_n37), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__7_ ( .D(oc8051_indi_addr1_n36), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__0_ ( .D(oc8051_indi_addr1_n91), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__1_ ( .D(oc8051_indi_addr1_n90), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__2_ ( .D(oc8051_indi_addr1_n89), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__3_ ( .D(oc8051_indi_addr1_n88), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__4_ ( .D(oc8051_indi_addr1_n87), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__5_ ( .D(oc8051_indi_addr1_n86), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__6_ ( .D(oc8051_indi_addr1_n85), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__7_ ( .D(oc8051_indi_addr1_n84), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__0_ ( .D(oc8051_indi_addr1_n59), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__1_ ( .D(oc8051_indi_addr1_n58), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__2_ ( .D(oc8051_indi_addr1_n57), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__3_ ( .D(oc8051_indi_addr1_n56), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__4_ ( .D(oc8051_indi_addr1_n55), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__5_ ( .D(oc8051_indi_addr1_n54), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__6_ ( .D(oc8051_indi_addr1_n53), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__7_ ( .D(oc8051_indi_addr1_n52), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_wr_bit_r_reg ( .D(bit_addr_o), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_wr_bit_r) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u833 ( .AN(mem_act[0]), .B(
        wbd_ack_i), .Y(oc8051_memory_interface1_n1290) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u832 ( .A(
        oc8051_memory_interface1_op1_5_), .Y(oc8051_memory_interface1_n649) );
  OR3_X0P5M_A12TS oc8051_memory_interface1_u831 ( .A(
        oc8051_memory_interface1_pc_wr_r2), .B(
        oc8051_memory_interface1_imem_wait), .C(
        oc8051_memory_interface1_dmem_wait), .Y(mem_wait) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u830 ( .A(rd), .Y(
        oc8051_memory_interface1_n258) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u829 ( .A(
        oc8051_memory_interface1_int_ack_t), .Y(oc8051_memory_interface1_n257)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u828 ( .A(n_logic0_), .B(ea_in), 
        .Y(oc8051_memory_interface1_n297) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u827 ( .A(
        oc8051_memory_interface1_n297), .Y(oc8051_memory_interface1_n242) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u826 ( .A(
        oc8051_memory_interface1_n242), .B(wbi_ack_i), .Y(
        oc8051_memory_interface1_n243) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u825 ( .A(
        oc8051_memory_interface1_n257), .B(oc8051_memory_interface1_n243), .Y(
        oc8051_memory_interface1_n597) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u824 ( .A(
        oc8051_memory_interface1_n258), .B(oc8051_memory_interface1_n597), .Y(
        oc8051_memory_interface1_n386) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u823 ( .A(
        oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n341) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u822 ( .A(
        oc8051_memory_interface1_n649), .B(mem_wait), .C(
        oc8051_memory_interface1_n341), .Y(oc8051_memory_interface1_n646) );
  OR3_X0P5M_A12TS oc8051_memory_interface1_u821 ( .A(
        oc8051_memory_interface1_op1_6_), .B(oc8051_memory_interface1_op1_7_), 
        .C(oc8051_memory_interface1_op1_3_), .Y(oc8051_memory_interface1_n648)
         );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u820 ( .A(
        oc8051_memory_interface1_n648), .B(oc8051_memory_interface1_op1_2_), 
        .C(oc8051_memory_interface1_op1_0_), .Y(oc8051_memory_interface1_n647)
         );
  AND4_X0P5M_A12TS oc8051_memory_interface1_u819 ( .A(
        oc8051_memory_interface1_op1_4_), .B(oc8051_memory_interface1_op1_1_), 
        .C(oc8051_memory_interface1_n646), .D(oc8051_memory_interface1_n647), 
        .Y(oc8051_memory_interface1_n1980) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u818 ( .AN(
        oc8051_memory_interface1_int_ack_buff), .B(
        oc8051_memory_interface1_int_ack_t), .Y(oc8051_memory_interface1_n3700) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u817 ( .A(
        oc8051_memory_interface1_cdone), .B(oc8051_memory_interface1_dack_ir), 
        .Y(oc8051_memory_interface1_n643) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u816 ( .AN(
        oc8051_memory_interface1_n643), .B(oc8051_memory_interface1_n597), .Y(
        oc8051_memory_interface1_n639) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u815 ( .AN(
        oc8051_memory_interface1_cdone), .B(oc8051_memory_interface1_dack_ir), 
        .Y(oc8051_memory_interface1_n640) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u814 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_6_), .B0(
        oc8051_memory_interface1_n639), .B1(oc8051_memory_interface1_op1_6_), 
        .C0(oc8051_memory_interface1_cdata_6_), .C1(
        oc8051_memory_interface1_n640), .Y(oc8051_memory_interface1_n602) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u813 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_0_), .B0(
        oc8051_memory_interface1_n639), .B1(oc8051_memory_interface1_op1_0_), 
        .C0(oc8051_memory_interface1_cdata_0_), .C1(
        oc8051_memory_interface1_n640), .Y(oc8051_memory_interface1_n618) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u812 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_3_), .B0(
        oc8051_memory_interface1_n639), .B1(oc8051_memory_interface1_op1_3_), 
        .C0(oc8051_memory_interface1_cdata_3_), .C1(
        oc8051_memory_interface1_n640), .Y(oc8051_memory_interface1_n611) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u811 ( .A(
        oc8051_memory_interface1_n611), .Y(op1_n[3]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u810 ( .A(
        oc8051_memory_interface1_n618), .B(op1_n[3]), .Y(
        oc8051_memory_interface1_n641) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u809 ( .A0(
        oc8051_memory_interface1_ddat_ir_4_), .A1(
        oc8051_memory_interface1_dack_ir), .B0(oc8051_memory_interface1_n640), 
        .B1(oc8051_memory_interface1_cdata_4_), .Y(
        oc8051_memory_interface1_n645) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u808 ( .A0(
        oc8051_memory_interface1_n597), .A1(oc8051_memory_interface1_op1_4_), 
        .B0(oc8051_memory_interface1_n643), .C0(oc8051_memory_interface1_n645), 
        .Y(oc8051_memory_interface1_n606) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u807 ( .A(
        oc8051_memory_interface1_n606), .Y(op1_n[4]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u806 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_2_), .B0(
        oc8051_memory_interface1_n639), .B1(oc8051_memory_interface1_op1_2_), 
        .C0(oc8051_memory_interface1_cdata_2_), .C1(
        oc8051_memory_interface1_n640), .Y(oc8051_memory_interface1_n632) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u805 ( .A(
        oc8051_memory_interface1_n632), .Y(op1_n[2]) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u804 ( .A0(
        oc8051_memory_interface1_ddat_ir_1_), .A1(
        oc8051_memory_interface1_dack_ir), .B0(oc8051_memory_interface1_n640), 
        .B1(oc8051_memory_interface1_cdata_1_), .Y(
        oc8051_memory_interface1_n644) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u803 ( .A0(
        oc8051_memory_interface1_n597), .A1(oc8051_memory_interface1_op1_1_), 
        .B0(oc8051_memory_interface1_n643), .C0(oc8051_memory_interface1_n644), 
        .Y(oc8051_memory_interface1_n613) );
  NAND4_X0P5A_A12TS oc8051_memory_interface1_u802 ( .A(
        oc8051_memory_interface1_n641), .B(op1_n[4]), .C(op1_n[2]), .D(
        oc8051_memory_interface1_n613), .Y(oc8051_memory_interface1_n642) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u801 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_7_), .B0(
        oc8051_memory_interface1_n639), .B1(oc8051_memory_interface1_op1_7_), 
        .C0(oc8051_memory_interface1_cdata_7_), .C1(
        oc8051_memory_interface1_n640), .Y(oc8051_memory_interface1_n604) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u800 ( .A(
        oc8051_memory_interface1_n641), .B(oc8051_memory_interface1_n642), 
        .S0(oc8051_memory_interface1_n604), .Y(oc8051_memory_interface1_n638)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u799 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_5_), .B0(
        oc8051_memory_interface1_n639), .B1(oc8051_memory_interface1_op1_5_), 
        .C0(oc8051_memory_interface1_cdata_5_), .C1(
        oc8051_memory_interface1_n640), .Y(oc8051_memory_interface1_n610) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u798 ( .A(
        oc8051_memory_interface1_n610), .Y(op1_n[5]) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u797 ( .A0(
        oc8051_memory_interface1_n632), .A1(oc8051_memory_interface1_n613), 
        .B0(oc8051_memory_interface1_n611), .Y(oc8051_memory_interface1_n635)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u796 ( .A0(
        oc8051_memory_interface1_n638), .A1(op1_n[5]), .B0(
        oc8051_memory_interface1_n635), .B1(oc8051_memory_interface1_n606), 
        .Y(oc8051_memory_interface1_n625) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u795 ( .A(
        oc8051_memory_interface1_n613), .Y(op1_n[1]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u794 ( .A(
        oc8051_memory_interface1_n606), .B(op1_n[5]), .Y(
        oc8051_memory_interface1_n605) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u793 ( .A(
        oc8051_memory_interface1_n602), .Y(op1_n[6]) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u792 ( .A(op1_n[6]), .B(op1_n[1]), 
        .C(op1_n[4]), .Y(oc8051_memory_interface1_n616) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u791 ( .A0(op1_n[1]), .A1(
        op1_n[4]), .B0(oc8051_memory_interface1_n605), .B1(op1_n[6]), .C0(
        oc8051_memory_interface1_n616), .Y(oc8051_memory_interface1_n636) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u790 ( .A(
        oc8051_memory_interface1_n606), .B(op1_n[6]), .Y(
        oc8051_memory_interface1_n624) );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u789 ( .A0(
        oc8051_memory_interface1_n606), .A1(oc8051_memory_interface1_n618), 
        .A2(op1_n[6]), .B0(oc8051_memory_interface1_n624), .B1(op1_n[5]), .Y(
        oc8051_memory_interface1_n637) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u788 ( .A0(op1_n[3]), .A1(
        oc8051_memory_interface1_n636), .B0(oc8051_memory_interface1_n637), 
        .C0(oc8051_memory_interface1_n632), .Y(oc8051_memory_interface1_n629)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u787 ( .A(
        oc8051_memory_interface1_n635), .Y(oc8051_memory_interface1_n603) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u786 ( .A(
        oc8051_memory_interface1_n611), .B(oc8051_memory_interface1_n613), .Y(
        oc8051_memory_interface1_n633) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u785 ( .A(
        oc8051_memory_interface1_n618), .B(oc8051_memory_interface1_n610), .Y(
        oc8051_memory_interface1_n617) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u784 ( .A(
        oc8051_memory_interface1_n617), .Y(oc8051_memory_interface1_n634) );
  AOI211_X0P5M_A12TS oc8051_memory_interface1_u783 ( .A0(
        oc8051_memory_interface1_n632), .A1(oc8051_memory_interface1_n618), 
        .B0(oc8051_memory_interface1_n633), .C0(oc8051_memory_interface1_n634), 
        .Y(oc8051_memory_interface1_n631) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u782 ( .A0(op1_n[5]), .A1(
        oc8051_memory_interface1_n603), .B0(op1_n[6]), .B1(
        oc8051_memory_interface1_n631), .Y(oc8051_memory_interface1_n630) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u781 ( .A(
        oc8051_memory_interface1_n629), .B(oc8051_memory_interface1_n630), 
        .S0(oc8051_memory_interface1_n604), .Y(oc8051_memory_interface1_n626)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u780 ( .A(
        oc8051_memory_interface1_n618), .Y(op1_n[0]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u779 ( .A(op1_n[2]), .B(op1_n[3]), 
        .Y(oc8051_memory_interface1_n612) );
  OAI31_X0P5M_A12TS oc8051_memory_interface1_u778 ( .A0(
        oc8051_memory_interface1_n617), .A1(op1_n[1]), .A2(op1_n[2]), .B0(
        oc8051_memory_interface1_n611), .Y(oc8051_memory_interface1_n628) );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u777 ( .A0(op1_n[1]), .A1(
        op1_n[0]), .A2(oc8051_memory_interface1_n612), .B0(
        oc8051_memory_interface1_n624), .B1(oc8051_memory_interface1_n628), 
        .Y(oc8051_memory_interface1_n627) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u776 ( .A0(
        oc8051_memory_interface1_n602), .A1(oc8051_memory_interface1_n625), 
        .B0(oc8051_memory_interface1_n626), .C0(oc8051_memory_interface1_n627), 
        .Y(oc8051_memory_interface1_n4250) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u775 ( .A0(op1_n[0]), .A1(
        oc8051_memory_interface1_n604), .B0(op1_n[6]), .Y(
        oc8051_memory_interface1_n622) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u774 ( .A(
        oc8051_memory_interface1_n624), .B(op1_n[5]), .S0(
        oc8051_memory_interface1_n604), .Y(oc8051_memory_interface1_n623) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u773 ( .A0(op1_n[5]), .A1(
        oc8051_memory_interface1_n618), .B0(oc8051_memory_interface1_n622), 
        .C0(oc8051_memory_interface1_n623), .Y(oc8051_memory_interface1_n614)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u772 ( .A(
        oc8051_memory_interface1_n604), .Y(op1_n[7]) );
  AOI31_X0P5M_A12TS oc8051_memory_interface1_u771 ( .A0(op1_n[0]), .A1(
        op1_n[5]), .A2(op1_n[4]), .B0(op1_n[7]), .Y(
        oc8051_memory_interface1_n620) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u770 ( .A(
        oc8051_memory_interface1_n604), .B(op1_n[0]), .Y(
        oc8051_memory_interface1_n621) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u769 ( .A(
        oc8051_memory_interface1_n620), .B(oc8051_memory_interface1_n621), 
        .S0(oc8051_memory_interface1_n602), .Y(oc8051_memory_interface1_n619)
         );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u768 ( .A0(
        oc8051_memory_interface1_n616), .A1(oc8051_memory_interface1_n617), 
        .B0(op1_n[1]), .B1(oc8051_memory_interface1_n618), .C0(
        oc8051_memory_interface1_n619), .Y(oc8051_memory_interface1_n615) );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u767 ( .A0(
        oc8051_memory_interface1_n611), .A1(oc8051_memory_interface1_n613), 
        .A2(oc8051_memory_interface1_n614), .B0(oc8051_memory_interface1_n612), 
        .B1(oc8051_memory_interface1_n615), .Y(oc8051_memory_interface1_n598)
         );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u766 ( .A(op1_n[7]), .B(
        oc8051_memory_interface1_n612), .Y(oc8051_memory_interface1_n608) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u765 ( .A(
        oc8051_memory_interface1_n611), .B(oc8051_memory_interface1_n604), .Y(
        oc8051_memory_interface1_n609) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u764 ( .A(
        oc8051_memory_interface1_n608), .B(oc8051_memory_interface1_n609), 
        .S0(oc8051_memory_interface1_n610), .Y(oc8051_memory_interface1_n607)
         );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u763 ( .A(
        oc8051_memory_interface1_n606), .B(oc8051_memory_interface1_n607), .Y(
        oc8051_memory_interface1_n600) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u762 ( .A(
        oc8051_memory_interface1_n603), .B(oc8051_memory_interface1_n604), .C(
        oc8051_memory_interface1_n605), .Y(oc8051_memory_interface1_n601) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u761 ( .A(
        oc8051_memory_interface1_n600), .B(oc8051_memory_interface1_n601), 
        .S0(oc8051_memory_interface1_n602), .Y(oc8051_memory_interface1_n599)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u760 ( .A(
        oc8051_memory_interface1_n598), .B(oc8051_memory_interface1_n599), .Y(
        oc8051_memory_interface1_n4260) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u759 ( .A(pc_wr_sel[2]), .Y(
        oc8051_memory_interface1_n397) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u758 ( .A(pc_wr_sel[1]), .Y(
        oc8051_memory_interface1_n361) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u757 ( .A(
        oc8051_memory_interface1_n397), .B(oc8051_memory_interface1_n361), .Y(
        oc8051_memory_interface1_n365) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u756 ( .A(
        oc8051_memory_interface1_n365), .Y(oc8051_memory_interface1_n576) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u755 ( .A(n_3_net_), .Y(
        oc8051_memory_interface1_n398) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u754 ( .A0(
        oc8051_memory_interface1_n576), .A1(pc_wr_sel[0]), .B0(
        oc8051_memory_interface1_n398), .Y(oc8051_memory_interface1_n5360) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u753 ( .A(ram_rd_sel[0]), .Y(
        oc8051_memory_interface1_n180) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u752 ( .A(
        oc8051_memory_interface1_n180), .B(ram_rd_sel[2]), .Y(
        oc8051_memory_interface1_n810) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u751 ( .A(ram_wr_sel[1]), .Y(
        oc8051_memory_interface1_n153) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u750 ( .A(
        oc8051_memory_interface1_n153), .B(ram_wr_sel[2]), .Y(wr_ind) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u749 ( .A0(
        oc8051_memory_interface1_op2_buff[7]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[7]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n359)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u748 ( .A(
        oc8051_memory_interface1_n359), .Y(op2_n[7]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u747 ( .A(
        oc8051_memory_interface1_n597), .B(rd), .Y(
        oc8051_memory_interface1_n342) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u746 ( .A0(
        oc8051_memory_interface1_op3[7]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_7_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[7]), .Y(
        oc8051_memory_interface1_n360) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u745 ( .A(
        oc8051_memory_interface1_n360), .Y(op3_n[7]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u744 ( .A(op2_n[7]), .B(op3_n[7]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n579) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u743 ( .A(
        oc8051_memory_interface1_n579), .Y(
        oc8051_memory_interface1_pcs_source_7_) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u742 ( .A(
        oc8051_memory_interface1_n380), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_10) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u741 ( .A(
        oc8051_memory_interface1_n379), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_11) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u740 ( .A(
        oc8051_memory_interface1_n378), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_12) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u739 ( .A(
        oc8051_memory_interface1_n377), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_13) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u738 ( .A(
        oc8051_memory_interface1_n383), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_14) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u737 ( .A(
        oc8051_memory_interface1_n384), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_15) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u736 ( .A(
        oc8051_memory_interface1_n382), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_8) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u735 ( .A(
        oc8051_memory_interface1_n381), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_u3_u7_z_9) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u734 ( .A(
        oc8051_memory_interface1_pc_buf_0_), .Y(oc8051_memory_interface1_n304)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u733 ( .A(
        oc8051_memory_interface1_iadr_t_0_), .Y(oc8051_memory_interface1_n594)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u732 ( .A(
        oc8051_memory_interface1_n304), .B(oc8051_memory_interface1_n594), 
        .S0(oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[0]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u731 ( .A(
        oc8051_memory_interface1_iadr_t_10_), .Y(oc8051_memory_interface1_n585) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u730 ( .A(
        oc8051_memory_interface1_n35), .B(oc8051_memory_interface1_n585), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[10]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u729 ( .A(
        oc8051_memory_interface1_iadr_t_11_), .Y(oc8051_memory_interface1_n584) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u728 ( .A(
        oc8051_memory_interface1_n41), .B(oc8051_memory_interface1_n584), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[11]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u727 ( .A(
        oc8051_memory_interface1_iadr_t_12_), .Y(oc8051_memory_interface1_n583) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u726 ( .A(
        oc8051_memory_interface1_n39), .B(oc8051_memory_interface1_n583), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[12]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u725 ( .A(
        oc8051_memory_interface1_iadr_t_13_), .Y(oc8051_memory_interface1_n582) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u724 ( .A(
        oc8051_memory_interface1_n38), .B(oc8051_memory_interface1_n582), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[13]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u723 ( .A(
        oc8051_memory_interface1_iadr_t_14_), .Y(oc8051_memory_interface1_n580) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u722 ( .A(
        oc8051_memory_interface1_n40), .B(oc8051_memory_interface1_n580), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[14]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u721 ( .A(
        oc8051_memory_interface1_pc_out_15_), .B(
        oc8051_memory_interface1_iadr_t_15_), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[15]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u720 ( .A(
        oc8051_memory_interface1_pc_buf_1_), .Y(oc8051_memory_interface1_n308)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u719 ( .A(
        oc8051_memory_interface1_iadr_t_1_), .Y(oc8051_memory_interface1_n593)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u718 ( .A(
        oc8051_memory_interface1_n308), .B(oc8051_memory_interface1_n593), 
        .S0(oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[1]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u717 ( .A(
        oc8051_memory_interface1_iadr_t_2_), .Y(oc8051_memory_interface1_n592)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u716 ( .A(
        oc8051_memory_interface1_n29), .B(oc8051_memory_interface1_n592), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[2]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u715 ( .A(
        oc8051_memory_interface1_iadr_t_3_), .Y(oc8051_memory_interface1_n591)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u714 ( .A(
        oc8051_memory_interface1_n30), .B(oc8051_memory_interface1_n591), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[3]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u713 ( .A(
        oc8051_memory_interface1_iadr_t_4_), .Y(oc8051_memory_interface1_n590)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u712 ( .A(
        oc8051_memory_interface1_n31), .B(oc8051_memory_interface1_n590), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[4]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u711 ( .A(
        oc8051_memory_interface1_iadr_t_5_), .Y(oc8051_memory_interface1_n589)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u710 ( .A(
        oc8051_memory_interface1_n33), .B(oc8051_memory_interface1_n589), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[5]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u709 ( .A(
        oc8051_memory_interface1_iadr_t_6_), .Y(oc8051_memory_interface1_n588)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u708 ( .A(
        oc8051_memory_interface1_n32), .B(oc8051_memory_interface1_n588), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[6]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u707 ( .A(
        oc8051_memory_interface1_pc_out_7_), .B(
        oc8051_memory_interface1_iadr_t_7_), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[7]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u706 ( .A(
        oc8051_memory_interface1_iadr_t_8_), .Y(oc8051_memory_interface1_n587)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u705 ( .A(
        oc8051_memory_interface1_n37), .B(oc8051_memory_interface1_n587), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[8]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u704 ( .A(
        oc8051_memory_interface1_iadr_t_9_), .Y(oc8051_memory_interface1_n586)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u703 ( .A(
        oc8051_memory_interface1_n36), .B(oc8051_memory_interface1_n586), .S0(
        oc8051_memory_interface1_istb_t), .Y(wbi_adr_o[9]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u702 ( .A(
        oc8051_memory_interface1_pc_wr_r2), .Y(oc8051_memory_interface1_n301)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u701 ( .A0(
        oc8051_memory_interface1_op_pos_1_), .A1(
        oc8051_memory_interface1_op_pos_0_), .B0(
        oc8051_memory_interface1_op_pos_2_), .C0(rd), .Y(
        oc8051_memory_interface1_n596) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u700 ( .A(
        oc8051_memory_interface1_n301), .B(oc8051_memory_interface1_n596), .Y(
        oc8051_memory_interface1_inc_pc) );
  NAND2B_X0P5M_A12TS oc8051_memory_interface1_u699 ( .AN(
        oc8051_memory_interface1_rd_ind), .B(
        oc8051_memory_interface1_rd_addr_r), .Y(oc8051_memory_interface1_n322)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u698 ( .A(
        oc8051_memory_interface1_n322), .Y(oc8051_memory_interface1_n674) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u697 ( .A(ram_data[0]), .B(
        sfr_out[0]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[0]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u696 ( .A(ram_data[1]), .B(
        sfr_out[1]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[1]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u695 ( .A(ram_data[2]), .B(
        sfr_out[2]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[2]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u694 ( .A(ram_data[3]), .B(
        sfr_out[3]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[3]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u693 ( .A(ram_data[4]), .B(
        sfr_out[4]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[4]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u692 ( .A(ram_data[5]), .B(
        sfr_out[5]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[5]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u691 ( .A(ram_data[6]), .B(
        sfr_out[6]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[6]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u690 ( .A(ram_data[7]), .B(
        sfr_out[7]), .S0(oc8051_memory_interface1_n674), .Y(ram_out[7]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u689 ( .A(
        oc8051_memory_interface1_istb_t), .B(oc8051_memory_interface1_n297), 
        .Y(oc8051_memory_interface1_n233) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u688 ( .A(istb), .B(
        oc8051_memory_interface1_n297), .Y(oc8051_memory_interface1_n595) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u687 ( .A0(wbi_ack_i), .A1(
        oc8051_memory_interface1_n233), .B0(oc8051_memory_interface1_n595), 
        .C0(wbd_cyc_o), .Y(oc8051_memory_interface1_istb_o) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u686 ( .A(
        oc8051_memory_interface1_ddat_ir_0_), .B(wbd_dat_i[0]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n401) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u685 ( .A(
        oc8051_memory_interface1_ddat_ir_1_), .B(wbd_dat_i[1]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n402) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u684 ( .A(
        oc8051_memory_interface1_ddat_ir_2_), .B(wbd_dat_i[2]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n403) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u683 ( .A(
        oc8051_memory_interface1_ddat_ir_3_), .B(wbd_dat_i[3]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n404) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u682 ( .A(
        oc8051_memory_interface1_ddat_ir_4_), .B(wbd_dat_i[4]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n405) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u681 ( .A(
        oc8051_memory_interface1_ddat_ir_5_), .B(wbd_dat_i[5]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n406) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u680 ( .A(
        oc8051_memory_interface1_ddat_ir_6_), .B(wbd_dat_i[6]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n407) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u679 ( .A(
        oc8051_memory_interface1_ddat_ir_7_), .B(wbd_dat_i[7]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n408) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u678 ( .A(
        oc8051_memory_interface1_int_vec_buff_0_), .B(int_src[0]), .S0(intr), 
        .Y(oc8051_memory_interface1_n409) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u677 ( .A(
        oc8051_memory_interface1_int_vec_buff_1_), .B(int_src[1]), .S0(intr), 
        .Y(oc8051_memory_interface1_n410) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u676 ( .A(
        oc8051_memory_interface1_int_vec_buff_2_), .B(n_logic0_), .S0(intr), 
        .Y(oc8051_memory_interface1_n411) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u675 ( .A(
        oc8051_memory_interface1_int_vec_buff_3_), .B(int_src[3]), .S0(intr), 
        .Y(oc8051_memory_interface1_n412) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u674 ( .A(
        oc8051_memory_interface1_int_vec_buff_4_), .B(int_src[4]), .S0(intr), 
        .Y(oc8051_memory_interface1_n413) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u673 ( .A(
        oc8051_memory_interface1_int_vec_buff_5_), .B(int_src[5]), .S0(intr), 
        .Y(oc8051_memory_interface1_n414) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u672 ( .A(
        oc8051_memory_interface1_int_vec_buff_6_), .B(n_logic0_), .S0(intr), 
        .Y(oc8051_memory_interface1_n415) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u671 ( .A(
        oc8051_memory_interface1_int_vec_buff_7_), .B(n_logic0_), .S0(intr), 
        .Y(oc8051_memory_interface1_n416) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u670 ( .A(des_acc[0]), .Y(
        oc8051_memory_interface1_n373) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u669 ( .A(mem_act[1]), .Y(
        oc8051_memory_interface1_n255) );
  NAND3B_X0P5M_A12TS oc8051_memory_interface1_u668 ( .AN(mem_act[0]), .B(
        oc8051_memory_interface1_n255), .C(mem_act[2]), .Y(
        oc8051_memory_interface1_n244) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u667 ( .A(
        oc8051_memory_interface1_n244), .Y(oc8051_memory_interface1_n581) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u666 ( .A(
        oc8051_memory_interface1_n594), .B(oc8051_memory_interface1_n373), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n425)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u665 ( .A(des_acc[1]), .Y(
        oc8051_memory_interface1_n390) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u664 ( .A(
        oc8051_memory_interface1_n593), .B(oc8051_memory_interface1_n390), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n426)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u663 ( .A(des_acc[2]), .Y(
        oc8051_memory_interface1_n395) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u662 ( .A(
        oc8051_memory_interface1_n592), .B(oc8051_memory_interface1_n395), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n427)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u661 ( .A(des_acc[3]), .Y(
        oc8051_memory_interface1_n421) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u660 ( .A(
        oc8051_memory_interface1_n591), .B(oc8051_memory_interface1_n421), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n428)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u659 ( .A(des_acc[4]), .Y(
        oc8051_memory_interface1_n442) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u658 ( .A(
        oc8051_memory_interface1_n590), .B(oc8051_memory_interface1_n442), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n429)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u657 ( .A(des_acc[5]), .Y(
        oc8051_memory_interface1_n533) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u656 ( .A(
        oc8051_memory_interface1_n589), .B(oc8051_memory_interface1_n533), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n430)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u655 ( .A(des_acc[6]), .Y(
        oc8051_memory_interface1_n570) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u654 ( .A(
        oc8051_memory_interface1_n588), .B(oc8051_memory_interface1_n570), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n431)
         );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u653 ( .A(des_acc[7]), .B(
        oc8051_memory_interface1_iadr_t_7_), .S0(oc8051_memory_interface1_n244), .Y(oc8051_memory_interface1_n432) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u652 ( .A(des2[0]), .Y(
        oc8051_memory_interface1_n372) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u651 ( .A(
        oc8051_memory_interface1_n587), .B(oc8051_memory_interface1_n372), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n433)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u650 ( .A(des2[1]), .Y(
        oc8051_memory_interface1_n389) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u649 ( .A(
        oc8051_memory_interface1_n586), .B(oc8051_memory_interface1_n389), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n434)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u648 ( .A(des2[2]), .Y(
        oc8051_memory_interface1_n394) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u647 ( .A(
        oc8051_memory_interface1_n585), .B(oc8051_memory_interface1_n394), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n435)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u646 ( .A(des2[3]), .Y(
        oc8051_memory_interface1_n420) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u645 ( .A(
        oc8051_memory_interface1_n584), .B(oc8051_memory_interface1_n420), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n436)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u644 ( .A(des2[4]), .Y(
        oc8051_memory_interface1_n441) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u643 ( .A(
        oc8051_memory_interface1_n583), .B(oc8051_memory_interface1_n441), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n437)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u642 ( .A(des2[5]), .Y(
        oc8051_memory_interface1_n531) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u641 ( .A(
        oc8051_memory_interface1_n582), .B(oc8051_memory_interface1_n531), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n438)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u640 ( .A(des2[6]), .Y(
        oc8051_memory_interface1_n541) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u639 ( .A(
        oc8051_memory_interface1_n580), .B(oc8051_memory_interface1_n541), 
        .S0(oc8051_memory_interface1_n581), .Y(oc8051_memory_interface1_n439)
         );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u638 ( .A(des2[7]), .B(
        oc8051_memory_interface1_iadr_t_15_), .S0(
        oc8051_memory_interface1_n244), .Y(oc8051_memory_interface1_n440) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u637 ( .A(pc_wr_sel[0]), .B(
        pc_wr_sel[1]), .C(oc8051_memory_interface1_n398), .Y(
        oc8051_memory_interface1_n399) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u636 ( .A(pc_wr_sel[2]), .B(
        pc_wr_sel[1]), .Y(oc8051_memory_interface1_n366) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u635 ( .A(
        oc8051_memory_interface1_n366), .Y(oc8051_memory_interface1_n575) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u634 ( .A(pc_wr_sel[2]), .B(
        oc8051_memory_interface1_n361), .Y(oc8051_memory_interface1_n400) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u633 ( .A(
        oc8051_memory_interface1_n361), .B(pc_wr_sel[2]), .Y(
        oc8051_memory_interface1_n337) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u632 ( .AN(
        oc8051_memory_interface1_n337), .B(
        oc8051_memory_interface1_pcs_source_7_), .Y(
        oc8051_memory_interface1_n385) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u631 ( .AN(
        oc8051_memory_interface1_n337), .B(oc8051_memory_interface1_n579), .Y(
        oc8051_memory_interface1_n375) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u630 ( .A0(
        oc8051_memory_interface1_n4060), .A1(oc8051_memory_interface1_n385), 
        .B0(oc8051_memory_interface1_n3900), .B1(oc8051_memory_interface1_n375), .Y(oc8051_memory_interface1_n578) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u629 ( .A0(
        oc8051_memory_interface1_n359), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n578), .Y(oc8051_memory_interface1_n577)
         );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u628 ( .A0(des2[7]), .A1(
        oc8051_memory_interface1_n575), .B0(oc8051_memory_interface1_n576), 
        .B1(des_acc[7]), .C0(oc8051_memory_interface1_n577), .Y(
        oc8051_memory_interface1_n574) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u627 ( .A(
        oc8051_memory_interface1_n574), .Y(oc8051_memory_interface1_n573) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u626 ( .A(
        oc8051_memory_interface1_n398), .B(oc8051_memory_interface1_n399), .Y(
        oc8051_memory_interface1_n418) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u625 ( .A0(
        oc8051_memory_interface1_pc_buf_15_), .A1(
        oc8051_memory_interface1_n399), .B0(oc8051_memory_interface1_n573), 
        .B1(oc8051_memory_interface1_n418), .C0(oc8051_memory_interface1_n398), 
        .C1(oc8051_memory_interface1_pc_out_15_), .Y(
        oc8051_memory_interface1_n572) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u624 ( .A(
        oc8051_memory_interface1_n572), .Y(oc8051_memory_interface1_n444) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u623 ( .A(
        oc8051_memory_interface1_n400), .Y(oc8051_memory_interface1_n362) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u622 ( .A0(
        oc8051_memory_interface1_op2_buff[6]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[6]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n170)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u621 ( .A(
        oc8051_memory_interface1_n170), .Y(op2_n[6]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u620 ( .A0(
        oc8051_memory_interface1_n3890), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n362), .B1(op2_n[6]), .C0(
        oc8051_memory_interface1_n4050), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n571) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u619 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n541), 
        .B0(oc8051_memory_interface1_n570), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n571), .Y(oc8051_memory_interface1_n539)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u618 ( .A0(
        oc8051_memory_interface1_n418), .A1(oc8051_memory_interface1_n539), 
        .B0(oc8051_memory_interface1_n399), .B1(
        oc8051_memory_interface1_pc_buf_14_), .Y(oc8051_memory_interface1_n537) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u617 ( .A0(n_3_net_), .A1(
        oc8051_memory_interface1_n40), .B0(oc8051_memory_interface1_n537), .Y(
        oc8051_memory_interface1_n445) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u616 ( .A0(
        oc8051_memory_interface1_op2_buff[5]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[5]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n176)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u615 ( .A(
        oc8051_memory_interface1_n176), .Y(op2_n[5]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u614 ( .A0(
        oc8051_memory_interface1_n3880), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n362), .B1(op2_n[5]), .C0(
        oc8051_memory_interface1_n4040), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n535) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u613 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n531), 
        .B0(oc8051_memory_interface1_n533), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n535), .Y(oc8051_memory_interface1_n529)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u612 ( .A0(
        oc8051_memory_interface1_n418), .A1(oc8051_memory_interface1_n529), 
        .B0(oc8051_memory_interface1_n399), .B1(
        oc8051_memory_interface1_pc_buf_13_), .Y(oc8051_memory_interface1_n527) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u611 ( .A0(n_3_net_), .A1(
        oc8051_memory_interface1_n38), .B0(oc8051_memory_interface1_n527), .Y(
        oc8051_memory_interface1_n446) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u610 ( .A0(
        oc8051_memory_interface1_op2_buff[4]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[4]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n181)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u609 ( .A(
        oc8051_memory_interface1_n181), .Y(op2_n[4]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u608 ( .A0(
        oc8051_memory_interface1_n3870), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n362), .B1(op2_n[4]), .C0(
        oc8051_memory_interface1_n4030), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n443) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u607 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n441), 
        .B0(oc8051_memory_interface1_n442), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n443), .Y(oc8051_memory_interface1_n424)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u606 ( .A0(
        oc8051_memory_interface1_n418), .A1(oc8051_memory_interface1_n424), 
        .B0(oc8051_memory_interface1_n399), .B1(
        oc8051_memory_interface1_pc_buf_12_), .Y(oc8051_memory_interface1_n423) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u605 ( .A0(n_3_net_), .A1(
        oc8051_memory_interface1_n39), .B0(oc8051_memory_interface1_n423), .Y(
        oc8051_memory_interface1_n447) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u604 ( .A0(
        oc8051_memory_interface1_op2_buff[3]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[3]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n185)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u603 ( .A(
        oc8051_memory_interface1_n185), .Y(op2_n[3]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u602 ( .A0(
        oc8051_memory_interface1_n3860), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n362), .B1(op2_n[3]), .C0(
        oc8051_memory_interface1_n4020), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n422) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u601 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n420), 
        .B0(oc8051_memory_interface1_n421), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n422), .Y(oc8051_memory_interface1_n419)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u600 ( .A0(
        oc8051_memory_interface1_n418), .A1(oc8051_memory_interface1_n419), 
        .B0(oc8051_memory_interface1_n399), .B1(
        oc8051_memory_interface1_pc_buf_11_), .Y(oc8051_memory_interface1_n417) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u599 ( .A0(n_3_net_), .A1(
        oc8051_memory_interface1_n41), .B0(oc8051_memory_interface1_n417), .Y(
        oc8051_memory_interface1_n448) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u598 ( .A(
        oc8051_memory_interface1_pc_buf_10_), .Y(oc8051_memory_interface1_n327) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u597 ( .A(pc_wr_sel[0]), .Y(
        oc8051_memory_interface1_n363) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u596 ( .A(
        oc8051_memory_interface1_n398), .B(oc8051_memory_interface1_n363), .Y(
        oc8051_memory_interface1_n364) );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u595 ( .A0(
        oc8051_memory_interface1_n364), .A1(pc_wr_sel[2]), .B0(
        oc8051_memory_interface1_n399), .C0(oc8051_memory_interface1_n400), 
        .Y(oc8051_memory_interface1_n367) );
  AND2_X0P5M_A12TS oc8051_memory_interface1_u594 ( .A(
        oc8051_memory_interface1_n399), .B(oc8051_memory_interface1_n367), .Y(
        oc8051_memory_interface1_n369) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u593 ( .AN(
        oc8051_memory_interface1_n367), .B(oc8051_memory_interface1_n398), .Y(
        oc8051_memory_interface1_n370) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u592 ( .A(
        oc8051_memory_interface1_n397), .B(oc8051_memory_interface1_n363), .Y(
        oc8051_memory_interface1_n376) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u591 ( .A0(
        oc8051_memory_interface1_op2_buff[2]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[2]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n188)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u590 ( .A(
        oc8051_memory_interface1_n188), .Y(op2_n[2]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u589 ( .A0(
        oc8051_memory_interface1_n3850), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n376), .B1(op2_n[2]), .C0(
        oc8051_memory_interface1_n4010), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n396) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u588 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n394), 
        .B0(oc8051_memory_interface1_n395), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n396), .Y(oc8051_memory_interface1_n393)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u587 ( .A0(
        oc8051_memory_interface1_n369), .A1(op1_n[7]), .B0(
        oc8051_memory_interface1_n370), .B1(oc8051_memory_interface1_n393), 
        .Y(oc8051_memory_interface1_n392) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u586 ( .A0(
        oc8051_memory_interface1_n327), .A1(oc8051_memory_interface1_n367), 
        .B0(n_3_net_), .B1(oc8051_memory_interface1_n35), .C0(
        oc8051_memory_interface1_n392), .Y(oc8051_memory_interface1_n449) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u585 ( .A(
        oc8051_memory_interface1_pc_buf_9_), .Y(oc8051_memory_interface1_n325)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u584 ( .A0(
        oc8051_memory_interface1_op2_buff[1]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[1]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n202)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u583 ( .A(
        oc8051_memory_interface1_n202), .Y(op2_n[1]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u582 ( .A0(
        oc8051_memory_interface1_n3840), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n376), .B1(op2_n[1]), .C0(
        oc8051_memory_interface1_n4000), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n391) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u581 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n389), 
        .B0(oc8051_memory_interface1_n390), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n391), .Y(oc8051_memory_interface1_n388)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u580 ( .A0(
        oc8051_memory_interface1_n369), .A1(op1_n[6]), .B0(
        oc8051_memory_interface1_n370), .B1(oc8051_memory_interface1_n388), 
        .Y(oc8051_memory_interface1_n387) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u579 ( .A0(
        oc8051_memory_interface1_n325), .A1(oc8051_memory_interface1_n367), 
        .B0(n_3_net_), .B1(oc8051_memory_interface1_n36), .C0(
        oc8051_memory_interface1_n387), .Y(oc8051_memory_interface1_n450) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u578 ( .A(
        oc8051_memory_interface1_pc_buf_8_), .Y(oc8051_memory_interface1_n323)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u577 ( .A0(
        oc8051_memory_interface1_op2_buff[0]), .A1(
        oc8051_memory_interface1_n258), .B0(oc8051_memory_interface1_op2[0]), 
        .B1(oc8051_memory_interface1_n386), .Y(oc8051_memory_interface1_n194)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u576 ( .A(
        oc8051_memory_interface1_n194), .Y(op2_n[0]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u575 ( .A0(
        oc8051_memory_interface1_n3830), .A1(oc8051_memory_interface1_n375), 
        .B0(oc8051_memory_interface1_n376), .B1(op2_n[0]), .C0(
        oc8051_memory_interface1_n3990), .C1(oc8051_memory_interface1_n385), 
        .Y(oc8051_memory_interface1_n374) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u574 ( .A0(
        oc8051_memory_interface1_n366), .A1(oc8051_memory_interface1_n372), 
        .B0(oc8051_memory_interface1_n373), .B1(oc8051_memory_interface1_n365), 
        .C0(oc8051_memory_interface1_n374), .Y(oc8051_memory_interface1_n371)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u573 ( .A0(
        oc8051_memory_interface1_n369), .A1(op1_n[5]), .B0(
        oc8051_memory_interface1_n370), .B1(oc8051_memory_interface1_n371), 
        .Y(oc8051_memory_interface1_n368) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u572 ( .A0(
        oc8051_memory_interface1_n323), .A1(oc8051_memory_interface1_n367), 
        .B0(n_3_net_), .B1(oc8051_memory_interface1_n37), .C0(
        oc8051_memory_interface1_n368), .Y(oc8051_memory_interface1_n451) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u571 ( .A(
        oc8051_memory_interface1_pc_buf_7_), .Y(oc8051_memory_interface1_n320)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u570 ( .A(
        oc8051_memory_interface1_n365), .B(oc8051_memory_interface1_n366), .Y(
        oc8051_memory_interface1_n336) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u569 ( .A(
        oc8051_memory_interface1_n364), .B(oc8051_memory_interface1_n336), .Y(
        oc8051_memory_interface1_n345) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u568 ( .A(
        oc8051_memory_interface1_n362), .B(oc8051_memory_interface1_n363), .Y(
        oc8051_memory_interface1_n339) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u567 ( .A(pc_wr_sel[0]), .B(
        oc8051_memory_interface1_n361), .Y(oc8051_memory_interface1_n340) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u566 ( .A0(
        oc8051_memory_interface1_n359), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n360), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n358) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u565 ( .A0(des_acc[7]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[7]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n358), 
        .Y(oc8051_memory_interface1_n356) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u564 ( .A(n_3_net_), .B(
        oc8051_memory_interface1_n345), .Y(oc8051_memory_interface1_n335) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u563 ( .A(
        oc8051_memory_interface1_pc_out_7_), .Y(oc8051_memory_interface1_n357)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u562 ( .A0(
        oc8051_memory_interface1_n320), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n356), .B1(oc8051_memory_interface1_n335), 
        .C0(n_3_net_), .C1(oc8051_memory_interface1_n357), .Y(
        oc8051_memory_interface1_n452) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u561 ( .A(
        oc8051_memory_interface1_pc_buf_6_), .Y(oc8051_memory_interface1_n318)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u560 ( .A0(
        oc8051_memory_interface1_op3[6]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_6_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[6]), .Y(
        oc8051_memory_interface1_n197) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u559 ( .A0(
        oc8051_memory_interface1_n170), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n355) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u558 ( .A0(des_acc[6]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[6]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n355), 
        .Y(oc8051_memory_interface1_n354) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u557 ( .A0(
        oc8051_memory_interface1_n318), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n354), .B1(oc8051_memory_interface1_n335), 
        .C0(n_3_net_), .C1(oc8051_memory_interface1_n32), .Y(
        oc8051_memory_interface1_n453) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u556 ( .A(
        oc8051_memory_interface1_pc_buf_5_), .Y(oc8051_memory_interface1_n316)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u555 ( .A0(
        oc8051_memory_interface1_op3[5]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_5_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[5]), .Y(
        oc8051_memory_interface1_n198) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u554 ( .A0(
        oc8051_memory_interface1_n176), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n198), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n353) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u553 ( .A0(des_acc[5]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[5]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n353), 
        .Y(oc8051_memory_interface1_n352) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u552 ( .A0(
        oc8051_memory_interface1_n316), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n352), .B1(oc8051_memory_interface1_n335), 
        .C0(n_3_net_), .C1(oc8051_memory_interface1_n33), .Y(
        oc8051_memory_interface1_n454) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u551 ( .A(
        oc8051_memory_interface1_pc_buf_4_), .Y(oc8051_memory_interface1_n314)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u550 ( .A0(
        oc8051_memory_interface1_op3[4]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_4_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[4]), .Y(
        oc8051_memory_interface1_n199) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u549 ( .A0(
        oc8051_memory_interface1_n181), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n199), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n351) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u548 ( .A0(des_acc[4]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[4]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n351), 
        .Y(oc8051_memory_interface1_n350) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u547 ( .A0(
        oc8051_memory_interface1_n314), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n350), .B1(oc8051_memory_interface1_n335), 
        .C0(n_3_net_), .C1(oc8051_memory_interface1_n31), .Y(
        oc8051_memory_interface1_n455) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u546 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .Y(oc8051_memory_interface1_n312)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u545 ( .A0(
        oc8051_memory_interface1_op3[3]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_3_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[3]), .Y(
        oc8051_memory_interface1_n200) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u544 ( .A0(
        oc8051_memory_interface1_n185), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n200), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n349) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u543 ( .A0(des_acc[3]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[3]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n349), 
        .Y(oc8051_memory_interface1_n348) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u542 ( .A0(
        oc8051_memory_interface1_n312), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n348), .B1(oc8051_memory_interface1_n335), 
        .C0(n_3_net_), .C1(oc8051_memory_interface1_n30), .Y(
        oc8051_memory_interface1_n456) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u541 ( .A(
        oc8051_memory_interface1_pc_buf_2_), .Y(oc8051_memory_interface1_n310)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u540 ( .A0(
        oc8051_memory_interface1_op3[2]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_2_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[2]), .Y(
        oc8051_memory_interface1_n201) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u539 ( .A0(
        oc8051_memory_interface1_n188), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n201), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n347) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u538 ( .A0(des_acc[2]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[2]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n347), 
        .Y(oc8051_memory_interface1_n346) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u537 ( .A0(
        oc8051_memory_interface1_n310), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n346), .B1(oc8051_memory_interface1_n335), 
        .C0(n_3_net_), .C1(oc8051_memory_interface1_n29), .Y(
        oc8051_memory_interface1_n457) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u536 ( .A0(
        oc8051_memory_interface1_op3[1]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_1_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[1]), .Y(
        oc8051_memory_interface1_n203) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u535 ( .A0(
        oc8051_memory_interface1_n202), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n203), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n344) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u534 ( .A0(des_acc[1]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[1]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n344), 
        .Y(oc8051_memory_interface1_n343) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u533 ( .A(
        oc8051_memory_interface1_n343), .B(oc8051_memory_interface1_n308), 
        .S0(oc8051_memory_interface1_n335), .Y(oc8051_memory_interface1_n458)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u532 ( .A0(
        oc8051_memory_interface1_op3[0]), .A1(oc8051_memory_interface1_n341), 
        .B0(oc8051_memory_interface1_int_vec_buff_0_), .B1(
        oc8051_memory_interface1_n342), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[0]), .Y(
        oc8051_memory_interface1_n204) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u531 ( .A0(
        oc8051_memory_interface1_n194), .A1(oc8051_memory_interface1_n339), 
        .B0(oc8051_memory_interface1_n204), .B1(oc8051_memory_interface1_n340), 
        .Y(oc8051_memory_interface1_n338) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u530 ( .A0(des_acc[0]), .A1(
        oc8051_memory_interface1_n336), .B0(
        oc8051_memory_interface1_pcs_result[0]), .B1(
        oc8051_memory_interface1_n337), .C0(oc8051_memory_interface1_n338), 
        .Y(oc8051_memory_interface1_n334) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u529 ( .A(
        oc8051_memory_interface1_n334), .B(oc8051_memory_interface1_n304), 
        .S0(oc8051_memory_interface1_n335), .Y(oc8051_memory_interface1_n459)
         );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u528 ( .A(
        oc8051_memory_interface1_int_ack_t), .B(
        oc8051_memory_interface1_pc_wr_r2), .C(oc8051_memory_interface1_n258), 
        .Y(oc8051_memory_interface1_n307) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u527 ( .A(
        oc8051_memory_interface1_n307), .B(oc8051_memory_interface1_pc_wr_r2), 
        .Y(oc8051_memory_interface1_n306) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u526 ( .A(
        oc8051_memory_interface1_n384), .Y(pc[15]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u525 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[15]), .B0(
        oc8051_memory_interface1_n4560), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n333) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u524 ( .B0(
        oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_pc_buf_15_), .A0N(
        oc8051_memory_interface1_n333), .Y(oc8051_memory_interface1_n460) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u523 ( .A(
        oc8051_memory_interface1_n383), .Y(pc[14]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u522 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[14]), .B0(
        oc8051_memory_interface1_n4550), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n332) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u521 ( .B0(
        oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_pc_buf_14_), .A0N(
        oc8051_memory_interface1_n332), .Y(oc8051_memory_interface1_n461) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u520 ( .A(
        oc8051_memory_interface1_n377), .Y(pc[13]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u519 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[13]), .B0(
        oc8051_memory_interface1_n4540), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n331) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u518 ( .B0(
        oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_pc_buf_13_), .A0N(
        oc8051_memory_interface1_n331), .Y(oc8051_memory_interface1_n462) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u516 ( .A(
        oc8051_memory_interface1_n378), .Y(pc[12]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u515 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[12]), .B0(
        oc8051_memory_interface1_n4530), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n330) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u514 ( .B0(
        oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_pc_buf_12_), .A0N(
        oc8051_memory_interface1_n330), .Y(oc8051_memory_interface1_n463) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u513 ( .A(
        oc8051_memory_interface1_n379), .Y(pc[11]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u512 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[11]), .B0(
        oc8051_memory_interface1_n4520), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n329) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u511 ( .B0(
        oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_pc_buf_11_), .A0N(
        oc8051_memory_interface1_n329), .Y(oc8051_memory_interface1_n464) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u510 ( .A(
        oc8051_memory_interface1_n380), .Y(pc[10]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u509 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[10]), .B0(
        oc8051_memory_interface1_n4510), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n328) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u508 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n327), 
        .B0(oc8051_memory_interface1_n328), .Y(oc8051_memory_interface1_n465)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u507 ( .A(
        oc8051_memory_interface1_n381), .Y(pc[9]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u506 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[9]), .B0(
        oc8051_memory_interface1_n4500), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n326) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u505 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n325), 
        .B0(oc8051_memory_interface1_n326), .Y(oc8051_memory_interface1_n466)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u504 ( .A(
        oc8051_memory_interface1_n382), .Y(pc[8]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u503 ( .A0(
        oc8051_memory_interface1_n306), .A1(pc[8]), .B0(
        oc8051_memory_interface1_n4490), .B1(oc8051_memory_interface1_n307), 
        .Y(oc8051_memory_interface1_n324) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u502 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n323), 
        .B0(oc8051_memory_interface1_n324), .Y(oc8051_memory_interface1_n467)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u501 ( .A0(pc[7]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4480), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n321)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u500 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n320), 
        .B0(oc8051_memory_interface1_n321), .Y(oc8051_memory_interface1_n468)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u499 ( .A0(pc[6]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4470), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n319)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u498 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n318), 
        .B0(oc8051_memory_interface1_n319), .Y(oc8051_memory_interface1_n469)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u497 ( .A0(pc[5]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4460), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n317)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u496 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n316), 
        .B0(oc8051_memory_interface1_n317), .Y(oc8051_memory_interface1_n470)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u495 ( .A0(pc[4]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4450), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n315)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u494 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n314), 
        .B0(oc8051_memory_interface1_n315), .Y(oc8051_memory_interface1_n471)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u493 ( .A0(pc[3]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4440), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n313)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u492 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n312), 
        .B0(oc8051_memory_interface1_n313), .Y(oc8051_memory_interface1_n472)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u491 ( .A0(pc[2]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4430), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n311)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u490 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n310), 
        .B0(oc8051_memory_interface1_n311), .Y(oc8051_memory_interface1_n473)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u489 ( .A0(pc[1]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4420), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n309)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u488 ( .A0(
        oc8051_memory_interface1_n301), .A1(oc8051_memory_interface1_n308), 
        .B0(oc8051_memory_interface1_n309), .Y(oc8051_memory_interface1_n474)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u487 ( .A0(pc[0]), .A1(
        oc8051_memory_interface1_n306), .B0(oc8051_memory_interface1_n4410), 
        .B1(oc8051_memory_interface1_n307), .Y(oc8051_memory_interface1_n305)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u486 ( .A0(
        oc8051_memory_interface1_n304), .A1(oc8051_memory_interface1_n301), 
        .B0(oc8051_memory_interface1_n305), .Y(oc8051_memory_interface1_n475)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u485 ( .A(
        oc8051_memory_interface1_op_pos_0_), .B(oc8051_memory_interface1_n4250), .Y(oc8051_memory_interface1_n303) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u484 ( .A(
        oc8051_memory_interface1_n4260), .B(oc8051_memory_interface1_op_pos_1_), .Y(oc8051_memory_interface1_n268) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u483 ( .A(
        oc8051_memory_interface1_n303), .B(oc8051_memory_interface1_n268), .Y(
        oc8051_memory_interface1_n302) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u482 ( .A(
        oc8051_memory_interface1_n302), .B(oc8051_memory_interface1_n301), .Y(
        oc8051_memory_interface1_n300) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u481 ( .A(
        oc8051_memory_interface1_op_pos_1_), .Y(oc8051_memory_interface1_n270)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u480 ( .A(
        oc8051_memory_interface1_n258), .B(oc8051_memory_interface1_n301), .Y(
        oc8051_memory_interface1_n267) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u479 ( .A(
        oc8051_memory_interface1_n267), .Y(oc8051_memory_interface1_n264) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u478 ( .A(
        oc8051_memory_interface1_n300), .B(oc8051_memory_interface1_n270), 
        .S0(oc8051_memory_interface1_n264), .Y(oc8051_memory_interface1_n476)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u477 ( .A(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n259)
         );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u476 ( .A(
        oc8051_memory_interface1_op_pos_0_), .B(oc8051_memory_interface1_n264), 
        .Y(oc8051_memory_interface1_n299) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u475 ( .A(
        oc8051_memory_interface1_n4250), .Y(oc8051_memory_interface1_n260) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u474 ( .A(
        oc8051_memory_interface1_n299), .B(oc8051_memory_interface1_op_pos_0_), 
        .S0(oc8051_memory_interface1_n260), .Y(oc8051_memory_interface1_n298)
         );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u473 ( .A0(
        oc8051_memory_interface1_n259), .A1(oc8051_memory_interface1_n267), 
        .B0(oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_n298), .Y(oc8051_memory_interface1_n477) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u472 ( .A(
        oc8051_memory_interface1_inc_pc), .Y(oc8051_memory_interface1_n266) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u471 ( .A(
        oc8051_memory_interface1_idat_old_31_), .B(
        oc8051_memory_interface1_idat_cur_31_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n478) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u470 ( .A(
        oc8051_memory_interface1_n209), .B(oc8051_memory_interface1_n297), .Y(
        oc8051_memory_interface1_n207) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u469 ( .A(
        oc8051_memory_interface1_n207), .Y(oc8051_memory_interface1_n272) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u468 ( .A(
        oc8051_memory_interface1_n242), .B(oc8051_memory_interface1_n209), .Y(
        oc8051_memory_interface1_n205) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u467 ( .A(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n273) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u466 ( .A0(wbi_dat_i[31]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n296) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u465 ( .A1N(
        oc8051_memory_interface1_idat_cur_31_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n296), 
        .Y(oc8051_memory_interface1_n479) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u464 ( .A(
        oc8051_memory_interface1_idat_old_30_), .B(
        oc8051_memory_interface1_idat_cur_30_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n480) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u463 ( .A0(wbi_dat_i[30]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n295) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u462 ( .A1N(
        oc8051_memory_interface1_idat_cur_30_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n295), 
        .Y(oc8051_memory_interface1_n481) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u461 ( .A(
        oc8051_memory_interface1_idat_old_29_), .B(
        oc8051_memory_interface1_idat_cur_29_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n482) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u460 ( .A0(wbi_dat_i[29]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n294) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u459 ( .A1N(
        oc8051_memory_interface1_idat_cur_29_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n294), 
        .Y(oc8051_memory_interface1_n483) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u458 ( .A(
        oc8051_memory_interface1_idat_old_28_), .B(
        oc8051_memory_interface1_idat_cur_28_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n484) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u457 ( .A0(wbi_dat_i[28]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n293) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u456 ( .A1N(
        oc8051_memory_interface1_idat_cur_28_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n293), 
        .Y(oc8051_memory_interface1_n485) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u455 ( .A(
        oc8051_memory_interface1_idat_old_27_), .B(
        oc8051_memory_interface1_idat_cur_27_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n486) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u454 ( .A0(wbi_dat_i[27]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n292) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u453 ( .A1N(
        oc8051_memory_interface1_idat_cur_27_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n292), 
        .Y(oc8051_memory_interface1_n487) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u452 ( .A(
        oc8051_memory_interface1_idat_old_26_), .B(
        oc8051_memory_interface1_idat_cur_26_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n488) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u451 ( .A0(wbi_dat_i[26]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n291) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u450 ( .A1N(
        oc8051_memory_interface1_idat_cur_26_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n291), 
        .Y(oc8051_memory_interface1_n489) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u449 ( .A(
        oc8051_memory_interface1_idat_old_25_), .B(
        oc8051_memory_interface1_idat_cur_25_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n490) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u448 ( .A0(wbi_dat_i[25]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n290) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u447 ( .A1N(
        oc8051_memory_interface1_idat_cur_25_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n290), 
        .Y(oc8051_memory_interface1_n491) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u446 ( .A(
        oc8051_memory_interface1_idat_old_24_), .B(
        oc8051_memory_interface1_idat_cur_24_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n492) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u445 ( .A0(wbi_dat_i[24]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n289) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u444 ( .A1N(
        oc8051_memory_interface1_idat_cur_24_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n289), 
        .Y(oc8051_memory_interface1_n493) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u443 ( .A(
        oc8051_memory_interface1_idat_old_23_), .B(
        oc8051_memory_interface1_idat_cur_23_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n494) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u442 ( .A0(wbi_dat_i[23]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n288) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u441 ( .A1N(
        oc8051_memory_interface1_idat_cur_23_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n288), 
        .Y(oc8051_memory_interface1_n495) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u440 ( .A(
        oc8051_memory_interface1_idat_old_22_), .B(
        oc8051_memory_interface1_idat_cur_22_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n496) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u439 ( .A0(wbi_dat_i[22]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n287) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u438 ( .A1N(
        oc8051_memory_interface1_idat_cur_22_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n287), 
        .Y(oc8051_memory_interface1_n497) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u437 ( .A(
        oc8051_memory_interface1_idat_old_21_), .B(
        oc8051_memory_interface1_idat_cur_21_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n498) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u436 ( .A0(wbi_dat_i[21]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n286) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u435 ( .A1N(
        oc8051_memory_interface1_idat_cur_21_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n499) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u434 ( .A(
        oc8051_memory_interface1_idat_old_20_), .B(
        oc8051_memory_interface1_idat_cur_20_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n500) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u433 ( .A0(wbi_dat_i[20]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n285) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u432 ( .A1N(
        oc8051_memory_interface1_idat_cur_20_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n285), 
        .Y(oc8051_memory_interface1_n501) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u431 ( .A(
        oc8051_memory_interface1_idat_old_19_), .B(
        oc8051_memory_interface1_idat_cur_19_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n502) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u430 ( .A0(wbi_dat_i[19]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n284) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u429 ( .A1N(
        oc8051_memory_interface1_idat_cur_19_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n284), 
        .Y(oc8051_memory_interface1_n503) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u428 ( .A(
        oc8051_memory_interface1_idat_old_18_), .B(
        oc8051_memory_interface1_idat_cur_18_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n504) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u427 ( .A0(wbi_dat_i[18]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n283) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u426 ( .A1N(
        oc8051_memory_interface1_idat_cur_18_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n283), 
        .Y(oc8051_memory_interface1_n505) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u425 ( .A(
        oc8051_memory_interface1_idat_old_17_), .B(
        oc8051_memory_interface1_idat_cur_17_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n506) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u424 ( .A0(wbi_dat_i[17]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n282) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u423 ( .A1N(
        oc8051_memory_interface1_idat_cur_17_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n282), 
        .Y(oc8051_memory_interface1_n507) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u422 ( .A(
        oc8051_memory_interface1_idat_old_16_), .B(
        oc8051_memory_interface1_idat_cur_16_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n508) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u421 ( .A0(wbi_dat_i[16]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n281) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u420 ( .A1N(
        oc8051_memory_interface1_idat_cur_16_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n281), 
        .Y(oc8051_memory_interface1_n509) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u419 ( .A(
        oc8051_memory_interface1_idat_old_15_), .B(
        oc8051_memory_interface1_idat_cur_15_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n510) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u418 ( .A0(wbi_dat_i[15]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n280) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u417 ( .A1N(
        oc8051_memory_interface1_idat_cur_15_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n280), 
        .Y(oc8051_memory_interface1_n511) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u416 ( .A(
        oc8051_memory_interface1_idat_old_14_), .B(
        oc8051_memory_interface1_idat_cur_14_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n512) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u415 ( .A0(wbi_dat_i[14]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n279) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u414 ( .A1N(
        oc8051_memory_interface1_idat_cur_14_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n279), 
        .Y(oc8051_memory_interface1_n513) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u413 ( .A(
        oc8051_memory_interface1_idat_old_13_), .B(
        oc8051_memory_interface1_idat_cur_13_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n514) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u412 ( .A0(wbi_dat_i[13]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n278) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u411 ( .A1N(
        oc8051_memory_interface1_idat_cur_13_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n278), 
        .Y(oc8051_memory_interface1_n515) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u410 ( .A(
        oc8051_memory_interface1_idat_old_12_), .B(
        oc8051_memory_interface1_idat_cur_12_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n516) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u409 ( .A0(wbi_dat_i[12]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n277) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u408 ( .A1N(
        oc8051_memory_interface1_idat_cur_12_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n277), 
        .Y(oc8051_memory_interface1_n517) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u407 ( .A(
        oc8051_memory_interface1_idat_old_11_), .B(
        oc8051_memory_interface1_idat_cur_11_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n518) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u406 ( .A0(wbi_dat_i[11]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n276) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u405 ( .A1N(
        oc8051_memory_interface1_idat_cur_11_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n276), 
        .Y(oc8051_memory_interface1_n519) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u404 ( .A(
        oc8051_memory_interface1_idat_old_10_), .B(
        oc8051_memory_interface1_idat_cur_10_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n520) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u403 ( .A0(wbi_dat_i[10]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n275) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u402 ( .A1N(
        oc8051_memory_interface1_idat_cur_10_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n275), 
        .Y(oc8051_memory_interface1_n521) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u401 ( .A(
        oc8051_memory_interface1_idat_old_9_), .B(
        oc8051_memory_interface1_idat_cur_9_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n522) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u400 ( .A0(wbi_dat_i[9]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n274) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u399 ( .A1N(
        oc8051_memory_interface1_idat_cur_9_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n274), 
        .Y(oc8051_memory_interface1_n523) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u398 ( .A(
        oc8051_memory_interface1_idat_old_8_), .B(
        oc8051_memory_interface1_idat_cur_8_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n524) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u397 ( .A0(wbi_dat_i[8]), .A1(
        oc8051_memory_interface1_n272), .B0(n_logic0_), .B1(
        oc8051_memory_interface1_n273), .Y(oc8051_memory_interface1_n271) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u396 ( .A1N(
        oc8051_memory_interface1_idat_cur_8_), .A0(
        oc8051_memory_interface1_n209), .B0(oc8051_memory_interface1_n271), 
        .Y(oc8051_memory_interface1_n525) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u395 ( .A(
        oc8051_memory_interface1_idat_old_7_), .B(
        oc8051_memory_interface1_idat_cur_7_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n526) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u394 ( .A(
        oc8051_memory_interface1_idat_old_6_), .B(
        oc8051_memory_interface1_idat_cur_6_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n528) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u393 ( .A(
        oc8051_memory_interface1_idat_old_5_), .B(
        oc8051_memory_interface1_idat_cur_5_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n530) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u392 ( .A(
        oc8051_memory_interface1_idat_old_4_), .B(
        oc8051_memory_interface1_idat_cur_4_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n532) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u391 ( .A(
        oc8051_memory_interface1_idat_old_3_), .B(
        oc8051_memory_interface1_idat_cur_3_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n534) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u390 ( .A(
        oc8051_memory_interface1_idat_old_2_), .B(
        oc8051_memory_interface1_idat_cur_2_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n536) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u389 ( .A(
        oc8051_memory_interface1_idat_old_1_), .B(
        oc8051_memory_interface1_idat_cur_1_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n538) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u388 ( .A(
        oc8051_memory_interface1_idat_old_0_), .B(
        oc8051_memory_interface1_idat_cur_0_), .S0(
        oc8051_memory_interface1_n209), .Y(oc8051_memory_interface1_n540) );
  AND3_X0P5M_A12TS oc8051_memory_interface1_u387 ( .A(
        oc8051_memory_interface1_op_pos_2_), .B(oc8051_memory_interface1_n270), 
        .C(oc8051_memory_interface1_n4260), .Y(oc8051_memory_interface1_n269)
         );
  AOI31_X0P5M_A12TS oc8051_memory_interface1_u386 ( .A0(
        oc8051_memory_interface1_n267), .A1(oc8051_memory_interface1_n266), 
        .A2(oc8051_memory_interface1_n268), .B0(oc8051_memory_interface1_n269), 
        .Y(oc8051_memory_interface1_n261) );
  AOI31_X0P5M_A12TS oc8051_memory_interface1_u385 ( .A0(
        oc8051_memory_interface1_op_pos_1_), .A1(oc8051_memory_interface1_n266), .A2(oc8051_memory_interface1_n4260), .B0(oc8051_memory_interface1_pc_wr_r2), 
        .Y(oc8051_memory_interface1_n265) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u384 ( .A(
        oc8051_memory_interface1_n265), .Y(oc8051_memory_interface1_n263) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u383 ( .A(
        oc8051_memory_interface1_n263), .B(oc8051_memory_interface1_op_pos_2_), 
        .S0(oc8051_memory_interface1_n264), .Y(oc8051_memory_interface1_n262)
         );
  OAI31_X0P5M_A12TS oc8051_memory_interface1_u382 ( .A0(
        oc8051_memory_interface1_n259), .A1(oc8051_memory_interface1_n260), 
        .A2(oc8051_memory_interface1_n261), .B0(oc8051_memory_interface1_n262), 
        .Y(oc8051_memory_interface1_n542) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u381 ( .A(
        oc8051_memory_interface1_n258), .B(oc8051_memory_interface1_pc_wr_r2), 
        .C(oc8051_memory_interface1_n243), .Y(oc8051_memory_interface1_n256)
         );
  OAI21B_X0P5M_A12TS oc8051_memory_interface1_u380 ( .A0(
        oc8051_memory_interface1_n256), .A1(oc8051_memory_interface1_n257), 
        .B0N(intr), .Y(oc8051_memory_interface1_n543) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u379 ( .A(wbd_ack_i), .B(
        mem_act[1]), .Y(oc8051_memory_interface1_n245) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u378 ( .A(
        oc8051_memory_interface1_n255), .B(wbd_ack_i), .Y(
        oc8051_memory_interface1_n247) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u377 ( .A0(dptr_lo[0]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[0]), .Y(oc8051_memory_interface1_n254) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u376 ( .B0(wbd_adr_o[0]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n254), .Y(
        oc8051_memory_interface1_n544) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u375 ( .A0(dptr_lo[1]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[1]), .Y(oc8051_memory_interface1_n253) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u374 ( .B0(wbd_adr_o[1]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n253), .Y(
        oc8051_memory_interface1_n545) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u373 ( .A0(dptr_lo[2]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[2]), .Y(oc8051_memory_interface1_n252) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u372 ( .B0(wbd_adr_o[2]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n252), .Y(
        oc8051_memory_interface1_n546) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u371 ( .A0(dptr_lo[3]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[3]), .Y(oc8051_memory_interface1_n251) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u370 ( .B0(wbd_adr_o[3]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n251), .Y(
        oc8051_memory_interface1_n547) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u369 ( .A0(dptr_lo[4]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[4]), .Y(oc8051_memory_interface1_n250) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u368 ( .B0(wbd_adr_o[4]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n250), .Y(
        oc8051_memory_interface1_n548) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u367 ( .A0(dptr_lo[5]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[5]), .Y(oc8051_memory_interface1_n249) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u366 ( .B0(wbd_adr_o[5]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n249), .Y(
        oc8051_memory_interface1_n549) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u365 ( .A0(dptr_lo[6]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[6]), .Y(oc8051_memory_interface1_n248) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u364 ( .B0(wbd_adr_o[6]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n248), .Y(
        oc8051_memory_interface1_n550) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u363 ( .A0(dptr_lo[7]), .A1(
        oc8051_memory_interface1_n245), .B0(oc8051_memory_interface1_n247), 
        .B1(ri[7]), .Y(oc8051_memory_interface1_n246) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u362 ( .B0(wbd_adr_o[7]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n246), .Y(
        oc8051_memory_interface1_n551) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u361 ( .A0(wbd_adr_o[8]), .A1(
        wbd_ack_i), .B0(dptr_hi[0]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n552) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u360 ( .A0(wbd_adr_o[9]), .A1(
        wbd_ack_i), .B0(dptr_hi[1]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n553) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u359 ( .A0(wbd_adr_o[10]), .A1(
        wbd_ack_i), .B0(dptr_hi[2]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n554) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u358 ( .A0(wbd_adr_o[11]), .A1(
        wbd_ack_i), .B0(dptr_hi[3]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n555) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u357 ( .A0(wbd_adr_o[12]), .A1(
        wbd_ack_i), .B0(dptr_hi[4]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n556) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u356 ( .A0(wbd_adr_o[13]), .A1(
        wbd_ack_i), .B0(dptr_hi[5]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n557) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u355 ( .A0(wbd_adr_o[14]), .A1(
        wbd_ack_i), .B0(dptr_hi[6]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n558) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u354 ( .A0(wbd_adr_o[15]), .A1(
        wbd_ack_i), .B0(dptr_hi[7]), .B1(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n559) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u353 ( .A0(wbd_dat_o[0]), .A1(
        wbd_ack_i), .B0(acc[0]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n560) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u352 ( .A0(wbd_dat_o[1]), .A1(
        wbd_ack_i), .B0(acc[1]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n561) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u351 ( .A0(wbd_dat_o[2]), .A1(
        wbd_ack_i), .B0(acc[2]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n562) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u350 ( .A0(wbd_dat_o[3]), .A1(
        wbd_ack_i), .B0(acc[3]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n563) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u349 ( .A0(wbd_dat_o[4]), .A1(
        wbd_ack_i), .B0(acc[4]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n564) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u348 ( .A0(wbd_dat_o[5]), .A1(
        wbd_ack_i), .B0(acc[5]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n565) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u347 ( .A0(wbd_dat_o[6]), .A1(
        wbd_ack_i), .B0(acc[6]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n566) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u346 ( .A0(wbd_dat_o[7]), .A1(
        wbd_ack_i), .B0(acc[7]), .B1(oc8051_memory_interface1_n1290), .Y(
        oc8051_memory_interface1_n567) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u345 ( .B0(
        oc8051_memory_interface1_istb_t), .B1(
        oc8051_memory_interface1_imem_wait), .A0N(
        oc8051_memory_interface1_n244), .Y(oc8051_memory_interface1_n568) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u344 ( .B0(
        oc8051_memory_interface1_n243), .B1(oc8051_memory_interface1_imem_wait), .A0N(oc8051_memory_interface1_n244), .Y(oc8051_memory_interface1_n569) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u343 ( .A(wbd_ack_i), .Y(
        oc8051_memory_interface1_n691) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u342 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n229) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u341 ( .A(
        oc8051_memory_interface1_istb_t), .B(oc8051_memory_interface1_n242), 
        .Y(oc8051_memory_interface1_n232) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u340 ( .A(wbi_dat_i[7]), .Y(
        oc8051_memory_interface1_n230) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u339 ( .A(
        oc8051_memory_interface1_cdata_7_), .Y(oc8051_memory_interface1_n241)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u338 ( .A0(
        oc8051_memory_interface1_n229), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n230), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n241), .Y(oc8051_memory_interface1_n682) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u337 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n226) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u336 ( .A(wbi_dat_i[6]), .Y(
        oc8051_memory_interface1_n227) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u335 ( .A(
        oc8051_memory_interface1_cdata_6_), .Y(oc8051_memory_interface1_n240)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u334 ( .A0(
        oc8051_memory_interface1_n226), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n227), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n240), .Y(oc8051_memory_interface1_n681) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u333 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n223) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u332 ( .A(wbi_dat_i[5]), .Y(
        oc8051_memory_interface1_n224) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u331 ( .A(
        oc8051_memory_interface1_cdata_5_), .Y(oc8051_memory_interface1_n239)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u330 ( .A0(
        oc8051_memory_interface1_n223), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n224), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n239), .Y(oc8051_memory_interface1_n680) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u329 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n220) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u328 ( .A(wbi_dat_i[4]), .Y(
        oc8051_memory_interface1_n221) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u327 ( .A(
        oc8051_memory_interface1_cdata_4_), .Y(oc8051_memory_interface1_n238)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u326 ( .A0(
        oc8051_memory_interface1_n220), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n221), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n238), .Y(oc8051_memory_interface1_n679) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u325 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n217) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u324 ( .A(wbi_dat_i[3]), .Y(
        oc8051_memory_interface1_n218) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u323 ( .A(
        oc8051_memory_interface1_cdata_3_), .Y(oc8051_memory_interface1_n237)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u322 ( .A0(
        oc8051_memory_interface1_n217), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n218), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n237), .Y(oc8051_memory_interface1_n678) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u321 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n214) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u320 ( .A(wbi_dat_i[2]), .Y(
        oc8051_memory_interface1_n215) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u319 ( .A(
        oc8051_memory_interface1_cdata_2_), .Y(oc8051_memory_interface1_n236)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u318 ( .A0(
        oc8051_memory_interface1_n214), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n215), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n236), .Y(oc8051_memory_interface1_n677) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u317 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n211) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u316 ( .A(wbi_dat_i[1]), .Y(
        oc8051_memory_interface1_n212) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u315 ( .A(
        oc8051_memory_interface1_cdata_1_), .Y(oc8051_memory_interface1_n235)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u314 ( .A0(
        oc8051_memory_interface1_n211), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n212), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n235), .Y(oc8051_memory_interface1_n676) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u313 ( .A(n_logic0_), .Y(
        oc8051_memory_interface1_n206) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u312 ( .A(wbi_dat_i[0]), .Y(
        oc8051_memory_interface1_n208) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u311 ( .A(
        oc8051_memory_interface1_cdata_0_), .Y(oc8051_memory_interface1_n234)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u310 ( .A0(
        oc8051_memory_interface1_n206), .A1(oc8051_memory_interface1_n232), 
        .B0(oc8051_memory_interface1_n208), .B1(oc8051_memory_interface1_n233), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n234), .Y(oc8051_memory_interface1_n675) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u309 ( .A(
        oc8051_memory_interface1_idat_cur_7_), .Y(
        oc8051_memory_interface1_n231) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u308 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n229), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n230), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n231), 
        .Y(oc8051_memory_interface1_n673) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u307 ( .A(
        oc8051_memory_interface1_idat_cur_6_), .Y(
        oc8051_memory_interface1_n228) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u306 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n226), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n227), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n228), 
        .Y(oc8051_memory_interface1_n672) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u305 ( .A(
        oc8051_memory_interface1_idat_cur_5_), .Y(
        oc8051_memory_interface1_n225) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u304 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n223), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n224), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n225), 
        .Y(oc8051_memory_interface1_n671) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u303 ( .A(
        oc8051_memory_interface1_idat_cur_4_), .Y(
        oc8051_memory_interface1_n222) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u302 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n220), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n221), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n222), 
        .Y(oc8051_memory_interface1_n670) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u301 ( .A(
        oc8051_memory_interface1_idat_cur_3_), .Y(
        oc8051_memory_interface1_n219) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u300 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n217), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n218), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n219), 
        .Y(oc8051_memory_interface1_n669) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u299 ( .A(
        oc8051_memory_interface1_idat_cur_2_), .Y(
        oc8051_memory_interface1_n216) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u298 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n214), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n215), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n216), 
        .Y(oc8051_memory_interface1_n668) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u297 ( .A(
        oc8051_memory_interface1_idat_cur_1_), .Y(
        oc8051_memory_interface1_n213) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u296 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n211), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n212), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n213), 
        .Y(oc8051_memory_interface1_n667) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u295 ( .A(
        oc8051_memory_interface1_idat_cur_0_), .Y(
        oc8051_memory_interface1_n210) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u294 ( .A0(
        oc8051_memory_interface1_n205), .A1(oc8051_memory_interface1_n206), 
        .B0(oc8051_memory_interface1_n207), .B1(oc8051_memory_interface1_n208), 
        .C0(oc8051_memory_interface1_n209), .C1(oc8051_memory_interface1_n210), 
        .Y(oc8051_memory_interface1_n666) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u293 ( .A(
        oc8051_memory_interface1_n204), .Y(op3_n[0]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u292 ( .A(
        oc8051_memory_interface1_n203), .Y(op3_n[1]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u291 ( .A(
        oc8051_memory_interface1_n201), .Y(op3_n[2]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u290 ( .A(
        oc8051_memory_interface1_n200), .Y(op3_n[3]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u289 ( .A(
        oc8051_memory_interface1_n199), .Y(op3_n[4]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u288 ( .A(
        oc8051_memory_interface1_n198), .Y(op3_n[5]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u287 ( .A(
        oc8051_memory_interface1_n197), .Y(op3_n[6]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u286 ( .A(
        oc8051_memory_interface1_n194), .B(oc8051_memory_interface1_n204), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_0_) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u285 ( .A(
        oc8051_memory_interface1_n202), .B(oc8051_memory_interface1_n203), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_1_) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u284 ( .A(
        oc8051_memory_interface1_n188), .B(oc8051_memory_interface1_n201), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_2_) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u283 ( .A(
        oc8051_memory_interface1_n185), .B(oc8051_memory_interface1_n200), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_3_) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u282 ( .A(
        oc8051_memory_interface1_n181), .B(oc8051_memory_interface1_n199), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_4_) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u281 ( .A(
        oc8051_memory_interface1_n176), .B(oc8051_memory_interface1_n198), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_5_) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u280 ( .A(
        oc8051_memory_interface1_n170), .B(oc8051_memory_interface1_n197), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_pcs_source_6_) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u279 ( .A(ram_rd_sel[2]), .Y(
        oc8051_memory_interface1_n166) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u278 ( .A(
        oc8051_memory_interface1_n180), .B(oc8051_memory_interface1_n166), .C(
        ram_rd_sel[1]), .Y(oc8051_memory_interface1_n171) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u277 ( .A(ram_rd_sel[1]), .Y(
        oc8051_memory_interface1_n172) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u276 ( .AN(
        oc8051_memory_interface1_n810), .B(oc8051_memory_interface1_n172), .Y(
        oc8051_memory_interface1_n168) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u275 ( .A(sp[0]), .B(
        oc8051_memory_interface1_n168), .Y(oc8051_memory_interface1_n195) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u274 ( .A(
        oc8051_memory_interface1_n810), .B(oc8051_memory_interface1_n172), .Y(
        oc8051_memory_interface1_n164) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u273 ( .A(
        oc8051_memory_interface1_n164), .Y(oc8051_memory_interface1_n174) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u272 ( .A(ram_rd_sel[1]), .B(
        ram_rd_sel[2]), .C(ram_rd_sel[0]), .Y(oc8051_memory_interface1_n184)
         );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u271 ( .A0(ram_rd_sel[0]), .A1(
        oc8051_memory_interface1_n172), .A2(ram_rd_sel[2]), .B0(ri[1]), .B1(
        oc8051_memory_interface1_n174), .Y(oc8051_memory_interface1_n191) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u270 ( .A(op1_cur[1]), .B(
        oc8051_memory_interface1_n184), .Y(oc8051_memory_interface1_n192) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u269 ( .A(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n169) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u268 ( .A0(sp[1]), .A1(
        oc8051_memory_interface1_n168), .B0(oc8051_memory_interface1_n169), 
        .B1(op2_n[1]), .Y(oc8051_memory_interface1_n193) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u267 ( .A(sp[2]), .B(
        oc8051_memory_interface1_n168), .Y(oc8051_memory_interface1_n189) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u266 ( .A(sp[3]), .B(
        oc8051_memory_interface1_n168), .Y(oc8051_memory_interface1_n186) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u265 ( .A0(ri[3]), .A1(
        oc8051_memory_interface1_n174), .B0(bank_sel[0]), .B1(
        oc8051_memory_interface1_n184), .Y(oc8051_memory_interface1_n187) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u264 ( .A0(
        oc8051_memory_interface1_n185), .A1(oc8051_memory_interface1_n171), 
        .B0(oc8051_memory_interface1_n186), .C0(oc8051_memory_interface1_n187), 
        .Y(rd_addr[3]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u263 ( .A(sp[4]), .B(
        oc8051_memory_interface1_n168), .Y(oc8051_memory_interface1_n182) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u262 ( .A(
        oc8051_memory_interface1_n166), .B(ram_rd_sel[0]), .Y(
        oc8051_memory_interface1_n175) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u261 ( .A0(bank_sel[1]), .A1(
        oc8051_memory_interface1_n184), .B0(ri[4]), .B1(
        oc8051_memory_interface1_n174), .C0(oc8051_memory_interface1_n175), 
        .Y(oc8051_memory_interface1_n183) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u260 ( .A0(
        oc8051_memory_interface1_n181), .A1(oc8051_memory_interface1_n171), 
        .B0(oc8051_memory_interface1_n182), .C0(oc8051_memory_interface1_n183), 
        .Y(rd_addr[4]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u259 ( .A(
        oc8051_memory_interface1_n180), .B(oc8051_memory_interface1_n166), .Y(
        oc8051_memory_interface1_n179) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u258 ( .A(
        oc8051_memory_interface1_n175), .B(oc8051_memory_interface1_n179), 
        .S0(ram_rd_sel[1]), .Y(oc8051_memory_interface1_n177) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u257 ( .A0(ri[5]), .A1(
        oc8051_memory_interface1_n174), .B0(sp[5]), .B1(
        oc8051_memory_interface1_n168), .Y(oc8051_memory_interface1_n178) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u256 ( .A0(
        oc8051_memory_interface1_n176), .A1(oc8051_memory_interface1_n171), 
        .B0(oc8051_memory_interface1_n177), .C0(oc8051_memory_interface1_n178), 
        .Y(rd_addr[5]) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u255 ( .A0(sp[6]), .A1(
        oc8051_memory_interface1_n168), .B0(ri[6]), .B1(
        oc8051_memory_interface1_n174), .C0(oc8051_memory_interface1_n175), 
        .Y(oc8051_memory_interface1_n173) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u254 ( .A0(
        oc8051_memory_interface1_n170), .A1(oc8051_memory_interface1_n171), 
        .B0(oc8051_memory_interface1_n172), .B1(oc8051_memory_interface1_n166), 
        .C0(oc8051_memory_interface1_n173), .Y(rd_addr[6]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u253 ( .A(ri[7]), .Y(
        oc8051_memory_interface1_n165) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u252 ( .A0(sp[7]), .A1(
        oc8051_memory_interface1_n168), .B0(oc8051_memory_interface1_n169), 
        .B1(op2_n[7]), .Y(oc8051_memory_interface1_n167) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u251 ( .A(
        oc8051_memory_interface1_n153), .B(ram_wr_sel[0]), .Y(
        oc8051_memory_interface1_n146) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u250 ( .A(ram_wr_sel[0]), .B(
        ram_wr_sel[1]), .Y(oc8051_memory_interface1_n154) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u249 ( .A0(
        oc8051_memory_interface1_ri_r[0]), .A1(oc8051_memory_interface1_n146), 
        .B0(oc8051_memory_interface1_rn_r[0]), .B1(
        oc8051_memory_interface1_n154), .Y(oc8051_memory_interface1_n161) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u248 ( .A(ram_wr_sel[0]), .Y(
        oc8051_memory_interface1_n163) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u247 ( .A(ram_wr_sel[1]), .B(
        ram_wr_sel[2]), .C(oc8051_memory_interface1_n163), .Y(
        oc8051_memory_interface1_n145) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u246 ( .AN(ram_wr_sel[2]), .B(
        ram_wr_sel[1]), .Y(oc8051_memory_interface1_n143) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u245 ( .AN(wr_ind), .B(
        oc8051_memory_interface1_n163), .Y(oc8051_memory_interface1_n142) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u244 ( .A0(
        oc8051_memory_interface1_ri_r[1]), .A1(oc8051_memory_interface1_n146), 
        .B0(oc8051_memory_interface1_rn_r[1]), .B1(
        oc8051_memory_interface1_n154), .Y(oc8051_memory_interface1_n159) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u243 ( .A0(
        oc8051_memory_interface1_ri_r[2]), .A1(oc8051_memory_interface1_n146), 
        .B0(oc8051_memory_interface1_rn_r[2]), .B1(
        oc8051_memory_interface1_n154), .Y(oc8051_memory_interface1_n157) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u242 ( .A0(
        oc8051_memory_interface1_ri_r[3]), .A1(oc8051_memory_interface1_n146), 
        .B0(oc8051_memory_interface1_rn_r[3]), .B1(
        oc8051_memory_interface1_n154), .Y(oc8051_memory_interface1_n155) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u241 ( .A0(
        oc8051_memory_interface1_imm_r[3]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_imm2_r[3]), .B1(
        oc8051_memory_interface1_n143), .C0(sp_w[3]), .C1(
        oc8051_memory_interface1_n142), .Y(oc8051_memory_interface1_n156) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u240 ( .A(
        oc8051_memory_interface1_n155), .B(oc8051_memory_interface1_n156), .Y(
        wr_addr[3]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u239 ( .A0(
        oc8051_memory_interface1_rn_r[4]), .A1(oc8051_memory_interface1_n154), 
        .B0(oc8051_memory_interface1_imm_r[4]), .B1(
        oc8051_memory_interface1_n145), .C0(oc8051_memory_interface1_ri_r[4]), 
        .C1(oc8051_memory_interface1_n146), .Y(oc8051_memory_interface1_n151)
         );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u238 ( .AN(ram_wr_sel[2]), .B(
        oc8051_memory_interface1_n153), .Y(oc8051_memory_interface1_n144) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u237 ( .A0(sp_w[4]), .A1(
        oc8051_memory_interface1_n142), .B0(oc8051_memory_interface1_imm2_r[4]), .B1(oc8051_memory_interface1_n143), .C0(oc8051_memory_interface1_n144), .Y(
        oc8051_memory_interface1_n152) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u236 ( .A(
        oc8051_memory_interface1_n151), .B(oc8051_memory_interface1_n152), .Y(
        wr_addr[4]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u235 ( .A0(
        oc8051_memory_interface1_imm_r[5]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_ri_r[5]), .B1(
        oc8051_memory_interface1_n146), .Y(oc8051_memory_interface1_n149) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u234 ( .A0(sp_w[5]), .A1(
        oc8051_memory_interface1_n142), .B0(oc8051_memory_interface1_imm2_r[5]), .B1(oc8051_memory_interface1_n143), .C0(oc8051_memory_interface1_n144), .Y(
        oc8051_memory_interface1_n150) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u233 ( .A(
        oc8051_memory_interface1_n149), .B(oc8051_memory_interface1_n150), .Y(
        wr_addr[5]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u232 ( .A0(
        oc8051_memory_interface1_imm_r[6]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_ri_r[6]), .B1(
        oc8051_memory_interface1_n146), .Y(oc8051_memory_interface1_n147) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u231 ( .A0(sp_w[6]), .A1(
        oc8051_memory_interface1_n142), .B0(oc8051_memory_interface1_imm2_r[6]), .B1(oc8051_memory_interface1_n143), .C0(oc8051_memory_interface1_n144), .Y(
        oc8051_memory_interface1_n148) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u230 ( .A(
        oc8051_memory_interface1_n147), .B(oc8051_memory_interface1_n148), .Y(
        wr_addr[6]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u229 ( .A0(
        oc8051_memory_interface1_imm_r[7]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_ri_r[7]), .B1(
        oc8051_memory_interface1_n146), .Y(oc8051_memory_interface1_n140) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u228 ( .A0(sp_w[7]), .A1(
        oc8051_memory_interface1_n142), .B0(oc8051_memory_interface1_imm2_r[7]), .B1(oc8051_memory_interface1_n143), .C0(oc8051_memory_interface1_n144), .Y(
        oc8051_memory_interface1_n141) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u227 ( .A(
        oc8051_memory_interface1_n140), .B(oc8051_memory_interface1_n141), .Y(
        wr_addr[7]) );
  AND2_X1M_A12TS oc8051_memory_interface1_u226 ( .A(
        oc8051_memory_interface1_n63), .B(oc8051_memory_interface1_pc_buf_10_), 
        .Y(oc8051_memory_interface1_n64) );
  AND2_X1M_A12TS oc8051_memory_interface1_u225 ( .A(
        oc8051_memory_interface1_n62), .B(oc8051_memory_interface1_pc_buf_9_), 
        .Y(oc8051_memory_interface1_n63) );
  AND2_X1M_A12TS oc8051_memory_interface1_u224 ( .A(
        oc8051_memory_interface1_n61), .B(oc8051_memory_interface1_pc_buf_8_), 
        .Y(oc8051_memory_interface1_n62) );
  AND2_X1M_A12TS oc8051_memory_interface1_u223 ( .A(
        oc8051_memory_interface1_n60), .B(oc8051_memory_interface1_pc_buf_7_), 
        .Y(oc8051_memory_interface1_n61) );
  AND2_X1M_A12TS oc8051_memory_interface1_u222 ( .A(
        oc8051_memory_interface1_n59), .B(oc8051_memory_interface1_pc_buf_6_), 
        .Y(oc8051_memory_interface1_n60) );
  AND2_X1M_A12TS oc8051_memory_interface1_u221 ( .A(
        oc8051_memory_interface1_n58), .B(oc8051_memory_interface1_pc_buf_5_), 
        .Y(oc8051_memory_interface1_n59) );
  AND2_X1M_A12TS oc8051_memory_interface1_u220 ( .A(
        oc8051_memory_interface1_n57), .B(oc8051_memory_interface1_pc_buf_4_), 
        .Y(oc8051_memory_interface1_n58) );
  AND2_X1M_A12TS oc8051_memory_interface1_u219 ( .A(
        oc8051_memory_interface1_n42), .B(oc8051_memory_interface1_pc_buf_3_), 
        .Y(oc8051_memory_interface1_n57) );
  AND2_X1M_A12TS oc8051_memory_interface1_u218 ( .A(
        oc8051_memory_interface1_n55), .B(oc8051_memory_interface1_pc_buf_13_), 
        .Y(oc8051_memory_interface1_n56) );
  AND2_X1M_A12TS oc8051_memory_interface1_u217 ( .A(
        oc8051_memory_interface1_n54), .B(oc8051_memory_interface1_pc_buf_12_), 
        .Y(oc8051_memory_interface1_n55) );
  AND2_X1M_A12TS oc8051_memory_interface1_u216 ( .A(
        oc8051_memory_interface1_n64), .B(oc8051_memory_interface1_pc_buf_11_), 
        .Y(oc8051_memory_interface1_n54) );
  AND2_X1M_A12TS oc8051_memory_interface1_u215 ( .A(
        oc8051_memory_interface1_pc_buf_10_), .B(oc8051_memory_interface1_n52), 
        .Y(oc8051_memory_interface1_n53) );
  AND2_X1M_A12TS oc8051_memory_interface1_u214 ( .A(
        oc8051_memory_interface1_pc_buf_9_), .B(oc8051_memory_interface1_n51), 
        .Y(oc8051_memory_interface1_n52) );
  AND2_X1M_A12TS oc8051_memory_interface1_u213 ( .A(
        oc8051_memory_interface1_pc_buf_8_), .B(oc8051_memory_interface1_n50), 
        .Y(oc8051_memory_interface1_n51) );
  AND2_X1M_A12TS oc8051_memory_interface1_u212 ( .A(
        oc8051_memory_interface1_pc_buf_7_), .B(oc8051_memory_interface1_n49), 
        .Y(oc8051_memory_interface1_n50) );
  AND2_X1M_A12TS oc8051_memory_interface1_u211 ( .A(
        oc8051_memory_interface1_pc_buf_6_), .B(oc8051_memory_interface1_n48), 
        .Y(oc8051_memory_interface1_n49) );
  AND2_X1M_A12TS oc8051_memory_interface1_u210 ( .A(
        oc8051_memory_interface1_pc_buf_5_), .B(oc8051_memory_interface1_n47), 
        .Y(oc8051_memory_interface1_n48) );
  AND2_X1M_A12TS oc8051_memory_interface1_u209 ( .A(
        oc8051_memory_interface1_pc_buf_4_), .B(oc8051_memory_interface1_n43), 
        .Y(oc8051_memory_interface1_n47) );
  AND2_X1M_A12TS oc8051_memory_interface1_u208 ( .A(
        oc8051_memory_interface1_pc_buf_13_), .B(oc8051_memory_interface1_n45), 
        .Y(oc8051_memory_interface1_n46) );
  AND2_X1M_A12TS oc8051_memory_interface1_u207 ( .A(
        oc8051_memory_interface1_pc_buf_12_), .B(oc8051_memory_interface1_n44), 
        .Y(oc8051_memory_interface1_n45) );
  AND2_X1M_A12TS oc8051_memory_interface1_u206 ( .A(
        oc8051_memory_interface1_pc_buf_11_), .B(oc8051_memory_interface1_n53), 
        .Y(oc8051_memory_interface1_n44) );
  AND2_X1M_A12TS oc8051_memory_interface1_u205 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .B(
        oc8051_memory_interface1_add_2_root_add_937_2_carry_3_), .Y(
        oc8051_memory_interface1_n43) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u204 ( .A(
        oc8051_memory_interface1_idat_old_1_), .B(
        oc8051_memory_interface1_idat_old_9_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n117)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u203 ( .A(
        oc8051_memory_interface1_idat_cur_9_), .Y(
        oc8051_memory_interface1_n125) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u202 ( .A(
        oc8051_memory_interface1_n117), .B(oc8051_memory_interface1_n71), .C(
        oc8051_memory_interface1_n72), .D(oc8051_memory_interface1_n125), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_1_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u201 ( .A(
        oc8051_memory_interface1_idat_old_4_), .B(
        oc8051_memory_interface1_idat_old_12_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n120)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u200 ( .A(
        oc8051_memory_interface1_idat_cur_12_), .Y(
        oc8051_memory_interface1_n128) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u199 ( .A(
        oc8051_memory_interface1_n120), .B(oc8051_memory_interface1_n80), .C(
        oc8051_memory_interface1_n81), .D(oc8051_memory_interface1_n128), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_4_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u198 ( .A(
        oc8051_memory_interface1_idat_old_2_), .B(
        oc8051_memory_interface1_idat_old_10_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n118)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u197 ( .A(
        oc8051_memory_interface1_idat_cur_10_), .Y(
        oc8051_memory_interface1_n126) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u196 ( .A(
        oc8051_memory_interface1_n118), .B(oc8051_memory_interface1_n74), .C(
        oc8051_memory_interface1_n75), .D(oc8051_memory_interface1_n126), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_2_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u195 ( .A(
        oc8051_memory_interface1_idat_old_0_), .B(
        oc8051_memory_interface1_idat_old_8_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n116)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u194 ( .A(
        oc8051_memory_interface1_idat_cur_8_), .Y(
        oc8051_memory_interface1_n124) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u193 ( .A(
        oc8051_memory_interface1_n116), .B(oc8051_memory_interface1_n68), .C(
        oc8051_memory_interface1_n69), .D(oc8051_memory_interface1_n124), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_0_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u192 ( .A(
        oc8051_memory_interface1_idat_old_5_), .B(
        oc8051_memory_interface1_idat_old_13_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n121)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u191 ( .A(
        oc8051_memory_interface1_idat_cur_13_), .Y(
        oc8051_memory_interface1_n129) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u190 ( .A(
        oc8051_memory_interface1_n121), .B(oc8051_memory_interface1_n83), .C(
        oc8051_memory_interface1_n84), .D(oc8051_memory_interface1_n129), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_5_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u189 ( .A(
        oc8051_memory_interface1_idat_old_7_), .B(
        oc8051_memory_interface1_idat_old_15_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n123)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u188 ( .A(
        oc8051_memory_interface1_idat_cur_15_), .Y(
        oc8051_memory_interface1_n131) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u187 ( .A(
        oc8051_memory_interface1_n123), .B(oc8051_memory_interface1_n89), .C(
        oc8051_memory_interface1_n90), .D(oc8051_memory_interface1_n131), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_7_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u186 ( .A(
        oc8051_memory_interface1_idat_old_6_), .B(
        oc8051_memory_interface1_idat_old_14_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n122)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u185 ( .A(
        oc8051_memory_interface1_idat_cur_14_), .Y(
        oc8051_memory_interface1_n130) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u184 ( .A(
        oc8051_memory_interface1_n122), .B(oc8051_memory_interface1_n86), .C(
        oc8051_memory_interface1_n87), .D(oc8051_memory_interface1_n130), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_6_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u183 ( .A(
        oc8051_memory_interface1_idat_old_3_), .B(
        oc8051_memory_interface1_idat_old_11_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n119)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u182 ( .A(
        oc8051_memory_interface1_idat_cur_11_), .Y(
        oc8051_memory_interface1_n127) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u181 ( .A(
        oc8051_memory_interface1_n119), .B(oc8051_memory_interface1_n77), .C(
        oc8051_memory_interface1_n78), .D(oc8051_memory_interface1_n127), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_3_) );
  AND2_X1M_A12TS oc8051_memory_interface1_u180 ( .A(
        oc8051_memory_interface1_pc_buf_2_), .B(
        oc8051_memory_interface1_inc_pc), .Y(oc8051_memory_interface1_n42) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u179 ( .A(
        oc8051_memory_interface1_pc_buf_11_), .B(oc8051_memory_interface1_n64), 
        .Y(oc8051_memory_interface1_n41) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u178 ( .A(
        oc8051_memory_interface1_pc_buf_14_), .B(oc8051_memory_interface1_n56), 
        .Y(oc8051_memory_interface1_n40) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u177 ( .A(
        oc8051_memory_interface1_pc_buf_12_), .B(oc8051_memory_interface1_n54), 
        .Y(oc8051_memory_interface1_n39) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u176 ( .A(
        oc8051_memory_interface1_pc_buf_13_), .B(oc8051_memory_interface1_n55), 
        .Y(oc8051_memory_interface1_n38) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u175 ( .A(
        oc8051_memory_interface1_pc_buf_8_), .B(oc8051_memory_interface1_n61), 
        .Y(oc8051_memory_interface1_n37) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u174 ( .A(
        oc8051_memory_interface1_pc_buf_9_), .B(oc8051_memory_interface1_n62), 
        .Y(oc8051_memory_interface1_n36) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u173 ( .A(
        oc8051_memory_interface1_pc_buf_10_), .B(oc8051_memory_interface1_n63), 
        .Y(oc8051_memory_interface1_n35) );
  AND2_X1M_A12TS oc8051_memory_interface1_u172 ( .A(
        oc8051_memory_interface1_op_pos_0_), .B(
        oc8051_memory_interface1_pc_buf_0_), .Y(oc8051_memory_interface1_n34)
         );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u171 ( .A(
        oc8051_memory_interface1_pc_buf_5_), .B(oc8051_memory_interface1_n58), 
        .Y(oc8051_memory_interface1_n33) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u170 ( .A(
        oc8051_memory_interface1_pc_buf_6_), .B(oc8051_memory_interface1_n59), 
        .Y(oc8051_memory_interface1_n32) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u169 ( .A(
        oc8051_memory_interface1_pc_buf_4_), .B(oc8051_memory_interface1_n57), 
        .Y(oc8051_memory_interface1_n31) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u168 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .B(oc8051_memory_interface1_n42), 
        .Y(oc8051_memory_interface1_n30) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u167 ( .A(
        oc8051_memory_interface1_inc_pc), .B(
        oc8051_memory_interface1_pc_buf_2_), .Y(oc8051_memory_interface1_n29)
         );
  NAND2_X1M_A12TS oc8051_memory_interface1_u166 ( .A(
        oc8051_memory_interface1_n56), .B(oc8051_memory_interface1_pc_buf_14_), 
        .Y(oc8051_memory_interface1_n67) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u165 ( .A(
        oc8051_memory_interface1_pc_buf_15_), .B(oc8051_memory_interface1_n67), 
        .Y(oc8051_memory_interface1_pc_out_15_) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u164 ( .A(
        oc8051_memory_interface1_pc_buf_7_), .B(oc8051_memory_interface1_n60), 
        .Y(oc8051_memory_interface1_pc_out_7_) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u163 ( .A(
        oc8051_memory_interface1_n4240), .B(oc8051_memory_interface1_n65), .Y(
        oc8051_memory_interface1_n4560) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u162 ( .A(
        oc8051_memory_interface1_n4230), .B(oc8051_memory_interface1_n25), .Y(
        oc8051_memory_interface1_n4550) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u161 ( .A(
        oc8051_memory_interface1_n4200), .B(oc8051_memory_interface1_n22), .Y(
        oc8051_memory_interface1_n4520) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u160 ( .A(
        oc8051_memory_interface1_n4210), .B(oc8051_memory_interface1_n23), .Y(
        oc8051_memory_interface1_n4530) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u159 ( .A(
        oc8051_memory_interface1_n4220), .B(oc8051_memory_interface1_n24), .Y(
        oc8051_memory_interface1_n4540) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u158 ( .A(
        oc8051_memory_interface1_pc_buf_14_), .B(oc8051_memory_interface1_n46), 
        .Y(oc8051_memory_interface1_n66) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u157 ( .A(
        oc8051_memory_interface1_pc_buf_15_), .B(oc8051_memory_interface1_n66), 
        .Y(oc8051_memory_interface1_n4240) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u156 ( .A(
        oc8051_memory_interface1_pcs_source_0_), .B(pc[0]), .Y(
        oc8051_memory_interface1_pcs_result[0]) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u155 ( .A(
        oc8051_memory_interface1_n4250), .B(oc8051_memory_interface1_n4090), 
        .Y(oc8051_memory_interface1_n4410) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u154 ( .A(
        oc8051_memory_interface1_n4110), .B(
        oc8051_memory_interface1_add_0_root_add_937_2_carry_2_), .Y(
        oc8051_memory_interface1_n4430) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u153 ( .A(
        oc8051_memory_interface1_n4120), .B(oc8051_memory_interface1_n26), .Y(
        oc8051_memory_interface1_n4440) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u152 ( .A(
        oc8051_memory_interface1_n4130), .B(oc8051_memory_interface1_n15), .Y(
        oc8051_memory_interface1_n4450) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u151 ( .A(
        oc8051_memory_interface1_n4140), .B(oc8051_memory_interface1_n16), .Y(
        oc8051_memory_interface1_n4460) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u150 ( .A(
        oc8051_memory_interface1_n4150), .B(oc8051_memory_interface1_n17), .Y(
        oc8051_memory_interface1_n4470) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u149 ( .A(
        oc8051_memory_interface1_n4160), .B(oc8051_memory_interface1_n18), .Y(
        oc8051_memory_interface1_n4480) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u148 ( .A(
        oc8051_memory_interface1_pc_buf_11_), .B(oc8051_memory_interface1_n53), 
        .Y(oc8051_memory_interface1_n4200) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u147 ( .A(
        oc8051_memory_interface1_pc_buf_10_), .B(oc8051_memory_interface1_n52), 
        .Y(oc8051_memory_interface1_n4190) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u146 ( .A(
        oc8051_memory_interface1_pc_buf_9_), .B(oc8051_memory_interface1_n51), 
        .Y(oc8051_memory_interface1_n4180) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u145 ( .A(
        oc8051_memory_interface1_pc_buf_8_), .B(oc8051_memory_interface1_n50), 
        .Y(oc8051_memory_interface1_n4170) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u144 ( .A(
        oc8051_memory_interface1_pc_buf_7_), .B(oc8051_memory_interface1_n49), 
        .Y(oc8051_memory_interface1_n4160) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u143 ( .A(
        oc8051_memory_interface1_pc_buf_6_), .B(oc8051_memory_interface1_n48), 
        .Y(oc8051_memory_interface1_n4150) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u142 ( .A(
        oc8051_memory_interface1_pc_buf_5_), .B(oc8051_memory_interface1_n47), 
        .Y(oc8051_memory_interface1_n4140) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u141 ( .A(
        oc8051_memory_interface1_pc_buf_14_), .B(oc8051_memory_interface1_n46), 
        .Y(oc8051_memory_interface1_n4230) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u140 ( .A(
        oc8051_memory_interface1_pc_buf_13_), .B(oc8051_memory_interface1_n45), 
        .Y(oc8051_memory_interface1_n4220) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u139 ( .A(
        oc8051_memory_interface1_pc_buf_12_), .B(oc8051_memory_interface1_n44), 
        .Y(oc8051_memory_interface1_n4210) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u138 ( .A(
        oc8051_memory_interface1_pc_buf_4_), .B(oc8051_memory_interface1_n43), 
        .Y(oc8051_memory_interface1_n4130) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u137 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .B(
        oc8051_memory_interface1_add_2_root_add_937_2_carry_3_), .Y(
        oc8051_memory_interface1_n4120) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u136 ( .A(
        oc8051_memory_interface1_idat_cur_0_), .B(
        oc8051_memory_interface1_idat_cur_8_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n69)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u135 ( .A(
        oc8051_memory_interface1_idat_cur_1_), .B(
        oc8051_memory_interface1_idat_cur_9_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n72)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u134 ( .A(
        oc8051_memory_interface1_idat_cur_2_), .B(
        oc8051_memory_interface1_idat_cur_10_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n75)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u133 ( .A(
        oc8051_memory_interface1_idat_cur_3_), .B(
        oc8051_memory_interface1_idat_cur_11_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n78)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u132 ( .A(
        oc8051_memory_interface1_idat_cur_4_), .B(
        oc8051_memory_interface1_idat_cur_12_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n81)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u131 ( .A(
        oc8051_memory_interface1_idat_cur_5_), .B(
        oc8051_memory_interface1_idat_cur_13_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n84)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u130 ( .A(
        oc8051_memory_interface1_idat_cur_6_), .B(
        oc8051_memory_interface1_idat_cur_14_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n87)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u129 ( .A(
        oc8051_memory_interface1_idat_cur_7_), .B(
        oc8051_memory_interface1_idat_cur_15_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n90)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u128 ( .A(
        oc8051_memory_interface1_idat_old_16_), .B(
        oc8051_memory_interface1_idat_old_24_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n68)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u127 ( .A(
        oc8051_memory_interface1_idat_old_17_), .B(
        oc8051_memory_interface1_idat_old_25_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n71)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u126 ( .A(
        oc8051_memory_interface1_idat_old_18_), .B(
        oc8051_memory_interface1_idat_old_26_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n74)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u125 ( .A(
        oc8051_memory_interface1_idat_old_19_), .B(
        oc8051_memory_interface1_idat_old_27_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n77)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u124 ( .A(
        oc8051_memory_interface1_idat_old_20_), .B(
        oc8051_memory_interface1_idat_old_28_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n80)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u123 ( .A(
        oc8051_memory_interface1_idat_old_21_), .B(
        oc8051_memory_interface1_idat_old_29_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n83)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u122 ( .A(
        oc8051_memory_interface1_idat_old_22_), .B(
        oc8051_memory_interface1_idat_old_30_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n86)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u121 ( .A(
        oc8051_memory_interface1_idat_old_23_), .B(
        oc8051_memory_interface1_idat_old_31_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n89)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u120 ( .A(
        oc8051_memory_interface1_idat_old_26_), .B(
        oc8051_memory_interface1_idat_cur_2_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n98)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u119 ( .A(
        oc8051_memory_interface1_idat_old_24_), .B(
        oc8051_memory_interface1_idat_cur_0_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n92)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u118 ( .A(
        oc8051_memory_interface1_idat_old_25_), .B(
        oc8051_memory_interface1_idat_cur_1_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n95)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u117 ( .A(
        oc8051_memory_interface1_idat_old_27_), .B(
        oc8051_memory_interface1_idat_cur_3_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n101)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u116 ( .A(
        oc8051_memory_interface1_idat_old_28_), .B(
        oc8051_memory_interface1_idat_cur_4_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n104)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u115 ( .A(
        oc8051_memory_interface1_idat_old_29_), .B(
        oc8051_memory_interface1_idat_cur_5_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n107)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u114 ( .A(
        oc8051_memory_interface1_idat_old_30_), .B(
        oc8051_memory_interface1_idat_cur_6_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n110)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u113 ( .A(
        oc8051_memory_interface1_idat_old_31_), .B(
        oc8051_memory_interface1_idat_cur_7_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n113)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u112 ( .A(
        oc8051_memory_interface1_n113), .B(
        oc8051_memory_interface1_idat_cur_23_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n115)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u111 ( .A(
        oc8051_memory_interface1_idat_old_15_), .B(
        oc8051_memory_interface1_idat_cur_15_), .C(
        oc8051_memory_interface1_idat_old_23_), .D(
        oc8051_memory_interface1_idat_cur_23_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n114)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u110 ( .A(
        oc8051_memory_interface1_n114), .B(oc8051_memory_interface1_n115), 
        .S0(oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[7]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u109 ( .A(
        oc8051_memory_interface1_n95), .B(
        oc8051_memory_interface1_idat_cur_17_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n97)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u108 ( .A(
        oc8051_memory_interface1_idat_old_9_), .B(
        oc8051_memory_interface1_idat_cur_9_), .C(
        oc8051_memory_interface1_idat_old_17_), .D(
        oc8051_memory_interface1_idat_cur_17_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n96)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u107 ( .A(
        oc8051_memory_interface1_n96), .B(oc8051_memory_interface1_n97), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[1]) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u106 ( .A(
        oc8051_memory_interface1_op_pos_0_), .B(
        oc8051_memory_interface1_pc_buf_0_), .Y(oc8051_memory_interface1_n4090) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u105 ( .A(
        oc8051_memory_interface1_n98), .B(
        oc8051_memory_interface1_idat_cur_18_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n100)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u104 ( .A(
        oc8051_memory_interface1_idat_old_10_), .B(
        oc8051_memory_interface1_idat_cur_10_), .C(
        oc8051_memory_interface1_idat_old_18_), .D(
        oc8051_memory_interface1_idat_cur_18_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n99)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u103 ( .A(
        oc8051_memory_interface1_n99), .B(oc8051_memory_interface1_n100), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[2]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u102 ( .A(
        oc8051_memory_interface1_n92), .B(
        oc8051_memory_interface1_idat_cur_16_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n94)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u101 ( .A(
        oc8051_memory_interface1_idat_old_8_), .B(
        oc8051_memory_interface1_idat_cur_8_), .C(
        oc8051_memory_interface1_idat_old_16_), .D(
        oc8051_memory_interface1_idat_cur_16_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n93)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u100 ( .A(
        oc8051_memory_interface1_n93), .B(oc8051_memory_interface1_n94), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[0]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u99 ( .A(
        oc8051_memory_interface1_n101), .B(
        oc8051_memory_interface1_idat_cur_19_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n103)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u98 ( .A(
        oc8051_memory_interface1_idat_old_11_), .B(
        oc8051_memory_interface1_idat_cur_11_), .C(
        oc8051_memory_interface1_idat_old_19_), .D(
        oc8051_memory_interface1_idat_cur_19_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n102)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u97 ( .A(
        oc8051_memory_interface1_n102), .B(oc8051_memory_interface1_n103), 
        .S0(oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[3]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u96 ( .A(
        oc8051_memory_interface1_n104), .B(
        oc8051_memory_interface1_idat_cur_20_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n106)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u95 ( .A(
        oc8051_memory_interface1_idat_old_12_), .B(
        oc8051_memory_interface1_idat_cur_12_), .C(
        oc8051_memory_interface1_idat_old_20_), .D(
        oc8051_memory_interface1_idat_cur_20_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n105)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u94 ( .A(
        oc8051_memory_interface1_n105), .B(oc8051_memory_interface1_n106), 
        .S0(oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[4]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u93 ( .A(
        oc8051_memory_interface1_n107), .B(
        oc8051_memory_interface1_idat_cur_21_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n109)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u92 ( .A(
        oc8051_memory_interface1_idat_old_13_), .B(
        oc8051_memory_interface1_idat_cur_13_), .C(
        oc8051_memory_interface1_idat_old_21_), .D(
        oc8051_memory_interface1_idat_cur_21_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n108)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u91 ( .A(
        oc8051_memory_interface1_n108), .B(oc8051_memory_interface1_n109), 
        .S0(oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[5]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u90 ( .A(
        oc8051_memory_interface1_n110), .B(
        oc8051_memory_interface1_idat_cur_22_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n112)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u89 ( .A(
        oc8051_memory_interface1_idat_old_14_), .B(
        oc8051_memory_interface1_idat_cur_14_), .C(
        oc8051_memory_interface1_idat_old_22_), .D(
        oc8051_memory_interface1_idat_cur_22_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n111)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u88 ( .A(
        oc8051_memory_interface1_n111), .B(oc8051_memory_interface1_n112), 
        .S0(oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[6]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u87 ( .A(
        oc8051_memory_interface1_idat_cur_23_), .B(
        oc8051_memory_interface1_idat_cur_31_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n91)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u86 ( .A(
        oc8051_memory_interface1_idat_cur_31_), .Y(
        oc8051_memory_interface1_n139) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u85 ( .A(
        oc8051_memory_interface1_n89), .B(oc8051_memory_interface1_n90), .C(
        oc8051_memory_interface1_n91), .D(oc8051_memory_interface1_n139), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[7]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u84 ( .A(
        oc8051_memory_interface1_idat_cur_16_), .B(
        oc8051_memory_interface1_idat_cur_24_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n70)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u83 ( .A(
        oc8051_memory_interface1_idat_cur_24_), .Y(
        oc8051_memory_interface1_n132) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u82 ( .A(
        oc8051_memory_interface1_n68), .B(oc8051_memory_interface1_n69), .C(
        oc8051_memory_interface1_n70), .D(oc8051_memory_interface1_n132), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[0]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u81 ( .A(
        oc8051_memory_interface1_idat_cur_17_), .B(
        oc8051_memory_interface1_idat_cur_25_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n73)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u80 ( .A(
        oc8051_memory_interface1_idat_cur_25_), .Y(
        oc8051_memory_interface1_n133) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u79 ( .A(
        oc8051_memory_interface1_n71), .B(oc8051_memory_interface1_n72), .C(
        oc8051_memory_interface1_n73), .D(oc8051_memory_interface1_n133), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[1]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u78 ( .A(
        oc8051_memory_interface1_idat_cur_18_), .B(
        oc8051_memory_interface1_idat_cur_26_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n76)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u77 ( .A(
        oc8051_memory_interface1_idat_cur_26_), .Y(
        oc8051_memory_interface1_n134) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u76 ( .A(
        oc8051_memory_interface1_n74), .B(oc8051_memory_interface1_n75), .C(
        oc8051_memory_interface1_n76), .D(oc8051_memory_interface1_n134), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[2]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u75 ( .A(
        oc8051_memory_interface1_idat_cur_19_), .B(
        oc8051_memory_interface1_idat_cur_27_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n79)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u74 ( .A(
        oc8051_memory_interface1_idat_cur_27_), .Y(
        oc8051_memory_interface1_n135) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u73 ( .A(
        oc8051_memory_interface1_n77), .B(oc8051_memory_interface1_n78), .C(
        oc8051_memory_interface1_n79), .D(oc8051_memory_interface1_n135), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[3]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u72 ( .A(
        oc8051_memory_interface1_idat_cur_20_), .B(
        oc8051_memory_interface1_idat_cur_28_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n82)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u71 ( .A(
        oc8051_memory_interface1_idat_cur_28_), .Y(
        oc8051_memory_interface1_n136) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u70 ( .A(
        oc8051_memory_interface1_n80), .B(oc8051_memory_interface1_n81), .C(
        oc8051_memory_interface1_n82), .D(oc8051_memory_interface1_n136), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[4]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u69 ( .A(
        oc8051_memory_interface1_idat_cur_21_), .B(
        oc8051_memory_interface1_idat_cur_29_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n85)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u68 ( .A(
        oc8051_memory_interface1_idat_cur_29_), .Y(
        oc8051_memory_interface1_n137) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u67 ( .A(
        oc8051_memory_interface1_n83), .B(oc8051_memory_interface1_n84), .C(
        oc8051_memory_interface1_n85), .D(oc8051_memory_interface1_n137), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[5]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u66 ( .A(
        oc8051_memory_interface1_idat_cur_22_), .B(
        oc8051_memory_interface1_idat_cur_30_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n88)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u65 ( .A(
        oc8051_memory_interface1_idat_cur_30_), .Y(
        oc8051_memory_interface1_n138) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u64 ( .A(
        oc8051_memory_interface1_n86), .B(oc8051_memory_interface1_n87), .C(
        oc8051_memory_interface1_n88), .D(oc8051_memory_interface1_n138), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[6]) );
  OR2_X1M_A12TS oc8051_memory_interface1_u63 ( .A(oc8051_memory_interface1_n13), .B(pc[14]), .Y(oc8051_memory_interface1_n28) );
  AND2_X1M_A12TS oc8051_memory_interface1_u62 ( .A(
        oc8051_memory_interface1_u3_u7_z_14), .B(oc8051_memory_interface1_n8), 
        .Y(oc8051_memory_interface1_n27) );
  AND2_X1M_A12TS oc8051_memory_interface1_u61 ( .A(
        oc8051_memory_interface1_n4110), .B(
        oc8051_memory_interface1_add_0_root_add_937_2_carry_2_), .Y(
        oc8051_memory_interface1_n26) );
  OR2_X1M_A12TS oc8051_memory_interface1_u60 ( .A(oc8051_memory_interface1_n24), .B(oc8051_memory_interface1_n4220), .Y(oc8051_memory_interface1_n25) );
  OR2_X1M_A12TS oc8051_memory_interface1_u59 ( .A(oc8051_memory_interface1_n23), .B(oc8051_memory_interface1_n4210), .Y(oc8051_memory_interface1_n24) );
  OR2_X1M_A12TS oc8051_memory_interface1_u58 ( .A(oc8051_memory_interface1_n22), .B(oc8051_memory_interface1_n4200), .Y(oc8051_memory_interface1_n23) );
  OR2_X1M_A12TS oc8051_memory_interface1_u57 ( .A(oc8051_memory_interface1_n21), .B(oc8051_memory_interface1_n4190), .Y(oc8051_memory_interface1_n22) );
  OR2_X1M_A12TS oc8051_memory_interface1_u56 ( .A(oc8051_memory_interface1_n20), .B(oc8051_memory_interface1_n4180), .Y(oc8051_memory_interface1_n21) );
  OR2_X1M_A12TS oc8051_memory_interface1_u55 ( .A(oc8051_memory_interface1_n19), .B(oc8051_memory_interface1_n4170), .Y(oc8051_memory_interface1_n20) );
  OR2_X1M_A12TS oc8051_memory_interface1_u54 ( .A(oc8051_memory_interface1_n18), .B(oc8051_memory_interface1_n4160), .Y(oc8051_memory_interface1_n19) );
  OR2_X1M_A12TS oc8051_memory_interface1_u53 ( .A(oc8051_memory_interface1_n17), .B(oc8051_memory_interface1_n4150), .Y(oc8051_memory_interface1_n18) );
  OR2_X1M_A12TS oc8051_memory_interface1_u52 ( .A(oc8051_memory_interface1_n16), .B(oc8051_memory_interface1_n4140), .Y(oc8051_memory_interface1_n17) );
  OR2_X1M_A12TS oc8051_memory_interface1_u51 ( .A(oc8051_memory_interface1_n15), .B(oc8051_memory_interface1_n4130), .Y(oc8051_memory_interface1_n16) );
  OR2_X1M_A12TS oc8051_memory_interface1_u50 ( .A(oc8051_memory_interface1_n26), .B(oc8051_memory_interface1_n4120), .Y(oc8051_memory_interface1_n15) );
  OR2_X1M_A12TS oc8051_memory_interface1_u49 ( .A(pc[8]), .B(
        oc8051_memory_interface1_n3990), .Y(oc8051_memory_interface1_n14) );
  NOR2_X1A_A12TS oc8051_memory_interface1_u48 ( .A(
        oc8051_memory_interface1_n25), .B(oc8051_memory_interface1_n4230), .Y(
        oc8051_memory_interface1_n65) );
  OR2_X1M_A12TS oc8051_memory_interface1_u47 ( .A(oc8051_memory_interface1_n12), .B(pc[13]), .Y(oc8051_memory_interface1_n13) );
  OR2_X1M_A12TS oc8051_memory_interface1_u46 ( .A(oc8051_memory_interface1_n11), .B(pc[12]), .Y(oc8051_memory_interface1_n12) );
  OR2_X1M_A12TS oc8051_memory_interface1_u45 ( .A(oc8051_memory_interface1_n10), .B(pc[11]), .Y(oc8051_memory_interface1_n11) );
  OR2_X1M_A12TS oc8051_memory_interface1_u44 ( .A(oc8051_memory_interface1_n9), 
        .B(pc[10]), .Y(oc8051_memory_interface1_n10) );
  OR2_X1M_A12TS oc8051_memory_interface1_u43 ( .A(oc8051_memory_interface1_n14), .B(pc[9]), .Y(oc8051_memory_interface1_n9) );
  AND2_X1M_A12TS oc8051_memory_interface1_u42 ( .A(
        oc8051_memory_interface1_u3_u7_z_13), .B(oc8051_memory_interface1_n7), 
        .Y(oc8051_memory_interface1_n8) );
  AND2_X1M_A12TS oc8051_memory_interface1_u41 ( .A(
        oc8051_memory_interface1_u3_u7_z_12), .B(oc8051_memory_interface1_n6), 
        .Y(oc8051_memory_interface1_n7) );
  AND2_X1M_A12TS oc8051_memory_interface1_u40 ( .A(
        oc8051_memory_interface1_u3_u7_z_11), .B(oc8051_memory_interface1_n5), 
        .Y(oc8051_memory_interface1_n6) );
  AND2_X1M_A12TS oc8051_memory_interface1_u39 ( .A(
        oc8051_memory_interface1_u3_u7_z_10), .B(oc8051_memory_interface1_n4), 
        .Y(oc8051_memory_interface1_n5) );
  AND2_X1M_A12TS oc8051_memory_interface1_u38 ( .A(
        oc8051_memory_interface1_u3_u7_z_9), .B(oc8051_memory_interface1_n3), 
        .Y(oc8051_memory_interface1_n4) );
  AND2_X1M_A12TS oc8051_memory_interface1_u37 ( .A(
        oc8051_memory_interface1_u3_u7_z_8), .B(
        oc8051_memory_interface1_r390_carry_8_), .Y(
        oc8051_memory_interface1_n3) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u36 ( .A(
        oc8051_memory_interface1_u3_u7_z_14), .B(oc8051_memory_interface1_n8), 
        .Y(oc8051_memory_interface1_n4050) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u35 ( .A(
        oc8051_memory_interface1_u3_u7_z_9), .B(oc8051_memory_interface1_n3), 
        .Y(oc8051_memory_interface1_n4000) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u34 ( .A(
        oc8051_memory_interface1_u3_u7_z_10), .B(oc8051_memory_interface1_n4), 
        .Y(oc8051_memory_interface1_n4010) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u33 ( .A(
        oc8051_memory_interface1_u3_u7_z_11), .B(oc8051_memory_interface1_n5), 
        .Y(oc8051_memory_interface1_n4020) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u32 ( .A(
        oc8051_memory_interface1_u3_u7_z_12), .B(oc8051_memory_interface1_n6), 
        .Y(oc8051_memory_interface1_n4030) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u31 ( .A(
        oc8051_memory_interface1_u3_u7_z_13), .B(oc8051_memory_interface1_n7), 
        .Y(oc8051_memory_interface1_n4040) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u30 ( .A(pc[9]), .B(
        oc8051_memory_interface1_n14), .Y(oc8051_memory_interface1_n3840) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u29 ( .A(pc[14]), .B(
        oc8051_memory_interface1_n13), .Y(oc8051_memory_interface1_n3890) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u28 ( .A(pc[10]), .B(
        oc8051_memory_interface1_n9), .Y(oc8051_memory_interface1_n3850) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u27 ( .A(pc[11]), .B(
        oc8051_memory_interface1_n10), .Y(oc8051_memory_interface1_n3860) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u26 ( .A(pc[12]), .B(
        oc8051_memory_interface1_n11), .Y(oc8051_memory_interface1_n3870) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u25 ( .A(pc[13]), .B(
        oc8051_memory_interface1_n12), .Y(oc8051_memory_interface1_n3880) );
  AND2_X1M_A12TS oc8051_memory_interface1_u24 ( .A(
        oc8051_memory_interface1_n4250), .B(oc8051_memory_interface1_n4090), 
        .Y(oc8051_memory_interface1_n2) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u23 ( .A(pc[15]), .B(
        oc8051_memory_interface1_n28), .Y(oc8051_memory_interface1_n3900) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u22 ( .A(
        oc8051_memory_interface1_u3_u7_z_15), .B(oc8051_memory_interface1_n27), 
        .Y(oc8051_memory_interface1_n4060) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u21 ( .A(
        oc8051_memory_interface1_n4170), .B(oc8051_memory_interface1_n19), .Y(
        oc8051_memory_interface1_n4490) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u20 ( .A(
        oc8051_memory_interface1_n4180), .B(oc8051_memory_interface1_n20), .Y(
        oc8051_memory_interface1_n4500) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u19 ( .A(
        oc8051_memory_interface1_n4190), .B(oc8051_memory_interface1_n21), .Y(
        oc8051_memory_interface1_n4510) );
  XNOR2_X1M_A12TS oc8051_memory_interface1_u18 ( .A(
        oc8051_memory_interface1_n3990), .B(pc[8]), .Y(
        oc8051_memory_interface1_n3830) );
  XOR2_X1M_A12TS oc8051_memory_interface1_u17 ( .A(
        oc8051_memory_interface1_u3_u7_z_8), .B(
        oc8051_memory_interface1_r390_carry_8_), .Y(
        oc8051_memory_interface1_n3990) );
  NAND3_X2M_A12TS oc8051_memory_interface1_u16 ( .A(
        oc8051_memory_interface1_n191), .B(oc8051_memory_interface1_n192), .C(
        oc8051_memory_interface1_n193), .Y(rd_addr[1]) );
  AOI222_X1M_A12TS oc8051_memory_interface1_u15 ( .A0(
        oc8051_memory_interface1_imm_r[0]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_imm2_r[0]), .B1(
        oc8051_memory_interface1_n143), .C0(sp_w[0]), .C1(
        oc8051_memory_interface1_n142), .Y(oc8051_memory_interface1_n162) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u14 ( .A(
        oc8051_memory_interface1_n161), .B(oc8051_memory_interface1_n162), .Y(
        wr_addr[0]) );
  AOI22_X1M_A12TS oc8051_memory_interface1_u13 ( .A0(ri[0]), .A1(
        oc8051_memory_interface1_n174), .B0(op1_cur[0]), .B1(
        oc8051_memory_interface1_n184), .Y(oc8051_memory_interface1_n196) );
  OAI211_X2M_A12TS oc8051_memory_interface1_u12 ( .A0(
        oc8051_memory_interface1_n194), .A1(oc8051_memory_interface1_n171), 
        .B0(oc8051_memory_interface1_n195), .C0(oc8051_memory_interface1_n196), 
        .Y(rd_addr[0]) );
  AOI222_X1M_A12TS oc8051_memory_interface1_u11 ( .A0(
        oc8051_memory_interface1_imm_r[1]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_imm2_r[1]), .B1(
        oc8051_memory_interface1_n143), .C0(sp_w[1]), .C1(
        oc8051_memory_interface1_n142), .Y(oc8051_memory_interface1_n160) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u10 ( .A(
        oc8051_memory_interface1_n159), .B(oc8051_memory_interface1_n160), .Y(
        wr_addr[1]) );
  AOI22_X1M_A12TS oc8051_memory_interface1_u9 ( .A0(ri[2]), .A1(
        oc8051_memory_interface1_n174), .B0(op1_cur[2]), .B1(
        oc8051_memory_interface1_n184), .Y(oc8051_memory_interface1_n190) );
  OAI211_X1M_A12TS oc8051_memory_interface1_u8 ( .A0(
        oc8051_memory_interface1_n188), .A1(oc8051_memory_interface1_n171), 
        .B0(oc8051_memory_interface1_n189), .C0(oc8051_memory_interface1_n190), 
        .Y(rd_addr[2]) );
  OAI211_X1M_A12TS oc8051_memory_interface1_u7 ( .A0(
        oc8051_memory_interface1_n164), .A1(oc8051_memory_interface1_n165), 
        .B0(oc8051_memory_interface1_n166), .C0(oc8051_memory_interface1_n167), 
        .Y(rd_addr[7]) );
  AOI222_X1M_A12TS oc8051_memory_interface1_u6 ( .A0(
        oc8051_memory_interface1_imm_r[2]), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_imm2_r[2]), .B1(
        oc8051_memory_interface1_n143), .C0(sp_w[2]), .C1(
        oc8051_memory_interface1_n142), .Y(oc8051_memory_interface1_n158) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u5 ( .A(
        oc8051_memory_interface1_n157), .B(oc8051_memory_interface1_n158), .Y(
        wr_addr[2]) );
  NOR2_X2M_A12TS oc8051_memory_interface1_u4 ( .A(
        oc8051_memory_interface1_n266), .B(oc8051_memory_interface1_n243), .Y(
        oc8051_memory_interface1_n209) );
  AND2_X1M_A12TS oc8051_memory_interface1_u3 ( .A(
        oc8051_memory_interface1_pcs_source_0_), .B(pc[0]), .Y(
        oc8051_memory_interface1_n1) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_wr_r_reg ( .D(
        oc8051_memory_interface1_n5360), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_wr_r) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op_pos_reg_0_ ( .D(
        oc8051_memory_interface1_n477), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_op_pos_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op_pos_reg_2_ ( .D(
        oc8051_memory_interface1_n542), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_op_pos_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dstb_o_reg ( .D(
        oc8051_memory_interface1_n691), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_cyc_o) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dwe_o_reg ( .D(
        oc8051_memory_interface1_n1290), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_we_o) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op_pos_reg_1_ ( .D(
        oc8051_memory_interface1_n476), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_op_pos_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_istb_t_reg ( .D(
        oc8051_memory_interface1_n568), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_istb_t) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_13_ ( .D(
        oc8051_memory_interface1_n446), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_12_ ( .D(
        oc8051_memory_interface1_n447), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_11_ ( .D(
        oc8051_memory_interface1_n448), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_14_ ( .D(
        oc8051_memory_interface1_n445), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_10_ ( .D(
        oc8051_memory_interface1_n449), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_9_ ( .D(
        oc8051_memory_interface1_n450), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_8_ ( .D(
        oc8051_memory_interface1_n451), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_7_ ( .D(
        oc8051_memory_interface1_n452), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_6_ ( .D(
        oc8051_memory_interface1_n453), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_5_ ( .D(
        oc8051_memory_interface1_n454), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_4_ ( .D(
        oc8051_memory_interface1_n455), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_3_ ( .D(
        oc8051_memory_interface1_n456), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_3_) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_13_ ( .D(
        oc8051_memory_interface1_n462), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n377) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_12_ ( .D(
        oc8051_memory_interface1_n463), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n378) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_11_ ( .D(
        oc8051_memory_interface1_n464), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n379) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_10_ ( .D(
        oc8051_memory_interface1_n465), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n380) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_9_ ( .D(
        oc8051_memory_interface1_n466), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n381) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_8_ ( .D(
        oc8051_memory_interface1_n467), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n382) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_14_ ( .D(
        oc8051_memory_interface1_n461), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n383) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_15_ ( .D(
        oc8051_memory_interface1_n460), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n384) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_16_ ( .D(
        oc8051_memory_interface1_n509), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_16_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_17_ ( .D(
        oc8051_memory_interface1_n507), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_17_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_18_ ( .D(
        oc8051_memory_interface1_n505), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_18_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_19_ ( .D(
        oc8051_memory_interface1_n503), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_19_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_20_ ( .D(
        oc8051_memory_interface1_n501), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_20_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_21_ ( .D(
        oc8051_memory_interface1_n499), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_21_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_22_ ( .D(
        oc8051_memory_interface1_n497), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_22_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_23_ ( .D(
        oc8051_memory_interface1_n495), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_23_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_2_ ( .D(
        oc8051_memory_interface1_n457), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_wr_r2_reg ( .D(
        oc8051_memory_interface1_pc_wr_r), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_wr_r2) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_8_ ( .D(
        oc8051_memory_interface1_n525), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_9_ ( .D(
        oc8051_memory_interface1_n523), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_10_ ( .D(
        oc8051_memory_interface1_n521), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_11_ ( .D(
        oc8051_memory_interface1_n519), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_12_ ( .D(
        oc8051_memory_interface1_n517), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_13_ ( .D(
        oc8051_memory_interface1_n515), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_14_ ( .D(
        oc8051_memory_interface1_n513), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_15_ ( .D(
        oc8051_memory_interface1_n511), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dack_ir_reg ( .D(wbd_ack_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_dack_ir) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_0_ ( .D(
        oc8051_memory_interface1_n666), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_1_ ( .D(
        oc8051_memory_interface1_n667), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_2_ ( .D(
        oc8051_memory_interface1_n668), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_3_ ( .D(
        oc8051_memory_interface1_n669), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_4_ ( .D(
        oc8051_memory_interface1_n670), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_5_ ( .D(
        oc8051_memory_interface1_n671), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_6_ ( .D(
        oc8051_memory_interface1_n672), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_7_ ( .D(
        oc8051_memory_interface1_n673), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_24_ ( .D(
        oc8051_memory_interface1_n493), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_24_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_25_ ( .D(
        oc8051_memory_interface1_n491), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_25_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_26_ ( .D(
        oc8051_memory_interface1_n489), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_26_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_27_ ( .D(
        oc8051_memory_interface1_n487), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_27_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_28_ ( .D(
        oc8051_memory_interface1_n485), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_28_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_29_ ( .D(
        oc8051_memory_interface1_n483), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_29_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_30_ ( .D(
        oc8051_memory_interface1_n481), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_30_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_31_ ( .D(
        oc8051_memory_interface1_n479), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_31_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_15_ ( .D(
        oc8051_memory_interface1_n444), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_0_ ( .D(
        oc8051_memory_interface1_n475), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[0])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_24_ ( .D(
        oc8051_memory_interface1_n492), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_24_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_25_ ( .D(
        oc8051_memory_interface1_n490), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_25_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_26_ ( .D(
        oc8051_memory_interface1_n488), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_26_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_27_ ( .D(
        oc8051_memory_interface1_n486), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_27_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_28_ ( .D(
        oc8051_memory_interface1_n484), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_28_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_29_ ( .D(
        oc8051_memory_interface1_n482), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_29_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_30_ ( .D(
        oc8051_memory_interface1_n480), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_30_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_31_ ( .D(
        oc8051_memory_interface1_n478), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_31_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_0_ ( .D(
        oc8051_memory_interface1_n459), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_8_ ( .D(
        oc8051_memory_interface1_n524), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_9_ ( .D(
        oc8051_memory_interface1_n522), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_10_ ( .D(
        oc8051_memory_interface1_n520), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_11_ ( .D(
        oc8051_memory_interface1_n518), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_12_ ( .D(
        oc8051_memory_interface1_n516), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_13_ ( .D(
        oc8051_memory_interface1_n514), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_14_ ( .D(
        oc8051_memory_interface1_n512), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_15_ ( .D(
        oc8051_memory_interface1_n510), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_16_ ( .D(
        oc8051_memory_interface1_n508), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_16_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_17_ ( .D(
        oc8051_memory_interface1_n506), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_17_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_18_ ( .D(
        oc8051_memory_interface1_n504), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_18_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_19_ ( .D(
        oc8051_memory_interface1_n502), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_19_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_20_ ( .D(
        oc8051_memory_interface1_n500), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_20_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_21_ ( .D(
        oc8051_memory_interface1_n498), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_21_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_22_ ( .D(
        oc8051_memory_interface1_n496), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_22_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_23_ ( .D(
        oc8051_memory_interface1_n494), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_23_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_7_ ( .D(
        oc8051_memory_interface1_n468), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[7])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_6_ ( .D(
        oc8051_memory_interface1_n469), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[6])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_5_ ( .D(
        oc8051_memory_interface1_n470), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[5])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_4_ ( .D(
        oc8051_memory_interface1_n471), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[4])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_3_ ( .D(
        oc8051_memory_interface1_n472), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[3])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_2_ ( .D(
        oc8051_memory_interface1_n473), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[2])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_1_ ( .D(
        oc8051_memory_interface1_n474), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[1])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_0_ ( .D(
        oc8051_memory_interface1_n540), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_1_ ( .D(
        oc8051_memory_interface1_n538), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_2_ ( .D(
        oc8051_memory_interface1_n536), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_3_ ( .D(
        oc8051_memory_interface1_n534), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_4_ ( .D(
        oc8051_memory_interface1_n532), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_5_ ( .D(
        oc8051_memory_interface1_n530), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_6_ ( .D(
        oc8051_memory_interface1_n528), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_7_ ( .D(
        oc8051_memory_interface1_n526), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_1_ ( .D(
        oc8051_memory_interface1_n458), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_ack_t_reg ( .D(
        oc8051_memory_interface1_n543), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_ack_t) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imem_wait_reg ( .D(
        oc8051_memory_interface1_n569), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_imem_wait) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_0_ ( .D(
        oc8051_memory_interface1_n675), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_2_ ( .D(
        oc8051_memory_interface1_n677), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_3_ ( .D(
        oc8051_memory_interface1_n678), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_5_ ( .D(
        oc8051_memory_interface1_n680), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_6_ ( .D(
        oc8051_memory_interface1_n681), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_7_ ( .D(
        oc8051_memory_interface1_n682), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_7_ ( .D(
        oc8051_memory_interface1_n432), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_15_ ( .D(
        oc8051_memory_interface1_n440), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdone_reg ( .D(
        oc8051_memory_interface1_istb_t), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdone) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_0_ ( .D(
        oc8051_memory_interface1_n401), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_2_ ( .D(
        oc8051_memory_interface1_n403), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_3_ ( .D(
        oc8051_memory_interface1_n404), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_5_ ( .D(
        oc8051_memory_interface1_n406), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_6_ ( .D(
        oc8051_memory_interface1_n407), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_7_ ( .D(
        oc8051_memory_interface1_n408), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_1_ ( .D(
        oc8051_memory_interface1_n676), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_4_ ( .D(
        oc8051_memory_interface1_n679), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_0_ ( .D(
        oc8051_memory_interface1_n409), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_1_ ( .D(
        oc8051_memory_interface1_n410), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_2_ ( .D(
        oc8051_memory_interface1_n411), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_3_ ( .D(
        oc8051_memory_interface1_n412), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_4_ ( .D(
        oc8051_memory_interface1_n413), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_5_ ( .D(
        oc8051_memory_interface1_n414), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_6_ ( .D(
        oc8051_memory_interface1_n415), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_7_ ( .D(
        oc8051_memory_interface1_n416), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_1_ ( .D(
        oc8051_memory_interface1_n402), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_4_ ( .D(
        oc8051_memory_interface1_n405), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dmem_wait_reg ( .D(
        oc8051_memory_interface1_n691), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_dmem_wait) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_reti_reg ( .D(
        oc8051_memory_interface1_n1980), .CK(wb_clk_i), .R(wb_rst_i), .Q(reti)
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_ack_reg ( .D(
        oc8051_memory_interface1_n3700), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        int_ack) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_0_ ( .D(
        oc8051_memory_interface1_n425), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_1_ ( .D(
        oc8051_memory_interface1_n426), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_2_ ( .D(
        oc8051_memory_interface1_n427), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_3_ ( .D(
        oc8051_memory_interface1_n428), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_4_ ( .D(
        oc8051_memory_interface1_n429), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_5_ ( .D(
        oc8051_memory_interface1_n430), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_6_ ( .D(
        oc8051_memory_interface1_n431), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_8_ ( .D(
        oc8051_memory_interface1_n433), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_9_ ( .D(
        oc8051_memory_interface1_n434), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_10_ ( .D(
        oc8051_memory_interface1_n435), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_11_ ( .D(
        oc8051_memory_interface1_n436), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_12_ ( .D(
        oc8051_memory_interface1_n437), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_13_ ( .D(
        oc8051_memory_interface1_n438), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_14_ ( .D(
        oc8051_memory_interface1_n439), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_7_ ( .D(op3_n[7]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[7])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_0_ ( .D(op3_n[0]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[0])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_1_ ( .D(op3_n[1]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[1])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_2_ ( .D(op3_n[2]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[2])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_3_ ( .D(op3_n[3]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[3])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_4_ ( .D(op3_n[4]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[4])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_5_ ( .D(op3_n[5]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[5])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_6_ ( .D(op3_n[6]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[6])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rd_addr_r_reg ( .D(rd_addr[7]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rd_addr_r) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_4_ ( .D(op3_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_5_ ( .D(op3_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_6_ ( .D(op3_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_7_ ( .D(op3_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_5_ ( .D(op2_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_6_ ( .D(op2_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_7_ ( .D(op2_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_0_ ( .D(ri[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_1_ ( .D(ri[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_2_ ( .D(ri[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_3_ ( .D(ri[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_7_ ( .D(op2_n[7]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[7])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_0_ ( .D(op2_n[0]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[0])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_1_ ( .D(op2_n[1]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[1])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_2_ ( .D(op2_n[2]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[2])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_3_ ( .D(op2_n[3]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[3])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_4_ ( .D(op2_n[4]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[4])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_5_ ( .D(op2_n[5]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[5])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_6_ ( .D(op2_n[6]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[6])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_5_ ( .D(ri[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_6_ ( .D(ri[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_7_ ( .D(ri[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_0_ ( .D(op1_cur[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_1_ ( .D(op1_cur[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_2_ ( .D(op1_cur[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_3_ ( .D(bank_sel[0]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_4_ ( .D(ri[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_0_ ( .D(op2_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_1_ ( .D(op2_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_2_ ( .D(op2_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_3_ ( .D(op2_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_4_ ( .D(bank_sel[1]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_0_ ( .D(op3_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_1_ ( .D(op3_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_2_ ( .D(op3_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_3_ ( .D(op3_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_4_ ( .D(op2_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_ack_buff_reg ( .D(
        oc8051_memory_interface1_int_ack_t), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_ack_buff) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rd_ind_reg ( .D(
        oc8051_memory_interface1_n810), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_rd_ind) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_8_ ( .D(
        oc8051_memory_interface1_n552), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[8]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_9_ ( .D(
        oc8051_memory_interface1_n553), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[9]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_10_ ( .D(
        oc8051_memory_interface1_n554), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[10]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_11_ ( .D(
        oc8051_memory_interface1_n555), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[11]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_12_ ( .D(
        oc8051_memory_interface1_n556), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[12]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_13_ ( .D(
        oc8051_memory_interface1_n557), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[13]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_14_ ( .D(
        oc8051_memory_interface1_n558), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[14]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_15_ ( .D(
        oc8051_memory_interface1_n559), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[15]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_0_ ( .D(
        oc8051_memory_interface1_n560), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_1_ ( .D(
        oc8051_memory_interface1_n561), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_2_ ( .D(
        oc8051_memory_interface1_n562), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_3_ ( .D(
        oc8051_memory_interface1_n563), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_4_ ( .D(
        oc8051_memory_interface1_n564), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_5_ ( .D(
        oc8051_memory_interface1_n565), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_6_ ( .D(
        oc8051_memory_interface1_n566), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_7_ ( .D(
        oc8051_memory_interface1_n567), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_0_ ( .D(
        oc8051_memory_interface1_n544), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_1_ ( .D(
        oc8051_memory_interface1_n545), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_2_ ( .D(
        oc8051_memory_interface1_n546), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_3_ ( .D(
        oc8051_memory_interface1_n547), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_4_ ( .D(
        oc8051_memory_interface1_n548), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_5_ ( .D(
        oc8051_memory_interface1_n549), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_6_ ( .D(
        oc8051_memory_interface1_n550), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_7_ ( .D(
        oc8051_memory_interface1_n551), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[7]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_7 ( .A(pc[7]), .B(
        oc8051_memory_interface1_pcs_source_7_), .CI(
        oc8051_memory_interface1_r390_carry_7_), .CO(
        oc8051_memory_interface1_r390_carry_8_), .S(
        oc8051_memory_interface1_pcs_result[7]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_6 ( .A(pc[6]), .B(
        oc8051_memory_interface1_pcs_source_6_), .CI(
        oc8051_memory_interface1_r390_carry_6_), .CO(
        oc8051_memory_interface1_r390_carry_7_), .S(
        oc8051_memory_interface1_pcs_result[6]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_5 ( .A(pc[5]), .B(
        oc8051_memory_interface1_pcs_source_5_), .CI(
        oc8051_memory_interface1_r390_carry_5_), .CO(
        oc8051_memory_interface1_r390_carry_6_), .S(
        oc8051_memory_interface1_pcs_result[5]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_4 ( .A(pc[4]), .B(
        oc8051_memory_interface1_pcs_source_4_), .CI(
        oc8051_memory_interface1_r390_carry_4_), .CO(
        oc8051_memory_interface1_r390_carry_5_), .S(
        oc8051_memory_interface1_pcs_result[4]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_3 ( .A(pc[3]), .B(
        oc8051_memory_interface1_pcs_source_3_), .CI(
        oc8051_memory_interface1_r390_carry_3_), .CO(
        oc8051_memory_interface1_r390_carry_4_), .S(
        oc8051_memory_interface1_pcs_result[3]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_2 ( .A(pc[2]), .B(
        oc8051_memory_interface1_pcs_source_2_), .CI(
        oc8051_memory_interface1_r390_carry_2_), .CO(
        oc8051_memory_interface1_r390_carry_3_), .S(
        oc8051_memory_interface1_pcs_result[2]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_r390_u1_1 ( .A(pc[1]), .B(
        oc8051_memory_interface1_pcs_source_1_), .CI(
        oc8051_memory_interface1_n1), .CO(
        oc8051_memory_interface1_r390_carry_2_), .S(
        oc8051_memory_interface1_pcs_result[1]) );
  ADDF_X1M_A12TS oc8051_memory_interface1_add_2_root_add_937_2_u1_2 ( .A(
        oc8051_memory_interface1_pc_buf_2_), .B(
        oc8051_memory_interface1_op_pos_2_), .CI(
        oc8051_memory_interface1_add_2_root_add_937_2_carry_2_), .CO(
        oc8051_memory_interface1_add_2_root_add_937_2_carry_3_), .S(
        oc8051_memory_interface1_n4110) );
  ADDF_X1M_A12TS oc8051_memory_interface1_add_2_root_add_937_2_u1_1 ( .A(
        oc8051_memory_interface1_pc_buf_1_), .B(
        oc8051_memory_interface1_op_pos_1_), .CI(oc8051_memory_interface1_n34), 
        .CO(oc8051_memory_interface1_add_2_root_add_937_2_carry_2_), .S(
        oc8051_memory_interface1_n4100) );
  ADDF_X1M_A12TS oc8051_memory_interface1_add_0_root_add_937_2_u1_1 ( .A(
        oc8051_memory_interface1_n4100), .B(oc8051_memory_interface1_n4260), 
        .CI(oc8051_memory_interface1_n2), .CO(
        oc8051_memory_interface1_add_0_root_add_937_2_carry_2_), .S(
        oc8051_memory_interface1_n4420) );
  AO22_X4M_A12TS oc8051_memory_interface1_u517 ( .A0(bit_data), .A1(
        oc8051_memory_interface1_n322), .B0(sfr_bit), .B1(
        oc8051_memory_interface1_n674), .Y(bit_out) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u279 ( .A(rd_addr[3]), .B(rd_addr[6]), .Y(
        oc8051_sfr1_n219) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u278 ( .A(rd_addr[2]), .B(rd_addr[5]), .C(
        rd_addr[4]), .Y(oc8051_sfr1_n257) );
  AND4_X0P5M_A12TS oc8051_sfr1_u277 ( .A(rd_addr[1]), .B(oc8051_sfr1_n219), 
        .C(rd_addr[7]), .D(oc8051_sfr1_n257), .Y(oc8051_sfr1_n231) );
  INV_X0P5B_A12TS oc8051_sfr1_u276 ( .A(rd_addr[0]), .Y(oc8051_sfr1_n174) );
  AND4_X0P5M_A12TS oc8051_sfr1_u275 ( .A(wr_sfr[1]), .B(wr_sfr[0]), .C(
        oc8051_sfr1_n231), .D(oc8051_sfr1_n174), .Y(oc8051_sfr1_n35) );
  INV_X0P5B_A12TS oc8051_sfr1_u274 ( .A(rd_addr[1]), .Y(oc8051_sfr1_n185) );
  INV_X0P5B_A12TS oc8051_sfr1_u273 ( .A(rd_addr[2]), .Y(oc8051_sfr1_n172) );
  INV_X0P5B_A12TS oc8051_sfr1_u272 ( .A(rd_addr[3]), .Y(oc8051_sfr1_n183) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u271 ( .A(oc8051_sfr1_n174), .B(
        oc8051_sfr1_n185), .C(oc8051_sfr1_n172), .D(oc8051_sfr1_n183), .Y(
        oc8051_sfr1_n227) );
  INV_X0P5B_A12TS oc8051_sfr1_u270 ( .A(rd_addr[4]), .Y(oc8051_sfr1_n182) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u269 ( .A(oc8051_sfr1_n182), .B(rd_addr[5]), 
        .Y(oc8051_sfr1_n181) );
  INV_X0P5B_A12TS oc8051_sfr1_u268 ( .A(rd_addr[6]), .Y(oc8051_sfr1_n168) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u267 ( .AN(oc8051_sfr1_n181), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n42) );
  OAI211_X0P5M_A12TS oc8051_sfr1_u266 ( .A0(psw_set[1]), .A1(psw_set[0]), .B0(
        rd_addr[7]), .C0(oc8051_sfr1_n42), .Y(oc8051_sfr1_n228) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u265 ( .A(oc8051_sfr1_n174), .B(
        oc8051_sfr1_n172), .Y(oc8051_sfr1_n170) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u264 ( .A(wr_addr[3]), .B(oc8051_sfr1_n183), 
        .Y(oc8051_sfr1_n251) );
  INV_X0P5B_A12TS oc8051_sfr1_u263 ( .A(wr_addr[6]), .Y(oc8051_sfr1_n203) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u262 ( .A(oc8051_sfr1_n203), .B(rd_addr[6]), 
        .Y(oc8051_sfr1_n252) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u261 ( .A(wr_addr[4]), .B(rd_addr[4]), .Y(
        oc8051_sfr1_n255) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u260 ( .A(wr_addr[5]), .B(rd_addr[5]), .Y(
        oc8051_sfr1_n256) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u259 ( .A(oc8051_sfr1_n255), .B(
        oc8051_sfr1_n256), .Y(oc8051_sfr1_n253) );
  INV_X0P5B_A12TS oc8051_sfr1_u258 ( .A(wr_addr[7]), .Y(oc8051_sfr1_n250) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u257 ( .A(rd_addr[7]), .B(oc8051_sfr1_n250), 
        .Y(oc8051_sfr1_n254) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u256 ( .A(oc8051_sfr1_n251), .B(
        oc8051_sfr1_n252), .C(oc8051_sfr1_n253), .D(oc8051_sfr1_n254), .Y(
        oc8051_sfr1_n249) );
  AOI211_X0P5M_A12TS oc8051_sfr1_u255 ( .A0(oc8051_sfr1_n170), .A1(rd_addr[1]), 
        .B0(oc8051_sfr1_n249), .C0(oc8051_sfr1_n250), .Y(oc8051_sfr1_n236) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u254 ( .A(wr_addr[0]), .B(oc8051_sfr1_n174), 
        .Y(oc8051_sfr1_n246) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u253 ( .A(wr_addr[2]), .B(oc8051_sfr1_n172), 
        .Y(oc8051_sfr1_n247) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u252 ( .A(wr_addr[1]), .B(oc8051_sfr1_n185), 
        .Y(oc8051_sfr1_n248) );
  INV_X0P5B_A12TS oc8051_sfr1_u251 ( .A(oc8051_sfr1_n249), .Y(oc8051_sfr1_n210) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u250 ( .A(oc8051_sfr1_n246), .B(
        oc8051_sfr1_n247), .C(oc8051_sfr1_n248), .D(oc8051_sfr1_n210), .Y(
        oc8051_sfr1_n214) );
  INV_X0P5B_A12TS oc8051_sfr1_u249 ( .A(oc8051_sfr1_n214), .Y(oc8051_sfr1_n245) );
  INV_X0P5B_A12TS oc8051_sfr1_u248 ( .A(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_n200) );
  AND4_X0P5M_A12TS oc8051_sfr1_u247 ( .A(oc8051_sfr1_n245), .B(n_5_net_), .C(
        wr_addr[7]), .D(oc8051_sfr1_n200), .Y(oc8051_sfr1_n187) );
  AOI31_X0P5M_A12TS oc8051_sfr1_u246 ( .A0(oc8051_sfr1_wr_bit_r), .A1(n_5_net_), .A2(oc8051_sfr1_n236), .B0(oc8051_sfr1_n187), .Y(oc8051_sfr1_n229) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u245 ( .AN(wr_sfr[1]), .B(wr_sfr[0]), .Y(
        oc8051_sfr1_n198) );
  INV_X0P5B_A12TS oc8051_sfr1_u244 ( .A(rd_addr[5]), .Y(oc8051_sfr1_n186) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u243 ( .A(oc8051_sfr1_n186), .B(rd_addr[4]), 
        .C(oc8051_sfr1_n168), .Y(oc8051_sfr1_n40) );
  AND3_X0P5M_A12TS oc8051_sfr1_u242 ( .A(rd_addr[7]), .B(oc8051_sfr1_n183), 
        .C(oc8051_sfr1_n40), .Y(oc8051_sfr1_n235) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u241 ( .AN(wr_sfr[0]), .B(wr_sfr[1]), .Y(
        oc8051_sfr1_n197) );
  AND2_X0P5M_A12TS oc8051_sfr1_u240 ( .A(oc8051_sfr1_n197), .B(
        oc8051_sfr1_n235), .Y(oc8051_sfr1_n209) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_u239 ( .A0(oc8051_sfr1_n198), .A1(
        oc8051_sfr1_n235), .B0(oc8051_sfr1_n209), .C0(oc8051_sfr1_n174), .Y(
        oc8051_sfr1_n234) );
  INV_X0P5B_A12TS oc8051_sfr1_u238 ( .A(oc8051_sfr1_n234), .Y(oc8051_sfr1_n232) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u237 ( .A(rd_addr[2]), .B(rd_addr[1]), .Y(
        oc8051_sfr1_n233) );
  AOI32_X0P5M_A12TS oc8051_sfr1_u236 ( .A0(wr_sfr[0]), .A1(oc8051_sfr1_n231), 
        .A2(wr_sfr[1]), .B0(oc8051_sfr1_n232), .B1(oc8051_sfr1_n233), .Y(
        oc8051_sfr1_n230) );
  OA211_X0P5M_A12TS oc8051_sfr1_u235 ( .A0(oc8051_sfr1_n227), .A1(
        oc8051_sfr1_n228), .B0(oc8051_sfr1_n229), .C0(oc8051_sfr1_n230), .Y(
        oc8051_sfr1_n226) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u234 ( .A(wait_data), .B(oc8051_sfr1_n35), .C(
        oc8051_sfr1_n226), .Y(oc8051_sfr1_n1020) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u233 ( .A(rd_addr[3]), .B(rd_addr[5]), .Y(
        oc8051_sfr1_n175) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u232 ( .A(oc8051_sfr1_n1350), .B(
        oc8051_sfr1_n1340), .S0(rd_addr[4]), .Y(oc8051_sfr1_n223) );
  NAND3_X0P5A_A12TS oc8051_sfr1_u231 ( .A(rd_addr[3]), .B(rd_addr[6]), .C(
        oc8051_sfr1_n1380), .Y(oc8051_sfr1_n224) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u230 ( .A(oc8051_sfr1_n186), .B(
        oc8051_sfr1_n182), .Y(oc8051_sfr1_n184) );
  NAND3_X0P5A_A12TS oc8051_sfr1_u229 ( .A(oc8051_sfr1_n184), .B(
        oc8051_sfr1_n219), .C(oc8051_sfr1_n1320), .Y(oc8051_sfr1_n225) );
  OAI211_X0P5M_A12TS oc8051_sfr1_u228 ( .A0(oc8051_sfr1_n175), .A1(
        oc8051_sfr1_n223), .B0(oc8051_sfr1_n224), .C0(oc8051_sfr1_n225), .Y(
        oc8051_sfr1_n215) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u227 ( .A(oc8051_sfr1_n183), .B(rd_addr[6]), 
        .Y(oc8051_sfr1_n173) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u226 ( .A0(oc8051_sfr1_n1360), .A1(
        oc8051_sfr1_n173), .B0(oc8051_sfr1_n1290), .B1(oc8051_sfr1_n183), .Y(
        oc8051_sfr1_n221) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u225 ( .A(oc8051_sfr1_n1370), .B(rd_addr[3]), 
        .Y(oc8051_sfr1_n222) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u224 ( .A(oc8051_sfr1_n221), .B(
        oc8051_sfr1_n222), .S0(rd_addr[4]), .Y(oc8051_sfr1_n220) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u223 ( .AN(oc8051_sfr1_n184), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n55) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u222 ( .A0(oc8051_sfr1_n220), .A1(
        oc8051_sfr1_n186), .B0(oc8051_sfr1_n1330), .B1(oc8051_sfr1_n55), .Y(
        oc8051_sfr1_n216) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u221 ( .A0(oc8051_sfr1_n1280), .A1(
        oc8051_sfr1_n42), .B0(oc8051_sfr1_n1270), .B1(oc8051_sfr1_n40), .Y(
        oc8051_sfr1_n217) );
  AND2_X0P5M_A12TS oc8051_sfr1_u220 ( .A(oc8051_sfr1_n181), .B(
        oc8051_sfr1_n219), .Y(oc8051_sfr1_n53) );
  AND3_X0P5M_A12TS oc8051_sfr1_u219 ( .A(oc8051_sfr1_n219), .B(
        oc8051_sfr1_n182), .C(rd_addr[5]), .Y(oc8051_sfr1_n41) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u218 ( .A0(oc8051_sfr1_n1300), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_n1310), .B1(oc8051_sfr1_n41), .Y(
        oc8051_sfr1_n218) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u217 ( .AN(oc8051_sfr1_n215), .B(
        oc8051_sfr1_n216), .C(oc8051_sfr1_n217), .D(oc8051_sfr1_n218), .Y(
        oc8051_sfr1_n212) );
  INV_X0P5B_A12TS oc8051_sfr1_u216 ( .A(n_5_net_), .Y(oc8051_sfr1_n204) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u215 ( .A(oc8051_sfr1_n200), .B(
        oc8051_sfr1_n214), .C(oc8051_sfr1_n204), .Y(oc8051_sfr1_n213) );
  AOI31_X0P5M_A12TS oc8051_sfr1_u214 ( .A0(wr_addr[2]), .A1(wr_addr[1]), .A2(
        wr_addr[0]), .B0(oc8051_sfr1_wr_bit_r), .Y(oc8051_sfr1_n211) );
  AND3_X0P5M_A12TS oc8051_sfr1_u213 ( .A(n_5_net_), .B(oc8051_sfr1_n210), .C(
        oc8051_sfr1_n211), .Y(oc8051_sfr1_n191) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u212 ( .A(oc8051_sfr1_n209), .B(
        oc8051_sfr1_n191), .Y(oc8051_sfr1_n208) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u211 ( .A(oc8051_sfr1_prescaler_1_), .B(
        oc8051_sfr1_prescaler_0_), .Y(oc8051_sfr1_n1500) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u210 ( .A(oc8051_sfr1_prescaler_1_), .B(
        oc8051_sfr1_prescaler_0_), .Y(oc8051_sfr1_n31) );
  INV_X0P5B_A12TS oc8051_sfr1_u209 ( .A(oc8051_sfr1_n31), .Y(oc8051_sfr1_n205)
         );
  INV_X0P5B_A12TS oc8051_sfr1_u208 ( .A(oc8051_sfr1_prescaler_3_), .Y(
        oc8051_sfr1_n30) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u207 ( .A(oc8051_sfr1_n205), .B(
        oc8051_sfr1_n30), .Y(oc8051_sfr1_n206) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u206 ( .A(oc8051_sfr1_n206), .B(
        oc8051_sfr1_n205), .S0(oc8051_sfr1_prescaler_2_), .Y(oc8051_sfr1_n1510) );
  INV_X0P5B_A12TS oc8051_sfr1_u205 ( .A(oc8051_sfr1_prescaler_2_), .Y(
        oc8051_sfr1_n207) );
  OAI22_X0P5M_A12TS oc8051_sfr1_u204 ( .A0(oc8051_sfr1_n205), .A1(
        oc8051_sfr1_n30), .B0(oc8051_sfr1_n206), .B1(oc8051_sfr1_n207), .Y(
        oc8051_sfr1_n1520) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u203 ( .A(comp_sel[1]), .B(wr_addr[5]), .S0(
        wr_addr[4]), .Y(oc8051_sfr1_n202) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u202 ( .A(oc8051_sfr1_n202), .B(
        oc8051_sfr1_n203), .C(oc8051_sfr1_n204), .Y(oc8051_sfr1_n192) );
  OR3_X0P5M_A12TS oc8051_sfr1_u201 ( .A(wr_addr[1]), .B(wr_addr[2]), .C(
        wr_addr[0]), .Y(oc8051_sfr1_n199) );
  OAI21_X0P5M_A12TS oc8051_sfr1_u200 ( .A0(comp_sel[1]), .A1(wr_addr[5]), .B0(
        wr_addr[7]), .Y(oc8051_sfr1_n201) );
  AOI211_X0P5M_A12TS oc8051_sfr1_u199 ( .A0(oc8051_sfr1_n199), .A1(
        oc8051_sfr1_n200), .B0(oc8051_sfr1_n201), .C0(wr_addr[3]), .Y(
        oc8051_sfr1_n193) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u198 ( .A(oc8051_sfr1_n197), .B(
        oc8051_sfr1_n198), .Y(oc8051_sfr1_n195) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u197 ( .A(psw_set[1]), .B(psw_set[0]), .Y(
        oc8051_sfr1_n196) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u196 ( .A(oc8051_sfr1_n195), .B(
        oc8051_sfr1_n196), .S0(comp_sel[1]), .Y(oc8051_sfr1_n194) );
  AOI21_X0P5M_A12TS oc8051_sfr1_u195 ( .A0(oc8051_sfr1_n192), .A1(
        oc8051_sfr1_n193), .B0(oc8051_sfr1_n194), .Y(oc8051_sfr1_n189) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u194 ( .A(comp_sel[1]), .B(oc8051_sfr1_n191), 
        .Y(oc8051_sfr1_n190) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u193 ( .A(oc8051_sfr1_n189), .B(
        oc8051_sfr1_n190), .S0(comp_sel[0]), .Y(oc8051_sfr1_n188) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u192 ( .A(oc8051_sfr1_n187), .B(
        oc8051_sfr1_n188), .Y(comp_wait) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u191 ( .A(oc8051_sfr1_n35), .B(
        oc8051_sfr1_n1020), .Y(oc8051_sfr1_n33) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u190 ( .A(oc8051_sfr1_n172), .B(
        oc8051_sfr1_n186), .Y(oc8051_sfr1_n71) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u189 ( .A(rd_addr[0]), .B(rd_addr[6]), .C(
        oc8051_sfr1_n172), .Y(oc8051_sfr1_n72) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u188 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(
        oc8051_sfr1_n183), .Y(oc8051_sfr1_n169) );
  AND3_X0P5M_A12TS oc8051_sfr1_u187 ( .A(rd_addr[0]), .B(oc8051_sfr1_n182), 
        .C(oc8051_sfr1_n169), .Y(oc8051_sfr1_n73) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u186 ( .A0(oc8051_sfr1_ip_7_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[7]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[7]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n176) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u185 ( .A(oc8051_sfr1_n185), .B(rd_addr[0]), 
        .Y(oc8051_sfr1_n167) );
  AND2_X0P5M_A12TS oc8051_sfr1_u184 ( .A(oc8051_sfr1_n173), .B(
        oc8051_sfr1_n167), .Y(oc8051_sfr1_n68) );
  AND4_X0P5M_A12TS oc8051_sfr1_u183 ( .A(oc8051_sfr1_n174), .B(
        oc8051_sfr1_n185), .C(oc8051_sfr1_n182), .D(oc8051_sfr1_n186), .Y(
        oc8051_sfr1_n171) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u182 ( .AN(oc8051_sfr1_n171), .B(rd_addr[3]), 
        .Y(oc8051_sfr1_n69) );
  AND2_X0P5M_A12TS oc8051_sfr1_u181 ( .A(oc8051_sfr1_n173), .B(
        oc8051_sfr1_n170), .Y(oc8051_sfr1_n70) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u180 ( .A0(oc8051_sfr1_tl0[7]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_7_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[7]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n177) );
  AND3_X0P5M_A12TS oc8051_sfr1_u179 ( .A(oc8051_sfr1_n172), .B(
        oc8051_sfr1_n168), .C(oc8051_sfr1_n184), .Y(oc8051_sfr1_n65) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u178 ( .A(rd_addr[1]), .B(rd_addr[3]), .C(
        oc8051_sfr1_n174), .Y(oc8051_sfr1_n66) );
  AND4_X0P5M_A12TS oc8051_sfr1_u177 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(
        oc8051_sfr1_n172), .D(oc8051_sfr1_n183), .Y(oc8051_sfr1_n67) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u176 ( .A0(oc8051_sfr1_p3_data_7_), .A1(
        oc8051_sfr1_n65), .B0(sp[7]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[7]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n178) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u175 ( .AN(oc8051_sfr1_n167), .B(rd_addr[3]), 
        .Y(oc8051_sfr1_n60) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u174 ( .A(oc8051_sfr1_n182), .B(rd_addr[0]), 
        .C(oc8051_sfr1_n183), .Y(oc8051_sfr1_n61) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u173 ( .AN(oc8051_sfr1_n181), .B(
        oc8051_sfr1_n174), .Y(oc8051_sfr1_n63) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u172 ( .A(rd_addr[3]), .B(rd_addr[5]), .C(
        oc8051_sfr1_n172), .Y(oc8051_sfr1_n64) );
  AO22_X0P5M_A12TS oc8051_sfr1_u171 ( .A0(oc8051_sfr1_sbuf[7]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[7]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n180) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u170 ( .A0(dptr_lo[7]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_7_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n180), 
        .Y(oc8051_sfr1_n179) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u169 ( .A(oc8051_sfr1_n176), .B(
        oc8051_sfr1_n177), .C(oc8051_sfr1_n178), .D(oc8051_sfr1_n179), .Y(
        oc8051_sfr1_n160) );
  INV_X0P5B_A12TS oc8051_sfr1_u168 ( .A(oc8051_sfr1_n175), .Y(oc8051_sfr1_n54)
         );
  AOI222_X0P5M_A12TS oc8051_sfr1_u167 ( .A0(oc8051_sfr1_p1_data_7_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_7_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_7_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n161) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u166 ( .A(oc8051_sfr1_n168), .B(rd_addr[2]), 
        .C(oc8051_sfr1_n174), .Y(oc8051_sfr1_n51) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u165 ( .A(oc8051_sfr1_n168), .B(rd_addr[0]), 
        .C(oc8051_sfr1_n172), .Y(oc8051_sfr1_n52) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u164 ( .A0(oc8051_sfr1_rcap2h[7]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[7]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n164) );
  AND3_X0P5M_A12TS oc8051_sfr1_u163 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(
        oc8051_sfr1_n173), .Y(oc8051_sfr1_n49) );
  AND3_X0P5M_A12TS oc8051_sfr1_u162 ( .A(oc8051_sfr1_n171), .B(
        oc8051_sfr1_n172), .C(oc8051_sfr1_n173), .Y(oc8051_sfr1_n50) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u161 ( .A0(oc8051_sfr1_tl1[7]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_7_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n165) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u160 ( .AN(oc8051_sfr1_n170), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n46) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u159 ( .AN(oc8051_sfr1_n169), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n47) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u158 ( .AN(oc8051_sfr1_n167), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n48) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u157 ( .A0(oc8051_sfr1_th2[7]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_7_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[7]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n166)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u156 ( .A(oc8051_sfr1_n164), .B(
        oc8051_sfr1_n165), .C(oc8051_sfr1_n166), .Y(oc8051_sfr1_n162) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u155 ( .A0(acc[7]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_7_), .B1(oc8051_sfr1_n41), .C0(cy), .C1(
        oc8051_sfr1_n42), .Y(oc8051_sfr1_n163) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u154 ( .AN(oc8051_sfr1_n160), .B(
        oc8051_sfr1_n161), .C(oc8051_sfr1_n162), .D(oc8051_sfr1_n163), .Y(
        oc8051_sfr1_n159) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u153 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n159), .B0(des_acc[7]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n158) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u152 ( .B0(sfr_out[7]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n158), .Y(oc8051_sfr1_n237) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u151 ( .A0(oc8051_sfr1_ip_6_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[6]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[6]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n153) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u150 ( .A0(oc8051_sfr1_tl0[6]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_6_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[6]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n154) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u149 ( .A0(oc8051_sfr1_p3_data_6_), .A1(
        oc8051_sfr1_n65), .B0(sp[6]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[6]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n155) );
  AO22_X0P5M_A12TS oc8051_sfr1_u148 ( .A0(oc8051_sfr1_sbuf[6]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[6]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n157) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u147 ( .A0(dptr_lo[6]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_6_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n157), 
        .Y(oc8051_sfr1_n156) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u146 ( .A(oc8051_sfr1_n153), .B(
        oc8051_sfr1_n154), .C(oc8051_sfr1_n155), .D(oc8051_sfr1_n156), .Y(
        oc8051_sfr1_n146) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u145 ( .A0(oc8051_sfr1_p1_data_6_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_6_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_6_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n147) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u144 ( .A0(oc8051_sfr1_rcap2h[6]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[6]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n150) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u143 ( .A0(oc8051_sfr1_tl1[6]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tr1), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n151) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u142 ( .A0(oc8051_sfr1_th2[6]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_6_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[6]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n152)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u141 ( .A(oc8051_sfr1_n150), .B(
        oc8051_sfr1_n151), .C(oc8051_sfr1_n152), .Y(oc8051_sfr1_n148) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u140 ( .A0(acc[6]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_6_), .B1(oc8051_sfr1_n41), .C0(srcac), .C1(
        oc8051_sfr1_n42), .Y(oc8051_sfr1_n149) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u139 ( .AN(oc8051_sfr1_n146), .B(
        oc8051_sfr1_n147), .C(oc8051_sfr1_n148), .D(oc8051_sfr1_n149), .Y(
        oc8051_sfr1_n145) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u138 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n145), .B0(des_acc[6]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n144) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u137 ( .B0(sfr_out[6]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n144), .Y(oc8051_sfr1_n238) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u136 ( .A0(oc8051_sfr1_ip_5_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[5]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[5]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n139) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u135 ( .A0(oc8051_sfr1_tl0[5]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_5_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[5]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n140) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u134 ( .A0(oc8051_sfr1_p3_data_5_), .A1(
        oc8051_sfr1_n65), .B0(sp[5]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[5]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n141) );
  AO22_X0P5M_A12TS oc8051_sfr1_u133 ( .A0(oc8051_sfr1_sbuf[5]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[5]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n143) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u132 ( .A0(dptr_lo[5]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_5_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n143), 
        .Y(oc8051_sfr1_n142) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u131 ( .A(oc8051_sfr1_n139), .B(
        oc8051_sfr1_n140), .C(oc8051_sfr1_n141), .D(oc8051_sfr1_n142), .Y(
        oc8051_sfr1_n132) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u130 ( .A0(oc8051_sfr1_p1_data_5_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_5_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_5_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n133) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u129 ( .A0(oc8051_sfr1_rcap2h[5]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[5]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n136) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u128 ( .A0(oc8051_sfr1_tl1[5]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_5_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n137) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u127 ( .A0(oc8051_sfr1_th2[5]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_rclk), .B1(oc8051_sfr1_n47), .C0(
        oc8051_sfr1_rcap2l[5]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n138) );
  AND3_X0P5M_A12TS oc8051_sfr1_u126 ( .A(oc8051_sfr1_n136), .B(
        oc8051_sfr1_n137), .C(oc8051_sfr1_n138), .Y(oc8051_sfr1_n134) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u125 ( .A0(acc[5]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_5_), .B1(oc8051_sfr1_n41), .C0(
        oc8051_sfr1_psw_5_), .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n135) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u124 ( .AN(oc8051_sfr1_n132), .B(
        oc8051_sfr1_n133), .C(oc8051_sfr1_n134), .D(oc8051_sfr1_n135), .Y(
        oc8051_sfr1_n131) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u123 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n131), .B0(des_acc[5]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n130) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u122 ( .B0(sfr_out[5]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n130), .Y(oc8051_sfr1_n239) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u121 ( .A0(oc8051_sfr1_ip_4_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[4]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[4]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n125) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u120 ( .A0(oc8051_sfr1_tl0[4]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_4_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[4]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n126) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u119 ( .A0(oc8051_sfr1_p3_data_4_), .A1(
        oc8051_sfr1_n65), .B0(sp[4]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[4]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n127) );
  AO22_X0P5M_A12TS oc8051_sfr1_u118 ( .A0(oc8051_sfr1_sbuf[4]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[4]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n129) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u117 ( .A0(dptr_lo[4]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_4_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n129), 
        .Y(oc8051_sfr1_n128) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u116 ( .A(oc8051_sfr1_n125), .B(
        oc8051_sfr1_n126), .C(oc8051_sfr1_n127), .D(oc8051_sfr1_n128), .Y(
        oc8051_sfr1_n118) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u115 ( .A0(oc8051_sfr1_p1_data_4_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_4_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_4_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n119) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u114 ( .A0(oc8051_sfr1_rcap2h[4]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[4]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n122) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u113 ( .A0(oc8051_sfr1_tl1[4]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tr0), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n123) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u112 ( .A0(oc8051_sfr1_th2[4]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_tclk), .B1(oc8051_sfr1_n47), .C0(
        oc8051_sfr1_rcap2l[4]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n124) );
  AND3_X0P5M_A12TS oc8051_sfr1_u111 ( .A(oc8051_sfr1_n122), .B(
        oc8051_sfr1_n123), .C(oc8051_sfr1_n124), .Y(oc8051_sfr1_n120) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u110 ( .A0(acc[4]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_4_), .B1(oc8051_sfr1_n41), .C0(
        oc8051_sfr1_psw_4_), .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n121) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u109 ( .AN(oc8051_sfr1_n118), .B(
        oc8051_sfr1_n119), .C(oc8051_sfr1_n120), .D(oc8051_sfr1_n121), .Y(
        oc8051_sfr1_n117) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u108 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n117), .B0(des_acc[4]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n116) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u107 ( .B0(sfr_out[4]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n116), .Y(oc8051_sfr1_n240) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u106 ( .A0(oc8051_sfr1_ip_3_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[3]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[3]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n111) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u105 ( .A0(oc8051_sfr1_tl0[3]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_3_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[3]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n112) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u104 ( .A0(oc8051_sfr1_p3_data_3_), .A1(
        oc8051_sfr1_n65), .B0(sp[3]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[3]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n113) );
  AO22_X0P5M_A12TS oc8051_sfr1_u103 ( .A0(oc8051_sfr1_sbuf[3]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[3]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n115) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u102 ( .A0(dptr_lo[3]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_3_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n115), 
        .Y(oc8051_sfr1_n114) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u101 ( .A(oc8051_sfr1_n111), .B(
        oc8051_sfr1_n112), .C(oc8051_sfr1_n113), .D(oc8051_sfr1_n114), .Y(
        oc8051_sfr1_n104) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u100 ( .A0(oc8051_sfr1_p1_data_3_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_3_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_3_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n105) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u99 ( .A0(oc8051_sfr1_rcap2h[3]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[3]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n108) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u98 ( .A0(oc8051_sfr1_tl1[3]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_3_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n109) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u97 ( .A0(oc8051_sfr1_th2[3]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_3_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[3]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n110)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u96 ( .A(oc8051_sfr1_n108), .B(oc8051_sfr1_n109), .C(oc8051_sfr1_n110), .Y(oc8051_sfr1_n106) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u95 ( .A0(acc[3]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_3_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_3_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n107) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u94 ( .AN(oc8051_sfr1_n104), .B(
        oc8051_sfr1_n105), .C(oc8051_sfr1_n106), .D(oc8051_sfr1_n107), .Y(
        oc8051_sfr1_n103) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u93 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n103), .B0(des_acc[3]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n102) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u92 ( .B0(sfr_out[3]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n102), .Y(oc8051_sfr1_n241) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u91 ( .A0(oc8051_sfr1_ip_2_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[2]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[2]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n97) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u90 ( .A0(oc8051_sfr1_tl0[2]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_2_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[2]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n98) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u89 ( .A0(oc8051_sfr1_p3_data_2_), .A1(
        oc8051_sfr1_n65), .B0(sp[2]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[2]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n99) );
  AO22_X0P5M_A12TS oc8051_sfr1_u88 ( .A0(oc8051_sfr1_sbuf[2]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[2]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n101) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u87 ( .A0(dptr_lo[2]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_2_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n101), 
        .Y(oc8051_sfr1_n100) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u86 ( .A(oc8051_sfr1_n97), .B(oc8051_sfr1_n98), 
        .C(oc8051_sfr1_n99), .D(oc8051_sfr1_n100), .Y(oc8051_sfr1_n90) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u85 ( .A0(oc8051_sfr1_p1_data_2_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_2_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_2_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n91) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u84 ( .A0(oc8051_sfr1_rcap2h[2]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[2]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n94) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u83 ( .A0(oc8051_sfr1_tl1[2]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_2_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n95) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u82 ( .A0(oc8051_sfr1_th2[2]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_2_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[2]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n96)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u81 ( .A(oc8051_sfr1_n94), .B(oc8051_sfr1_n95), 
        .C(oc8051_sfr1_n96), .Y(oc8051_sfr1_n92) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u80 ( .A0(acc[2]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_2_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_2_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n93) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u79 ( .AN(oc8051_sfr1_n90), .B(
        oc8051_sfr1_n91), .C(oc8051_sfr1_n92), .D(oc8051_sfr1_n93), .Y(
        oc8051_sfr1_n89) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u78 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n89), .B0(des_acc[2]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n88) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u77 ( .B0(sfr_out[2]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n88), .Y(oc8051_sfr1_n242) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u76 ( .A0(oc8051_sfr1_ip_1_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[1]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[1]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n83) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u75 ( .A0(oc8051_sfr1_tl0[1]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_1_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[1]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n84) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u74 ( .A0(oc8051_sfr1_p3_data_1_), .A1(
        oc8051_sfr1_n65), .B0(sp[1]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[1]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n85) );
  AO22_X0P5M_A12TS oc8051_sfr1_u73 ( .A0(oc8051_sfr1_sbuf[1]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[1]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n87) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u72 ( .A0(dptr_lo[1]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_1_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n87), 
        .Y(oc8051_sfr1_n86) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u71 ( .A(oc8051_sfr1_n83), .B(oc8051_sfr1_n84), 
        .C(oc8051_sfr1_n85), .D(oc8051_sfr1_n86), .Y(oc8051_sfr1_n76) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u70 ( .A0(oc8051_sfr1_p1_data_1_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_1_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_1_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n77) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u69 ( .A0(oc8051_sfr1_rcap2h[1]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[1]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n80) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u68 ( .A0(oc8051_sfr1_tl1[1]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_1_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n81) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u67 ( .A0(oc8051_sfr1_th2[1]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_1_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[1]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n82)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u66 ( .A(oc8051_sfr1_n80), .B(oc8051_sfr1_n81), 
        .C(oc8051_sfr1_n82), .Y(oc8051_sfr1_n78) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u65 ( .A0(acc[1]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_1_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_1_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n79) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u64 ( .AN(oc8051_sfr1_n76), .B(
        oc8051_sfr1_n77), .C(oc8051_sfr1_n78), .D(oc8051_sfr1_n79), .Y(
        oc8051_sfr1_n75) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u63 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n75), .B0(des_acc[1]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n74) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u62 ( .B0(sfr_out[1]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n74), .Y(oc8051_sfr1_n243) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u61 ( .A0(oc8051_sfr1_ip_0_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[0]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[0]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n56) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u60 ( .A0(oc8051_sfr1_tl0[0]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_0_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[0]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n57) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u59 ( .A0(oc8051_sfr1_p3_data_0_), .A1(
        oc8051_sfr1_n65), .B0(sp[0]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[0]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n58) );
  AO22_X0P5M_A12TS oc8051_sfr1_u58 ( .A0(oc8051_sfr1_sbuf[0]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[0]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n62) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u57 ( .A0(dptr_lo[0]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_0_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n62), 
        .Y(oc8051_sfr1_n59) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u56 ( .A(oc8051_sfr1_n56), .B(oc8051_sfr1_n57), 
        .C(oc8051_sfr1_n58), .D(oc8051_sfr1_n59), .Y(oc8051_sfr1_n36) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u55 ( .A0(oc8051_sfr1_p1_data_0_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_0_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_0_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n37) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u54 ( .A0(oc8051_sfr1_rcap2h[0]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[0]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n43) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u53 ( .A0(oc8051_sfr1_tl1[0]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_0_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n44) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u52 ( .A0(oc8051_sfr1_th2[0]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_0_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[0]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n45)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u51 ( .A(oc8051_sfr1_n43), .B(oc8051_sfr1_n44), 
        .C(oc8051_sfr1_n45), .Y(oc8051_sfr1_n38) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u50 ( .A0(acc[0]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_0_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_0_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n39) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u49 ( .AN(oc8051_sfr1_n36), .B(
        oc8051_sfr1_n37), .C(oc8051_sfr1_n38), .D(oc8051_sfr1_n39), .Y(
        oc8051_sfr1_n34) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u48 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n34), .B0(des_acc[0]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n32) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u47 ( .B0(sfr_out[0]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n32), .Y(oc8051_sfr1_n244) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u46 ( .A(oc8051_sfr1_n30), .B(
        oc8051_sfr1_prescaler_2_), .C(oc8051_sfr1_n31), .Y(oc8051_sfr1_n259)
         );
  INV_X0P5B_A12TS oc8051_sfr1_u45 ( .A(oc8051_sfr1_prescaler_0_), .Y(
        oc8051_sfr1_n258) );
  MXT4_X1M_A12TS oc8051_sfr1_u44 ( .A(oc8051_sfr1_tclk), .B(
        oc8051_sfr1_t2con_6_), .C(oc8051_sfr1_rclk), .D(oc8051_sfr1_t2con_7_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n17) );
  MXT4_X1M_A12TS oc8051_sfr1_u43 ( .A(oc8051_sfr1_t2con_0_), .B(
        oc8051_sfr1_t2con_2_), .C(oc8051_sfr1_t2con_1_), .D(
        oc8051_sfr1_t2con_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n16) );
  MXT2_X1M_A12TS oc8051_sfr1_u42 ( .A(oc8051_sfr1_n16), .B(oc8051_sfr1_n17), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1380) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u41 ( .A(oc8051_sfr1_ip_0_), .B(
        oc8051_sfr1_ip_2_), .C(oc8051_sfr1_ip_1_), .D(oc8051_sfr1_ip_3_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n22) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u40 ( .A(oc8051_sfr1_scon_0_), .B(
        oc8051_sfr1_scon_2_), .C(oc8051_sfr1_scon_1_), .D(oc8051_sfr1_scon_3_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n18) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u39 ( .A(oc8051_sfr1_ie_4_), .B(
        oc8051_sfr1_ie_6_), .C(oc8051_sfr1_ie_5_), .D(oc8051_sfr1_ie_7_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n21) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u38 ( .A(oc8051_sfr1_ip_4_), .B(
        oc8051_sfr1_ip_6_), .C(oc8051_sfr1_ip_5_), .D(oc8051_sfr1_ip_7_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n23) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u37 ( .A(oc8051_sfr1_scon_4_), .B(
        oc8051_sfr1_scon_6_), .C(oc8051_sfr1_scon_5_), .D(oc8051_sfr1_scon_7_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n19) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u36 ( .A(oc8051_sfr1_ie_0_), .B(
        oc8051_sfr1_ie_2_), .C(oc8051_sfr1_ie_1_), .D(oc8051_sfr1_ie_3_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n20) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u35 ( .A(oc8051_sfr1_n22), .B(oc8051_sfr1_n23), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1340) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u34 ( .A(oc8051_sfr1_n20), .B(oc8051_sfr1_n21), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1350) );
  MXT4_X1M_A12TS oc8051_sfr1_u33 ( .A(oc8051_sfr1_b_reg_4_), .B(
        oc8051_sfr1_b_reg_6_), .C(oc8051_sfr1_b_reg_5_), .D(
        oc8051_sfr1_b_reg_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n15) );
  MXT4_X1M_A12TS oc8051_sfr1_u32 ( .A(oc8051_sfr1_b_reg_0_), .B(
        oc8051_sfr1_b_reg_2_), .C(oc8051_sfr1_b_reg_1_), .D(
        oc8051_sfr1_b_reg_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n14) );
  MXT2_X1M_A12TS oc8051_sfr1_u31 ( .A(oc8051_sfr1_n14), .B(oc8051_sfr1_n15), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1330) );
  MXT4_X1M_A12TS oc8051_sfr1_u30 ( .A(acc[4]), .B(acc[6]), .C(acc[5]), .D(
        acc[7]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n13) );
  MXT4_X1M_A12TS oc8051_sfr1_u29 ( .A(acc[0]), .B(acc[2]), .C(acc[1]), .D(
        acc[3]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n12) );
  MXT2_X1M_A12TS oc8051_sfr1_u28 ( .A(oc8051_sfr1_n12), .B(oc8051_sfr1_n13), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1270) );
  MXT4_X1M_A12TS oc8051_sfr1_u27 ( .A(oc8051_sfr1_psw_4_), .B(srcac), .C(
        oc8051_sfr1_psw_5_), .D(cy), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n11) );
  MXT4_X1M_A12TS oc8051_sfr1_u26 ( .A(oc8051_sfr1_psw_0_), .B(
        oc8051_sfr1_psw_2_), .C(oc8051_sfr1_psw_1_), .D(oc8051_sfr1_psw_3_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n10) );
  MXT2_X1M_A12TS oc8051_sfr1_u25 ( .A(oc8051_sfr1_n10), .B(oc8051_sfr1_n11), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1280) );
  MXT4_X1M_A12TS oc8051_sfr1_u24 ( .A(oc8051_sfr1_tr0), .B(oc8051_sfr1_tr1), 
        .C(oc8051_sfr1_tcon_5_), .D(oc8051_sfr1_tcon_7_), .S0(rd_addr[1]), 
        .S1(rd_addr[0]), .Y(oc8051_sfr1_n9) );
  MXT4_X1M_A12TS oc8051_sfr1_u23 ( .A(oc8051_sfr1_tcon_0_), .B(
        oc8051_sfr1_tcon_2_), .C(oc8051_sfr1_tcon_1_), .D(oc8051_sfr1_tcon_3_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n8) );
  MXT2_X1M_A12TS oc8051_sfr1_u22 ( .A(oc8051_sfr1_n8), .B(oc8051_sfr1_n9), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1360) );
  MXIT2_X0P7M_A12TS oc8051_sfr1_u21 ( .A(oc8051_sfr1_n212), .B(descy), .S0(
        oc8051_sfr1_n213), .Y(oc8051_sfr1_n7) );
  MXT2_X1M_A12TS oc8051_sfr1_u20 ( .A(oc8051_sfr1_n28), .B(oc8051_sfr1_n29), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n6) );
  MXIT2_X0P7M_A12TS oc8051_sfr1_u19 ( .A(oc8051_sfr1_n6), .B(oc8051_sfr1_n7), 
        .S0(oc8051_sfr1_n208), .Y(oc8051_sfr1_n1400) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u18 ( .A(oc8051_sfr1_n18), .B(oc8051_sfr1_n19), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1370) );
  MXT4_X1M_A12TS oc8051_sfr1_u17 ( .A(oc8051_sfr1_p3_data_4_), .B(
        oc8051_sfr1_p3_data_6_), .C(oc8051_sfr1_p3_data_5_), .D(
        oc8051_sfr1_p3_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n5) );
  MXT4_X1M_A12TS oc8051_sfr1_u16 ( .A(oc8051_sfr1_p3_data_0_), .B(
        oc8051_sfr1_p3_data_2_), .C(oc8051_sfr1_p3_data_1_), .D(
        oc8051_sfr1_p3_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n4) );
  MXT2_X1M_A12TS oc8051_sfr1_u15 ( .A(oc8051_sfr1_n4), .B(oc8051_sfr1_n5), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1320) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u14 ( .A(wr_dat[0]), .B(wr_dat[2]), .C(
        wr_dat[1]), .D(wr_dat[3]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n28) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u13 ( .A(oc8051_sfr1_p1_data_0_), .B(
        oc8051_sfr1_p1_data_2_), .C(oc8051_sfr1_p1_data_1_), .D(
        oc8051_sfr1_p1_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n26) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u12 ( .A(oc8051_sfr1_p2_data_4_), .B(
        oc8051_sfr1_p2_data_6_), .C(oc8051_sfr1_p2_data_5_), .D(
        oc8051_sfr1_p2_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n25) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u11 ( .A(oc8051_sfr1_p1_data_4_), .B(
        oc8051_sfr1_p1_data_6_), .C(oc8051_sfr1_p1_data_5_), .D(
        oc8051_sfr1_p1_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n27) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u10 ( .A(oc8051_sfr1_p2_data_0_), .B(
        oc8051_sfr1_p2_data_2_), .C(oc8051_sfr1_p2_data_1_), .D(
        oc8051_sfr1_p2_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n24) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u9 ( .A(oc8051_sfr1_n26), .B(oc8051_sfr1_n27), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1300) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u8 ( .A(oc8051_sfr1_n24), .B(oc8051_sfr1_n25), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1310) );
  MXT4_X1M_A12TS oc8051_sfr1_u7 ( .A(oc8051_sfr1_p0_data_4_), .B(
        oc8051_sfr1_p0_data_6_), .C(oc8051_sfr1_p0_data_5_), .D(
        oc8051_sfr1_p0_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n3) );
  MXT4_X1M_A12TS oc8051_sfr1_u6 ( .A(oc8051_sfr1_p0_data_0_), .B(
        oc8051_sfr1_p0_data_2_), .C(oc8051_sfr1_p0_data_1_), .D(
        oc8051_sfr1_p0_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n2) );
  MXT2_X1M_A12TS oc8051_sfr1_u5 ( .A(oc8051_sfr1_n2), .B(oc8051_sfr1_n3), .S0(
        rd_addr[2]), .Y(oc8051_sfr1_n1290) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u4 ( .A(wr_dat[4]), .B(wr_dat[6]), .C(
        wr_dat[5]), .D(wr_dat[7]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n29) );
  TIELO_X1M_A12TS oc8051_sfr1_u3 ( .Y(oc8051_sfr1_int_src_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_bit_out_reg ( .D(oc8051_sfr1_n1400), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_bit) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_wr_bit_r_reg ( .D(bit_addr_o), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_wr_bit_r) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_wait_data_reg ( .D(oc8051_sfr1_n1020), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(wait_data) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_pres_ow_reg ( .D(oc8051_sfr1_n259), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_pres_ow) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_2_ ( .D(oc8051_sfr1_n1510), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_0_ ( .D(oc8051_sfr1_n258), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_1_ ( .D(oc8051_sfr1_n1500), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_7_ ( .D(oc8051_sfr1_n237), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_6_ ( .D(oc8051_sfr1_n238), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_5_ ( .D(oc8051_sfr1_n239), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_4_ ( .D(oc8051_sfr1_n240), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_3_ ( .D(oc8051_sfr1_n241), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_2_ ( .D(oc8051_sfr1_n242), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_1_ ( .D(oc8051_sfr1_n243), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_0_ ( .D(oc8051_sfr1_n244), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_3_ ( .D(oc8051_sfr1_n1520), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_3_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u77 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_acc1_n61) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u76 ( .A(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_acc1_n60) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u75 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_acc1_n11) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u74 ( .A(
        oc8051_sfr1_oc8051_acc1_n61), .B(oc8051_sfr1_oc8051_acc1_n60), .C(
        oc8051_sfr1_oc8051_acc1_n11), .Y(oc8051_sfr1_oc8051_acc1_n62) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u73 ( .A(n_5_net_), .Y(
        oc8051_sfr1_oc8051_acc1_n66) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u72 ( .A(
        oc8051_sfr1_oc8051_acc1_n66), .B(wr_addr[4]), .C(wr_addr[3]), .Y(
        oc8051_sfr1_oc8051_acc1_n65) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u71 ( .A(wr_addr[6]), .B(
        wr_addr[5]), .C(wr_addr[7]), .D(oc8051_sfr1_oc8051_acc1_n65), .Y(
        oc8051_sfr1_oc8051_acc1_n63) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u70 ( .AN(wr_sfr[1]), .B(
        wr_sfr[0]), .Y(oc8051_sfr1_oc8051_acc1_n64) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u69 ( .A0(
        oc8051_sfr1_oc8051_acc1_n62), .A1(oc8051_sfr1_wr_bit_r), .A2(
        oc8051_sfr1_oc8051_acc1_n63), .B0(oc8051_sfr1_oc8051_acc1_n64), .Y(
        oc8051_sfr1_oc8051_acc1_n57) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u68 ( .AN(wr_sfr[1]), .B(wr_sfr[0]), .Y(oc8051_sfr1_oc8051_acc1_n9) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u67 ( .AN(
        oc8051_sfr1_oc8051_acc1_n63), .B(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_acc1_n59) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u66 ( .A(
        oc8051_sfr1_oc8051_acc1_n57), .B(oc8051_sfr1_oc8051_acc1_n9), .C(
        oc8051_sfr1_oc8051_acc1_n59), .Y(oc8051_sfr1_oc8051_acc1_n33) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u65 ( .A(descy), .B(
        oc8051_sfr1_oc8051_acc1_n33), .Y(oc8051_sfr1_oc8051_acc1_n19) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u64 ( .A(oc8051_sfr1_oc8051_acc1_n19), .Y(oc8051_sfr1_oc8051_acc1_n32) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u63 ( .A(oc8051_sfr1_oc8051_acc1_n62), .Y(oc8051_sfr1_oc8051_acc1_n53) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u62 ( .A0(
        oc8051_sfr1_oc8051_acc1_n32), .A1(oc8051_sfr1_oc8051_acc1_n53), .B0(
        des2[0]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n54) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u61 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_acc1_n60), .C(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_acc1_n49) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u60 ( .A(
        oc8051_sfr1_oc8051_acc1_n11), .B(oc8051_sfr1_oc8051_acc1_n60), .C(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_acc1_n45) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u59 ( .A(
        oc8051_sfr1_oc8051_acc1_n61), .B(oc8051_sfr1_oc8051_acc1_n60), .C(
        wr_addr[0]), .Y(oc8051_sfr1_oc8051_acc1_n47) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u58 ( .A(
        oc8051_sfr1_oc8051_acc1_n49), .B(oc8051_sfr1_oc8051_acc1_n45), .C(
        oc8051_sfr1_oc8051_acc1_n47), .Y(oc8051_sfr1_oc8051_acc1_n34) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u57 ( .A(
        oc8051_sfr1_oc8051_acc1_n11), .B(oc8051_sfr1_oc8051_acc1_n61), .C(
        wr_addr[2]), .Y(oc8051_sfr1_oc8051_acc1_n46) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u56 ( .A(oc8051_sfr1_oc8051_acc1_n46), .Y(oc8051_sfr1_oc8051_acc1_n31) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u55 ( .A(
        oc8051_sfr1_oc8051_acc1_n34), .B(oc8051_sfr1_oc8051_acc1_n31), .Y(
        oc8051_sfr1_oc8051_acc1_n24) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u54 ( .A(oc8051_sfr1_oc8051_acc1_n33), .Y(oc8051_sfr1_oc8051_acc1_n25) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u53 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_acc1_n33), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_acc1_n23) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u52 ( .A(
        oc8051_sfr1_oc8051_acc1_n60), .B(wr_addr[1]), .C(
        oc8051_sfr1_oc8051_acc1_n11), .Y(oc8051_sfr1_oc8051_acc1_n27) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u51 ( .A(oc8051_sfr1_oc8051_acc1_n59), .Y(oc8051_sfr1_oc8051_acc1_n58) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u50 ( .A(
        oc8051_sfr1_oc8051_acc1_n58), .B(oc8051_sfr1_oc8051_acc1_n9), .C(
        oc8051_sfr1_oc8051_acc1_n57), .Y(oc8051_sfr1_oc8051_acc1_n22) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u49 ( .A0(
        oc8051_sfr1_oc8051_acc1_n33), .A1(oc8051_sfr1_oc8051_acc1_n27), .B0(
        oc8051_sfr1_oc8051_acc1_n22), .Y(oc8051_sfr1_oc8051_acc1_n17) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u48 ( .A0(
        oc8051_sfr1_oc8051_acc1_n24), .A1(oc8051_sfr1_oc8051_acc1_n25), .B0(
        oc8051_sfr1_oc8051_acc1_n23), .C0(oc8051_sfr1_oc8051_acc1_n17), .Y(
        oc8051_sfr1_oc8051_acc1_n56) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u47 ( .AN(
        oc8051_sfr1_oc8051_acc1_n57), .B(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n8) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u46 ( .A0(acc[0]), .A1(
        oc8051_sfr1_oc8051_acc1_n56), .B0(des_acc[0]), .B1(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n55) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u45 ( .A(
        oc8051_sfr1_oc8051_acc1_n54), .B(oc8051_sfr1_oc8051_acc1_n55), .Y(
        oc8051_sfr1_oc8051_acc1_acc_0_) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u44 ( .A(
        oc8051_sfr1_oc8051_acc1_n49), .B(oc8051_sfr1_oc8051_acc1_n45), .C(
        oc8051_sfr1_oc8051_acc1_n46), .Y(oc8051_sfr1_oc8051_acc1_n52) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u43 ( .A(
        oc8051_sfr1_oc8051_acc1_n33), .B(oc8051_sfr1_oc8051_acc1_n53), .Y(
        oc8051_sfr1_oc8051_acc1_n26) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u42 ( .A(
        oc8051_sfr1_oc8051_acc1_n26), .B(oc8051_sfr1_oc8051_acc1_n23), .C(
        oc8051_sfr1_oc8051_acc1_n17), .Y(oc8051_sfr1_oc8051_acc1_n35) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u41 ( .A0(
        oc8051_sfr1_oc8051_acc1_n33), .A1(oc8051_sfr1_oc8051_acc1_n52), .B0(
        oc8051_sfr1_oc8051_acc1_n35), .C0(acc[1]), .Y(
        oc8051_sfr1_oc8051_acc1_n50) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u40 ( .A0(des_acc[1]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[1]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n51) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u39 ( .A0(
        oc8051_sfr1_oc8051_acc1_n19), .A1(oc8051_sfr1_oc8051_acc1_n47), .B0(
        oc8051_sfr1_oc8051_acc1_n50), .C0(oc8051_sfr1_oc8051_acc1_n51), .Y(
        oc8051_sfr1_oc8051_acc1_acc_1_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u38 ( .A(des_acc[2]), .B(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n42) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u37 ( .A(oc8051_sfr1_oc8051_acc1_n49), .Y(oc8051_sfr1_oc8051_acc1_n39) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u36 ( .A(oc8051_sfr1_oc8051_acc1_n35), .Y(oc8051_sfr1_oc8051_acc1_n48) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u35 ( .A0(
        oc8051_sfr1_oc8051_acc1_n46), .A1(oc8051_sfr1_oc8051_acc1_n47), .B0(
        oc8051_sfr1_oc8051_acc1_n25), .C0(oc8051_sfr1_oc8051_acc1_n48), .Y(
        oc8051_sfr1_oc8051_acc1_n41) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u34 ( .A0(
        oc8051_sfr1_oc8051_acc1_n39), .A1(oc8051_sfr1_oc8051_acc1_n33), .B0(
        oc8051_sfr1_oc8051_acc1_n41), .C0(acc[2]), .Y(
        oc8051_sfr1_oc8051_acc1_n43) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u33 ( .A(oc8051_sfr1_oc8051_acc1_n45), .Y(oc8051_sfr1_oc8051_acc1_n40) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u32 ( .A0(
        oc8051_sfr1_oc8051_acc1_n32), .A1(oc8051_sfr1_oc8051_acc1_n40), .B0(
        des2[2]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n44) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u31 ( .A(
        oc8051_sfr1_oc8051_acc1_n42), .B(oc8051_sfr1_oc8051_acc1_n43), .C(
        oc8051_sfr1_oc8051_acc1_n44), .Y(oc8051_sfr1_oc8051_acc1_acc_2_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u30 ( .A(des_acc[3]), .B(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n36) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u29 ( .A0(
        oc8051_sfr1_oc8051_acc1_n40), .A1(oc8051_sfr1_oc8051_acc1_n33), .B0(
        oc8051_sfr1_oc8051_acc1_n41), .C0(acc[3]), .Y(
        oc8051_sfr1_oc8051_acc1_n37) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u28 ( .A0(
        oc8051_sfr1_oc8051_acc1_n39), .A1(oc8051_sfr1_oc8051_acc1_n32), .B0(
        des2[3]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n38) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u27 ( .A(
        oc8051_sfr1_oc8051_acc1_n36), .B(oc8051_sfr1_oc8051_acc1_n37), .C(
        oc8051_sfr1_oc8051_acc1_n38), .Y(oc8051_sfr1_oc8051_acc1_acc_3_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u26 ( .A(des_acc[4]), .B(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n28) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u25 ( .A0(
        oc8051_sfr1_oc8051_acc1_n33), .A1(oc8051_sfr1_oc8051_acc1_n34), .B0(
        oc8051_sfr1_oc8051_acc1_n35), .C0(acc[4]), .Y(
        oc8051_sfr1_oc8051_acc1_n29) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u24 ( .A0(
        oc8051_sfr1_oc8051_acc1_n31), .A1(oc8051_sfr1_oc8051_acc1_n32), .B0(
        des2[4]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n30) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u23 ( .A(
        oc8051_sfr1_oc8051_acc1_n28), .B(oc8051_sfr1_oc8051_acc1_n29), .C(
        oc8051_sfr1_oc8051_acc1_n30), .Y(oc8051_sfr1_oc8051_acc1_acc_4_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u22 ( .A(oc8051_sfr1_oc8051_acc1_n27), .Y(oc8051_sfr1_oc8051_acc1_n18) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u21 ( .A0(
        oc8051_sfr1_oc8051_acc1_n24), .A1(oc8051_sfr1_oc8051_acc1_n25), .B0(
        oc8051_sfr1_oc8051_acc1_n26), .Y(oc8051_sfr1_oc8051_acc1_n16) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u20 ( .A(oc8051_sfr1_oc8051_acc1_n23), .Y(oc8051_sfr1_oc8051_acc1_n10) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u19 ( .A0(
        oc8051_sfr1_oc8051_acc1_n16), .A1(oc8051_sfr1_oc8051_acc1_n10), .A2(
        oc8051_sfr1_oc8051_acc1_n22), .B0(acc[5]), .Y(
        oc8051_sfr1_oc8051_acc1_n20) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u18 ( .A0(des_acc[5]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[5]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n21) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u17 ( .A0(
        oc8051_sfr1_oc8051_acc1_n18), .A1(oc8051_sfr1_oc8051_acc1_n19), .B0(
        oc8051_sfr1_oc8051_acc1_n20), .C0(oc8051_sfr1_oc8051_acc1_n21), .Y(
        oc8051_sfr1_oc8051_acc1_acc_5_) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u16 ( .AN(
        oc8051_sfr1_oc8051_acc1_n16), .B(oc8051_sfr1_oc8051_acc1_n17), .Y(
        oc8051_sfr1_oc8051_acc1_n12) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u15 ( .A0(
        oc8051_sfr1_oc8051_acc1_n10), .A1(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_acc1_n12), .C0(acc[6]), .Y(
        oc8051_sfr1_oc8051_acc1_n13) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u14 ( .A(descy), .B(
        oc8051_sfr1_oc8051_acc1_n11), .C(oc8051_sfr1_oc8051_acc1_n10), .Y(
        oc8051_sfr1_oc8051_acc1_n14) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u13 ( .A0(des_acc[6]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[6]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n15) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u12 ( .A(
        oc8051_sfr1_oc8051_acc1_n13), .B(oc8051_sfr1_oc8051_acc1_n14), .C(
        oc8051_sfr1_oc8051_acc1_n15), .Y(oc8051_sfr1_oc8051_acc1_acc_6_) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u11 ( .A0(
        oc8051_sfr1_oc8051_acc1_n10), .A1(oc8051_sfr1_oc8051_acc1_n11), .B0(
        oc8051_sfr1_oc8051_acc1_n12), .C0(acc[7]), .Y(
        oc8051_sfr1_oc8051_acc1_n5) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u10 ( .A(descy), .B(wr_addr[0]), 
        .C(oc8051_sfr1_oc8051_acc1_n10), .Y(oc8051_sfr1_oc8051_acc1_n6) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u9 ( .A0(des_acc[7]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[7]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n7) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u8 ( .A(oc8051_sfr1_oc8051_acc1_n5), .B(oc8051_sfr1_oc8051_acc1_n6), .C(oc8051_sfr1_oc8051_acc1_n7), .Y(
        oc8051_sfr1_oc8051_acc1_acc_7_) );
  XNOR2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u7 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_1_), .B(oc8051_sfr1_oc8051_acc1_acc_0_), 
        .Y(oc8051_sfr1_oc8051_acc1_n4) );
  XNOR3_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u6 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_2_), .B(oc8051_sfr1_oc8051_acc1_acc_3_), 
        .C(oc8051_sfr1_oc8051_acc1_n4), .Y(oc8051_sfr1_oc8051_acc1_n1) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u5 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_5_), .B(oc8051_sfr1_oc8051_acc1_acc_4_), 
        .Y(oc8051_sfr1_oc8051_acc1_n3) );
  XOR3_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u4 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_7_), .B(oc8051_sfr1_oc8051_acc1_n3), .C(
        oc8051_sfr1_oc8051_acc1_acc_6_), .Y(oc8051_sfr1_oc8051_acc1_n2) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u3 ( .A(oc8051_sfr1_oc8051_acc1_n1), 
        .B(oc8051_sfr1_oc8051_acc1_n2), .Y(oc8051_sfr1_psw_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_0_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_2_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_6_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_1_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_4_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_3_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_7_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_5_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[5]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_b_register_u37 ( .A(oc8051_sfr1_wr_bit_r), 
        .Y(oc8051_sfr1_oc8051_b_register_n5) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u36 ( .AN(wr_addr[4]), .B(
        wr_addr[3]), .Y(oc8051_sfr1_oc8051_b_register_n28) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u35 ( .A(wr_addr[7]), .B(
        wr_addr[6]), .C(oc8051_sfr1_oc8051_b_register_n28), .D(wr_addr[5]), 
        .Y(oc8051_sfr1_oc8051_b_register_n25) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u34 ( .A(
        oc8051_sfr1_oc8051_b_register_n25), .B(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_b_register_n27) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_b_register_u33 ( .A(descy), .B(
        oc8051_sfr1_oc8051_b_register_n27), .Y(
        oc8051_sfr1_oc8051_b_register_n6) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u32 ( .B0(des_acc[0]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n23) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_b_register_u31 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_b_register_n9) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_b_register_u30 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_b_register_n12) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u29 ( .A(n_5_net_), .B(
        oc8051_sfr1_oc8051_b_register_n27), .Y(
        oc8051_sfr1_oc8051_b_register_n15) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u28 ( .AN(
        oc8051_sfr1_oc8051_b_register_n15), .B(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_b_register_n18) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_b_register_u27 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_wr_bit_r), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_b_register_n26) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u26 ( .A(
        oc8051_sfr1_oc8051_b_register_n25), .B(
        oc8051_sfr1_oc8051_b_register_n9), .C(n_5_net_), .D(
        oc8051_sfr1_oc8051_b_register_n26), .Y(
        oc8051_sfr1_oc8051_b_register_n4) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u25 ( .A0(
        oc8051_sfr1_oc8051_b_register_n9), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(
        oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n24) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u24 ( .A(
        oc8051_sfr1_oc8051_b_register_n23), .B(oc8051_sfr1_b_reg_0_), .S0(
        oc8051_sfr1_oc8051_b_register_n24), .Y(
        oc8051_sfr1_oc8051_b_register_n32) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u23 ( .B0(des_acc[1]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n21) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u22 ( .A0(wr_addr[0]), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(
        oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n22) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u21 ( .A(
        oc8051_sfr1_oc8051_b_register_n21), .B(oc8051_sfr1_b_reg_1_), .S0(
        oc8051_sfr1_oc8051_b_register_n22), .Y(
        oc8051_sfr1_oc8051_b_register_n33) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u20 ( .B0(des_acc[2]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n19) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u19 ( .A0(wr_addr[1]), .A1(
        oc8051_sfr1_oc8051_b_register_n9), .A2(
        oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n20) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u18 ( .A(
        oc8051_sfr1_oc8051_b_register_n19), .B(oc8051_sfr1_b_reg_2_), .S0(
        oc8051_sfr1_oc8051_b_register_n20), .Y(
        oc8051_sfr1_oc8051_b_register_n34) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u17 ( .B0(des_acc[3]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n16) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u16 ( .A0(wr_addr[1]), .A1(
        wr_addr[0]), .A2(oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n17) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u15 ( .A(
        oc8051_sfr1_oc8051_b_register_n16), .B(oc8051_sfr1_b_reg_3_), .S0(
        oc8051_sfr1_oc8051_b_register_n17), .Y(
        oc8051_sfr1_oc8051_b_register_n35) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u14 ( .B0(des_acc[4]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n13) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u13 ( .A(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_b_register_n15), .Y(
        oc8051_sfr1_oc8051_b_register_n3) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u12 ( .A0(
        oc8051_sfr1_oc8051_b_register_n9), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(
        oc8051_sfr1_oc8051_b_register_n3), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n14) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u11 ( .A(
        oc8051_sfr1_oc8051_b_register_n13), .B(oc8051_sfr1_b_reg_4_), .S0(
        oc8051_sfr1_oc8051_b_register_n14), .Y(
        oc8051_sfr1_oc8051_b_register_n36) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u10 ( .B0(des_acc[5]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n10) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u9 ( .A0(
        oc8051_sfr1_oc8051_b_register_n3), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n11) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u8 ( .A(
        oc8051_sfr1_oc8051_b_register_n10), .B(oc8051_sfr1_b_reg_5_), .S0(
        oc8051_sfr1_oc8051_b_register_n11), .Y(
        oc8051_sfr1_oc8051_b_register_n37) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u7 ( .B0(des_acc[6]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(oc8051_sfr1_oc8051_b_register_n7) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u6 ( .A0(
        oc8051_sfr1_oc8051_b_register_n3), .A1(
        oc8051_sfr1_oc8051_b_register_n9), .A2(wr_addr[1]), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(oc8051_sfr1_oc8051_b_register_n8) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u5 ( .A(
        oc8051_sfr1_oc8051_b_register_n7), .B(oc8051_sfr1_b_reg_6_), .S0(
        oc8051_sfr1_oc8051_b_register_n8), .Y(
        oc8051_sfr1_oc8051_b_register_n38) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u4 ( .B0(des_acc[7]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(oc8051_sfr1_oc8051_b_register_n1) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u3 ( .A0(wr_addr[0]), .A1(
        oc8051_sfr1_oc8051_b_register_n3), .A2(wr_addr[1]), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(oc8051_sfr1_oc8051_b_register_n2) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u2 ( .A(
        oc8051_sfr1_oc8051_b_register_n1), .B(oc8051_sfr1_b_reg_7_), .S0(
        oc8051_sfr1_oc8051_b_register_n2), .Y(
        oc8051_sfr1_oc8051_b_register_n39) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_b_register_n34), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_b_register_n38), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_b_register_n32), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_b_register_n36), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_b_register_n33), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_b_register_n37), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_b_register_n35), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_b_register_n39), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_7_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u34 ( .A(ram_rd_sel[2]), .Y(
        oc8051_sfr1_oc8051_sp1_n4) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u33 ( .A(oc8051_sfr1_oc8051_sp1_n4), 
        .B(ram_rd_sel[0]), .C(ram_rd_sel[1]), .Y(oc8051_sfr1_oc8051_sp1_n22)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u32 ( .A(wb_rst_i), .Y(
        oc8051_sfr1_oc8051_sp1_n5) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_sp1_u31 ( .A(oc8051_sfr1_oc8051_sp1_pop), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(oc8051_sfr1_oc8051_sp1_r313_b_as_0_) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_sp1_u30 ( .A(wr_addr[2]), .B(wr_addr[1]), 
        .Y(oc8051_sfr1_oc8051_sp1_n3) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_sp1_u29 ( .A(wr_addr[7]), .B(wr_addr[0]), .C(oc8051_sfr1_oc8051_sp1_n3), .D(n_5_net_), .Y(oc8051_sfr1_oc8051_sp1_n2)
         );
  OR6_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u28 ( .A(oc8051_sfr1_wr_bit_r), .B(
        wr_addr[6]), .C(wr_addr[5]), .D(wr_addr[4]), .E(wr_addr[3]), .F(
        oc8051_sfr1_oc8051_sp1_n2), .Y(oc8051_sfr1_oc8051_sp1_n1) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u27 ( .A(wr_dat[0]), .B(
        oc8051_sfr1_oc8051_sp1_n24), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[0])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u26 ( .A(wr_dat[1]), .B(
        oc8051_sfr1_oc8051_sp1_n25), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[1])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u25 ( .A(wr_dat[2]), .B(
        oc8051_sfr1_oc8051_sp1_n26), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[2])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u24 ( .A(wr_dat[3]), .B(
        oc8051_sfr1_oc8051_sp1_n27), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[3])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u23 ( .A(wr_dat[4]), .B(
        oc8051_sfr1_oc8051_sp1_n28), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[4])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u22 ( .A(wr_dat[5]), .B(
        oc8051_sfr1_oc8051_sp1_n29), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[5])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u21 ( .A(wr_dat[6]), .B(
        oc8051_sfr1_oc8051_sp1_n30), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[6])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u20 ( .A(wr_dat[7]), .B(
        oc8051_sfr1_oc8051_sp1_n31), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(sp[7])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u19 ( .A(wr_dat[0]), .B(
        oc8051_sfr1_oc8051_sp1_sp_0_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[0]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u18 ( .A(wr_dat[1]), .B(
        oc8051_sfr1_oc8051_sp1_sp_1_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[1]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u17 ( .A(wr_dat[2]), .B(
        oc8051_sfr1_oc8051_sp1_sp_2_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[2]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u16 ( .A(wr_dat[3]), .B(
        oc8051_sfr1_oc8051_sp1_sp_3_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[3]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u15 ( .A(wr_dat[4]), .B(
        oc8051_sfr1_oc8051_sp1_sp_4_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[4]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u14 ( .A(wr_dat[5]), .B(
        oc8051_sfr1_oc8051_sp1_sp_5_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[5]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u13 ( .A(wr_dat[6]), .B(
        oc8051_sfr1_oc8051_sp1_sp_6_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[6]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u12 ( .A(wr_dat[7]), .B(
        oc8051_sfr1_oc8051_sp1_sp_7_), .S0(oc8051_sfr1_oc8051_sp1_n1), .Y(
        oc8051_sfr1_oc8051_sp1_sp_t[7]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u11 ( .A(oc8051_sfr1_oc8051_sp1_n13), 
        .B(oc8051_sfr1_oc8051_sp1_sp_0_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[0]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u10 ( .A(oc8051_sfr1_oc8051_sp1_n14), 
        .B(oc8051_sfr1_oc8051_sp1_sp_1_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[1]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u9 ( .A(oc8051_sfr1_oc8051_sp1_n15), 
        .B(oc8051_sfr1_oc8051_sp1_sp_2_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[2]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u8 ( .A(oc8051_sfr1_oc8051_sp1_n16), 
        .B(oc8051_sfr1_oc8051_sp1_sp_3_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[3]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u7 ( .A(oc8051_sfr1_oc8051_sp1_n17), 
        .B(oc8051_sfr1_oc8051_sp1_sp_4_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[4]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u6 ( .A(oc8051_sfr1_oc8051_sp1_n18), 
        .B(oc8051_sfr1_oc8051_sp1_sp_5_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[5]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u5 ( .A(oc8051_sfr1_oc8051_sp1_n19), 
        .B(oc8051_sfr1_oc8051_sp1_sp_6_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[6]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u4 ( .A(oc8051_sfr1_oc8051_sp1_n20), 
        .B(oc8051_sfr1_oc8051_sp1_sp_7_), .S0(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .Y(sp_w[7]) );
  NAND3B_X1M_A12TS oc8051_sfr1_oc8051_sp1_u3 ( .AN(ram_wr_sel[2]), .B(
        ram_wr_sel[0]), .C(ram_wr_sel[1]), .Y(oc8051_sfr1_oc8051_sp1_u3_u2_z_0) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_0_ ( .D(sp[0]), .CK(wb_clk_i), 
        .SN(oc8051_sfr1_oc8051_sp1_n5), .Q(oc8051_sfr1_oc8051_sp1_sp_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_6_ ( .D(sp[6]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_5_ ( .D(sp[5]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_4_ ( .D(sp[4]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_3_ ( .D(sp[3]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_3_) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_2_ ( .D(sp[2]), .CK(wb_clk_i), 
        .SN(oc8051_sfr1_oc8051_sp1_n5), .Q(oc8051_sfr1_oc8051_sp1_sp_2_) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_1_ ( .D(sp[1]), .CK(wb_clk_i), 
        .SN(oc8051_sfr1_oc8051_sp1_n5), .Q(oc8051_sfr1_oc8051_sp1_sp_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_7_ ( .D(sp[7]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_pop_reg ( .D(
        oc8051_sfr1_oc8051_sp1_n22), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_sp1_pop) );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_7 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[7]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_7_), .CO(), .S(
        oc8051_sfr1_oc8051_sp1_n31) );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_6 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[6]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_6_), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_7_), .S(oc8051_sfr1_oc8051_sp1_n30)
         );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_5 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[5]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_5_), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_6_), .S(oc8051_sfr1_oc8051_sp1_n29)
         );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_4 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[4]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_4_), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_5_), .S(oc8051_sfr1_oc8051_sp1_n28)
         );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_3 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[3]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_3_), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_4_), .S(oc8051_sfr1_oc8051_sp1_n27)
         );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_2 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[2]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_2_), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_3_), .S(oc8051_sfr1_oc8051_sp1_n26)
         );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_1 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[1]), .B(oc8051_sfr1_oc8051_sp1_u3_u2_z_0), 
        .CI(oc8051_sfr1_oc8051_sp1_r313_carry_1_), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_2_), .S(oc8051_sfr1_oc8051_sp1_n25)
         );
  ADDF_X1M_A12TS oc8051_sfr1_oc8051_sp1_r313_u1_0 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_t[0]), .B(
        oc8051_sfr1_oc8051_sp1_r313_b_as_0_), .CI(
        oc8051_sfr1_oc8051_sp1_u3_u2_z_0), .CO(
        oc8051_sfr1_oc8051_sp1_r313_carry_1_), .S(oc8051_sfr1_oc8051_sp1_n24)
         );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u2 ( .A(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[7]), .B(
        oc8051_sfr1_oc8051_sp1_sp_7_), .Y(oc8051_sfr1_oc8051_sp1_n20) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_0_), .Y(oc8051_sfr1_oc8051_sp1_n13) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_1 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_1_), .B(oc8051_sfr1_oc8051_sp1_sp_0_), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[2]), .S(
        oc8051_sfr1_oc8051_sp1_n14) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_5 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_5_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[5]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[6]), .S(
        oc8051_sfr1_oc8051_sp1_n18) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_4 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_4_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[4]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[5]), .S(
        oc8051_sfr1_oc8051_sp1_n17) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_3 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_3_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[3]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[4]), .S(
        oc8051_sfr1_oc8051_sp1_n16) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_2 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_2_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[2]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[3]), .S(
        oc8051_sfr1_oc8051_sp1_n15) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_6 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_6_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[6]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[7]), .S(
        oc8051_sfr1_oc8051_sp1_n19) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u32 ( .A(wr_sfr[1]), .B(wr_sfr[0]), 
        .Y(oc8051_sfr1_oc8051_dptr1_n4) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u31 ( .AN(wr_addr[2]), .B(
        wr_addr[1]), .C(n_5_net_), .D(wr_addr[7]), .Y(
        oc8051_sfr1_oc8051_dptr1_n15) );
  OR6_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u30 ( .A(oc8051_sfr1_wr_bit_r), .B(
        wr_addr[6]), .C(wr_addr[5]), .D(wr_addr[4]), .E(wr_addr[3]), .F(
        oc8051_sfr1_oc8051_dptr1_n15), .Y(oc8051_sfr1_oc8051_dptr1_n2) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_dptr1_u29 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_dptr1_n3) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_dptr1_u28 ( .A(
        oc8051_sfr1_oc8051_dptr1_n2), .B(oc8051_sfr1_oc8051_dptr1_n4), .C(
        oc8051_sfr1_oc8051_dptr1_n3), .Y(oc8051_sfr1_oc8051_dptr1_n7) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_dptr1_u27 ( .A(
        oc8051_sfr1_oc8051_dptr1_n4), .B(oc8051_sfr1_oc8051_dptr1_n7), .Y(
        oc8051_sfr1_oc8051_dptr1_n6) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u26 ( .A0(dptr_hi[0]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[0]), .Y(oc8051_sfr1_oc8051_dptr1_n14) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u25 ( .B0(des2[0]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n14), .Y(
        oc8051_sfr1_oc8051_dptr1_n18) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u24 ( .A0(dptr_hi[1]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[1]), .Y(oc8051_sfr1_oc8051_dptr1_n13) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u23 ( .B0(des2[1]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n13), .Y(
        oc8051_sfr1_oc8051_dptr1_n19) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u22 ( .A0(dptr_hi[2]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[2]), .Y(oc8051_sfr1_oc8051_dptr1_n12) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u21 ( .B0(des2[2]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n12), .Y(
        oc8051_sfr1_oc8051_dptr1_n20) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u20 ( .A0(dptr_hi[3]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[3]), .Y(oc8051_sfr1_oc8051_dptr1_n11) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u19 ( .B0(des2[3]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n11), .Y(
        oc8051_sfr1_oc8051_dptr1_n21) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u18 ( .A0(dptr_hi[4]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[4]), .Y(oc8051_sfr1_oc8051_dptr1_n10) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u17 ( .B0(des2[4]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n10), .Y(
        oc8051_sfr1_oc8051_dptr1_n22) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u16 ( .A0(dptr_hi[5]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[5]), .Y(oc8051_sfr1_oc8051_dptr1_n9) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u15 ( .B0(des2[5]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n9), .Y(
        oc8051_sfr1_oc8051_dptr1_n23) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u14 ( .A0(dptr_hi[6]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[6]), .Y(oc8051_sfr1_oc8051_dptr1_n8) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u13 ( .B0(des2[6]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n8), .Y(
        oc8051_sfr1_oc8051_dptr1_n24) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u12 ( .A0(dptr_hi[7]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[7]), .Y(oc8051_sfr1_oc8051_dptr1_n5) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u11 ( .B0(des2[7]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n5), .Y(
        oc8051_sfr1_oc8051_dptr1_n25) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u10 ( .A1N(
        oc8051_sfr1_oc8051_dptr1_n2), .A0(oc8051_sfr1_oc8051_dptr1_n3), .B0(
        oc8051_sfr1_oc8051_dptr1_n4), .Y(oc8051_sfr1_oc8051_dptr1_n1) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u9 ( .A(des_acc[0]), .B(dptr_lo[0]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n26) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u8 ( .A(des_acc[1]), .B(dptr_lo[1]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n27) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u7 ( .A(des_acc[2]), .B(dptr_lo[2]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n28) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u6 ( .A(des_acc[3]), .B(dptr_lo[3]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n29) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u5 ( .A(des_acc[4]), .B(dptr_lo[4]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n30) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u4 ( .A(des_acc[5]), .B(dptr_lo[5]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n31) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u3 ( .A(des_acc[6]), .B(dptr_lo[6]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n32) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u2 ( .A(des_acc[7]), .B(dptr_lo[7]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n33) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_0_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n18), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_1_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n19), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_2_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n20), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_3_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n21), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_4_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n22), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_5_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n23), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_6_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n24), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_7_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n25), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_0_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n26), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_1_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n27), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_2_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n28), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_3_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n29), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_4_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n30), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_5_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n31), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_6_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n32), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_7_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n33), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[7]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u51 ( .A(n_5_net_), .Y(
        oc8051_sfr1_oc8051_psw1_n40) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u50 ( .A(
        oc8051_sfr1_oc8051_psw1_n40), .B(wr_addr[5]), .C(wr_addr[3]), .Y(
        oc8051_sfr1_oc8051_psw1_n39) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u49 ( .A(wr_addr[6]), .B(wr_addr[4]), .C(wr_addr[7]), .D(oc8051_sfr1_oc8051_psw1_n39), .Y(
        oc8051_sfr1_oc8051_psw1_n37) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u48 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_psw1_n10) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u47 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_wr_bit_r), .C(wr_addr[2]), .Y(oc8051_sfr1_oc8051_psw1_n38)
         );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u46 ( .A(
        oc8051_sfr1_oc8051_psw1_n37), .B(oc8051_sfr1_oc8051_psw1_n10), .C(
        oc8051_sfr1_oc8051_psw1_n38), .Y(oc8051_sfr1_oc8051_psw1_n16) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u45 ( .A(wr_dat[4]), .B(
        oc8051_sfr1_psw_4_), .S0(oc8051_sfr1_oc8051_psw1_n16), .Y(bank_sel[1])
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u44 ( .A(oc8051_sfr1_oc8051_psw1_n16), .Y(oc8051_sfr1_oc8051_psw1_n7) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u43 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_psw1_n37), .Y(oc8051_sfr1_oc8051_psw1_n36) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u42 ( .A(oc8051_sfr1_oc8051_psw1_n36), .Y(oc8051_sfr1_oc8051_psw1_n24) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u41 ( .A(descy), .B(
        oc8051_sfr1_oc8051_psw1_n24), .Y(oc8051_sfr1_oc8051_psw1_n20) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u40 ( .B0(wr_dat[1]), .B1(
        oc8051_sfr1_oc8051_psw1_n7), .A0N(oc8051_sfr1_oc8051_psw1_n20), .Y(
        oc8051_sfr1_oc8051_psw1_n34) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u39 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_psw1_n8) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u38 ( .A(
        oc8051_sfr1_oc8051_psw1_n36), .B(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_psw1_n28) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u37 ( .A0(wr_addr[0]), .A1(
        oc8051_sfr1_oc8051_psw1_n8), .A2(oc8051_sfr1_oc8051_psw1_n28), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n35) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u36 ( .A(
        oc8051_sfr1_oc8051_psw1_n34), .B(oc8051_sfr1_psw_1_), .S0(
        oc8051_sfr1_oc8051_psw1_n35), .Y(oc8051_sfr1_oc8051_psw1_n43) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u35 ( .B0(wr_dat[2]), .B1(
        oc8051_sfr1_oc8051_psw1_n7), .A0N(oc8051_sfr1_oc8051_psw1_n20), .Y(
        oc8051_sfr1_oc8051_psw1_n31) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u34 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_psw1_n8), .Y(oc8051_sfr1_oc8051_psw1_n33) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u33 ( .A(oc8051_sfr1_oc8051_psw1_n7), .B(oc8051_sfr1_oc8051_psw1_n24), .Y(oc8051_sfr1_oc8051_psw1_n6) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u32 ( .A(oc8051_sfr1_oc8051_psw1_n6), .B(psw_set[1]), .Y(oc8051_sfr1_oc8051_psw1_n14) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u31 ( .A0(
        oc8051_sfr1_oc8051_psw1_n33), .A1(oc8051_sfr1_oc8051_psw1_n28), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .C0(oc8051_sfr1_oc8051_psw1_n14), .Y(
        oc8051_sfr1_oc8051_psw1_n32) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u30 ( .A(
        oc8051_sfr1_oc8051_psw1_n31), .B(oc8051_sfr1_psw_2_), .S0(
        oc8051_sfr1_oc8051_psw1_n32), .Y(oc8051_sfr1_oc8051_psw1_n29) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u29 ( .A(
        oc8051_sfr1_oc8051_psw1_n6), .B(psw_set[1]), .C(desov), .Y(
        oc8051_sfr1_oc8051_psw1_n30) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u28 ( .A(
        oc8051_sfr1_oc8051_psw1_n29), .B(oc8051_sfr1_oc8051_psw1_n30), .Y(
        oc8051_sfr1_oc8051_psw1_n44) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u27 ( .A(oc8051_sfr1_oc8051_psw1_n20), .Y(oc8051_sfr1_oc8051_psw1_n11) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u26 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_psw1_n7), .B0(oc8051_sfr1_oc8051_psw1_n11), .Y(
        oc8051_sfr1_oc8051_psw1_n25) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u25 ( .A(oc8051_sfr1_psw_3_), .Y(
        oc8051_sfr1_oc8051_psw1_n26) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u24 ( .A0(wr_addr[1]), .A1(
        wr_addr[0]), .A2(oc8051_sfr1_oc8051_psw1_n28), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n27) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u23 ( .A(
        oc8051_sfr1_oc8051_psw1_n25), .B(oc8051_sfr1_oc8051_psw1_n26), .S0(
        oc8051_sfr1_oc8051_psw1_n27), .Y(oc8051_sfr1_oc8051_psw1_n45) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u22 ( .A(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_psw1_n24), .Y(oc8051_sfr1_oc8051_psw1_n9) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u21 ( .A(oc8051_sfr1_oc8051_psw1_n9), .B(wr_addr[1]), .Y(oc8051_sfr1_oc8051_psw1_n19) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u20 ( .A(
        oc8051_sfr1_oc8051_psw1_n19), .B(oc8051_sfr1_oc8051_psw1_n10), .Y(
        oc8051_sfr1_oc8051_psw1_n21) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u19 ( .A(
        oc8051_sfr1_oc8051_psw1_n21), .B(oc8051_sfr1_psw_4_), .Y(
        oc8051_sfr1_oc8051_psw1_n23) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u18 ( .A(
        oc8051_sfr1_oc8051_psw1_n23), .B(wr_dat[4]), .S0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n22) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u17 ( .A0(
        oc8051_sfr1_oc8051_psw1_n21), .A1(oc8051_sfr1_oc8051_psw1_n20), .B0(
        oc8051_sfr1_oc8051_psw1_n22), .Y(oc8051_sfr1_oc8051_psw1_n46) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u16 ( .B0(wr_dat[5]), .B1(
        oc8051_sfr1_oc8051_psw1_n7), .A0N(oc8051_sfr1_oc8051_psw1_n20), .Y(
        oc8051_sfr1_oc8051_psw1_n17) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u15 ( .A0(
        oc8051_sfr1_oc8051_psw1_n19), .A1(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n18) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u14 ( .A(
        oc8051_sfr1_oc8051_psw1_n17), .B(oc8051_sfr1_psw_5_), .S0(
        oc8051_sfr1_oc8051_psw1_n18), .Y(oc8051_sfr1_oc8051_psw1_n47) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u13 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_psw1_n7), .B0(desac), .B1(
        oc8051_sfr1_oc8051_psw1_n6), .C0(oc8051_sfr1_oc8051_psw1_n11), .Y(
        oc8051_sfr1_oc8051_psw1_n12) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u12 ( .A0(
        oc8051_sfr1_oc8051_psw1_n8), .A1(wr_addr[0]), .A2(
        oc8051_sfr1_oc8051_psw1_n9), .B0(oc8051_sfr1_oc8051_psw1_n16), .Y(
        oc8051_sfr1_oc8051_psw1_n15) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u11 ( .A0(psw_set[0]), .A1(
        oc8051_sfr1_oc8051_psw1_n14), .B0(oc8051_sfr1_oc8051_psw1_n15), .Y(
        oc8051_sfr1_oc8051_psw1_n13) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u10 ( .A(
        oc8051_sfr1_oc8051_psw1_n12), .B(oc8051_sfr1_oc8051_psw1_n1), .S0(
        oc8051_sfr1_oc8051_psw1_n13), .Y(oc8051_sfr1_oc8051_psw1_n48) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u9 ( .A0(
        oc8051_sfr1_oc8051_psw1_n6), .A1(descy), .B0(wr_dat[7]), .B1(
        oc8051_sfr1_oc8051_psw1_n7), .C0(oc8051_sfr1_oc8051_psw1_n11), .Y(
        oc8051_sfr1_oc8051_psw1_n2) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u8 ( .A(cy), .Y(
        oc8051_sfr1_oc8051_psw1_n3) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u7 ( .A(oc8051_sfr1_oc8051_psw1_n8), 
        .B(oc8051_sfr1_oc8051_psw1_n9), .C(oc8051_sfr1_oc8051_psw1_n10), .Y(
        oc8051_sfr1_oc8051_psw1_n5) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u6 ( .A(oc8051_sfr1_oc8051_psw1_n5), 
        .B(oc8051_sfr1_oc8051_psw1_n6), .C(oc8051_sfr1_oc8051_psw1_n7), .Y(
        oc8051_sfr1_oc8051_psw1_n4) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u5 ( .A(oc8051_sfr1_oc8051_psw1_n2), .B(oc8051_sfr1_oc8051_psw1_n3), .S0(oc8051_sfr1_oc8051_psw1_n4), .Y(
        oc8051_sfr1_oc8051_psw1_n49) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u4 ( .A(oc8051_sfr1_oc8051_psw1_n1), 
        .Y(srcac) );
  MXT2_X1M_A12TS oc8051_sfr1_oc8051_psw1_u3 ( .A(wr_dat[3]), .B(
        oc8051_sfr1_psw_3_), .S0(oc8051_sfr1_oc8051_psw1_n16), .Y(bank_sel[0])
         );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_6_ ( .D(
        oc8051_sfr1_oc8051_psw1_n48), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_psw1_n1) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_7_ ( .D(
        oc8051_sfr1_oc8051_psw1_n49), .CK(wb_clk_i), .R(wb_rst_i), .Q(cy) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_3_ ( .D(
        oc8051_sfr1_oc8051_psw1_n45), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_4_ ( .D(
        oc8051_sfr1_oc8051_psw1_n46), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_2_ ( .D(
        oc8051_sfr1_oc8051_psw1_n44), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_1_ ( .D(
        oc8051_sfr1_oc8051_psw1_n43), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_5_ ( .D(
        oc8051_sfr1_oc8051_psw1_n47), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_5_) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u171 ( .AN(oc8051_sfr1_wr_bit_r), .B(n_5_net_), .Y(oc8051_sfr1_oc8051_ports1_n48) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u170 ( .A(
        oc8051_sfr1_oc8051_ports1_n48), .Y(oc8051_sfr1_oc8051_ports1_n45) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u169 ( .A(wr_addr[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n81) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u168 ( .A(
        oc8051_sfr1_oc8051_ports1_n45), .B(oc8051_sfr1_oc8051_ports1_n81), .C(
        wr_addr[4]), .Y(oc8051_sfr1_oc8051_ports1_n82) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u167 ( .A(n_5_net_), .B(
        oc8051_sfr1_oc8051_ports1_n81), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u166 ( .A(
        oc8051_sfr1_oc8051_ports1_n85), .Y(oc8051_sfr1_oc8051_ports1_n88) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u165 ( .A(wr_addr[1]), .B(
        wr_addr[2]), .C(wr_addr[0]), .Y(oc8051_sfr1_oc8051_ports1_n43) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u164 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n43), .Y(
        oc8051_sfr1_oc8051_ports1_n103) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u163 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(descy), .Y(oc8051_sfr1_oc8051_ports1_n105) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u162 ( .A(
        oc8051_sfr1_oc8051_ports1_n105), .Y(oc8051_sfr1_oc8051_ports1_n86) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u161 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_ports1_n105), .Y(oc8051_sfr1_oc8051_ports1_n87)
         );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u160 ( .A0(wr_dat[0]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n40) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u159 ( .A(
        oc8051_sfr1_oc8051_ports1_n43), .Y(oc8051_sfr1_oc8051_ports1_n42) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u158 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n42), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n104) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u157 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n103), 
        .B0(oc8051_sfr1_oc8051_ports1_n40), .C0(oc8051_sfr1_oc8051_ports1_n104), .Y(oc8051_sfr1_oc8051_ports1_n132) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u156 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n91) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u155 ( .A(wr_addr[1]), .B(
        wr_addr[2]), .C(oc8051_sfr1_oc8051_ports1_n91), .Y(
        oc8051_sfr1_oc8051_ports1_n38) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u154 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n38), .Y(
        oc8051_sfr1_oc8051_ports1_n101) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u153 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n35) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u152 ( .A(
        oc8051_sfr1_oc8051_ports1_n38), .Y(oc8051_sfr1_oc8051_ports1_n37) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u151 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n37), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n102) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u150 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n101), 
        .B0(oc8051_sfr1_oc8051_ports1_n35), .C0(oc8051_sfr1_oc8051_ports1_n102), .Y(oc8051_sfr1_oc8051_ports1_n133) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u149 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n94) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u148 ( .A(wr_addr[0]), .B(
        wr_addr[2]), .C(oc8051_sfr1_oc8051_ports1_n94), .Y(
        oc8051_sfr1_oc8051_ports1_n33) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u147 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n33), .Y(
        oc8051_sfr1_oc8051_ports1_n99) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u146 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n30) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u145 ( .A(
        oc8051_sfr1_oc8051_ports1_n33), .Y(oc8051_sfr1_oc8051_ports1_n32) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u144 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n32), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n100) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u143 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n99), 
        .B0(oc8051_sfr1_oc8051_ports1_n30), .C0(oc8051_sfr1_oc8051_ports1_n100), .Y(oc8051_sfr1_oc8051_ports1_n134) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u142 ( .A(
        oc8051_sfr1_oc8051_ports1_n91), .B(wr_addr[2]), .C(
        oc8051_sfr1_oc8051_ports1_n94), .Y(oc8051_sfr1_oc8051_ports1_n28) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u141 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n28), .Y(
        oc8051_sfr1_oc8051_ports1_n97) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u140 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n25) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u139 ( .A(
        oc8051_sfr1_oc8051_ports1_n28), .Y(oc8051_sfr1_oc8051_ports1_n27) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u138 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n27), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n98) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u137 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n97), 
        .B0(oc8051_sfr1_oc8051_ports1_n25), .C0(oc8051_sfr1_oc8051_ports1_n98), 
        .Y(oc8051_sfr1_oc8051_ports1_n135) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u136 ( .A(
        oc8051_sfr1_oc8051_ports1_n91), .B(oc8051_sfr1_oc8051_ports1_n94), .C(
        wr_addr[2]), .Y(oc8051_sfr1_oc8051_ports1_n22) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u135 ( .A(
        oc8051_sfr1_oc8051_ports1_n22), .Y(oc8051_sfr1_oc8051_ports1_n23) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u134 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n23), .Y(
        oc8051_sfr1_oc8051_ports1_n95) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u133 ( .A0(wr_dat[4]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n20) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u132 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n22), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n96) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u131 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n95), 
        .B0(oc8051_sfr1_oc8051_ports1_n20), .C0(oc8051_sfr1_oc8051_ports1_n96), 
        .Y(oc8051_sfr1_oc8051_ports1_n136) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u130 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_ports1_n94), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u129 ( .A(
        oc8051_sfr1_oc8051_ports1_n17), .Y(oc8051_sfr1_oc8051_ports1_n18) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u128 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n18), .Y(
        oc8051_sfr1_oc8051_ports1_n92) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u127 ( .A0(wr_dat[5]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n15) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u126 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n17), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n93) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u125 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n92), 
        .B0(oc8051_sfr1_oc8051_ports1_n15), .C0(oc8051_sfr1_oc8051_ports1_n93), 
        .Y(oc8051_sfr1_oc8051_ports1_n137) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u124 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_ports1_n91), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n12) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u123 ( .A(
        oc8051_sfr1_oc8051_ports1_n12), .Y(oc8051_sfr1_oc8051_ports1_n13) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u122 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n13), .Y(
        oc8051_sfr1_oc8051_ports1_n89) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u121 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n10) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u120 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n12), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n90) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u119 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n89), 
        .B0(oc8051_sfr1_oc8051_ports1_n10), .C0(oc8051_sfr1_oc8051_ports1_n90), 
        .Y(oc8051_sfr1_oc8051_ports1_n138) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u118 ( .A(wr_addr[1]), .B(
        wr_addr[0]), .C(wr_addr[2]), .Y(oc8051_sfr1_oc8051_ports1_n5) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u117 ( .A(
        oc8051_sfr1_oc8051_ports1_n5), .Y(oc8051_sfr1_oc8051_ports1_n8) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u116 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n8), .Y(
        oc8051_sfr1_oc8051_ports1_n83) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u115 ( .A0(wr_dat[7]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n3) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u114 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n5), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n84) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u113 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n83), 
        .B0(oc8051_sfr1_oc8051_ports1_n3), .C0(oc8051_sfr1_oc8051_ports1_n84), 
        .Y(oc8051_sfr1_oc8051_ports1_n139) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u112 ( .A(p0_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n79) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u111 ( .A(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n44) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u110 ( .A(
        oc8051_sfr1_oc8051_ports1_n44), .B(oc8051_sfr1_oc8051_ports1_n81), .C(
        n_5_net_), .Y(oc8051_sfr1_oc8051_ports1_n66) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u109 ( .A0(
        oc8051_sfr1_oc8051_ports1_n42), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n80)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u108 ( .A(
        oc8051_sfr1_oc8051_ports1_n79), .B(oc8051_sfr1_oc8051_ports1_n40), 
        .S0(oc8051_sfr1_oc8051_ports1_n80), .Y(oc8051_sfr1_oc8051_ports1_n140)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u107 ( .A(p0_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n77) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u106 ( .A0(
        oc8051_sfr1_oc8051_ports1_n37), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n78)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u105 ( .A(
        oc8051_sfr1_oc8051_ports1_n77), .B(oc8051_sfr1_oc8051_ports1_n35), 
        .S0(oc8051_sfr1_oc8051_ports1_n78), .Y(oc8051_sfr1_oc8051_ports1_n141)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u104 ( .A(p0_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n75) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u103 ( .A0(
        oc8051_sfr1_oc8051_ports1_n32), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n76)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u102 ( .A(
        oc8051_sfr1_oc8051_ports1_n75), .B(oc8051_sfr1_oc8051_ports1_n30), 
        .S0(oc8051_sfr1_oc8051_ports1_n76), .Y(oc8051_sfr1_oc8051_ports1_n142)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u101 ( .A(p0_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n73) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u100 ( .A0(
        oc8051_sfr1_oc8051_ports1_n27), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n74)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u99 ( .A(
        oc8051_sfr1_oc8051_ports1_n73), .B(oc8051_sfr1_oc8051_ports1_n25), 
        .S0(oc8051_sfr1_oc8051_ports1_n74), .Y(oc8051_sfr1_oc8051_ports1_n143)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u98 ( .A(p0_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n71) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u97 ( .A0(
        oc8051_sfr1_oc8051_ports1_n22), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n72)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u96 ( .A(
        oc8051_sfr1_oc8051_ports1_n71), .B(oc8051_sfr1_oc8051_ports1_n20), 
        .S0(oc8051_sfr1_oc8051_ports1_n72), .Y(oc8051_sfr1_oc8051_ports1_n144)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u95 ( .A(p0_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n69) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u94 ( .A0(
        oc8051_sfr1_oc8051_ports1_n17), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n70)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u93 ( .A(
        oc8051_sfr1_oc8051_ports1_n69), .B(oc8051_sfr1_oc8051_ports1_n15), 
        .S0(oc8051_sfr1_oc8051_ports1_n70), .Y(oc8051_sfr1_oc8051_ports1_n145)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u92 ( .A(p0_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n67) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u91 ( .A0(
        oc8051_sfr1_oc8051_ports1_n12), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n68)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u90 ( .A(
        oc8051_sfr1_oc8051_ports1_n67), .B(oc8051_sfr1_oc8051_ports1_n10), 
        .S0(oc8051_sfr1_oc8051_ports1_n68), .Y(oc8051_sfr1_oc8051_ports1_n146)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u89 ( .A(p0_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n64) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u88 ( .A0(
        oc8051_sfr1_oc8051_ports1_n5), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n65)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u87 ( .A(
        oc8051_sfr1_oc8051_ports1_n64), .B(oc8051_sfr1_oc8051_ports1_n3), .S0(
        oc8051_sfr1_oc8051_ports1_n65), .Y(oc8051_sfr1_oc8051_ports1_n147) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u86 ( .A(p3_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n62) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u85 ( .A(wr_addr[5]), .B(
        n_5_net_), .C(wr_addr[4]), .Y(oc8051_sfr1_oc8051_ports1_n49) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u84 ( .A0(
        oc8051_sfr1_oc8051_ports1_n42), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n63)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u83 ( .A(
        oc8051_sfr1_oc8051_ports1_n62), .B(oc8051_sfr1_oc8051_ports1_n40), 
        .S0(oc8051_sfr1_oc8051_ports1_n63), .Y(oc8051_sfr1_oc8051_ports1_n148)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u82 ( .A(p3_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n60) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u81 ( .A0(
        oc8051_sfr1_oc8051_ports1_n37), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n61)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u80 ( .A(
        oc8051_sfr1_oc8051_ports1_n60), .B(oc8051_sfr1_oc8051_ports1_n35), 
        .S0(oc8051_sfr1_oc8051_ports1_n61), .Y(oc8051_sfr1_oc8051_ports1_n149)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u79 ( .A(p3_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n58) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u78 ( .A0(
        oc8051_sfr1_oc8051_ports1_n32), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n59)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u77 ( .A(
        oc8051_sfr1_oc8051_ports1_n58), .B(oc8051_sfr1_oc8051_ports1_n30), 
        .S0(oc8051_sfr1_oc8051_ports1_n59), .Y(oc8051_sfr1_oc8051_ports1_n150)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u76 ( .A(p3_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n56) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u75 ( .A0(
        oc8051_sfr1_oc8051_ports1_n27), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n57)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u74 ( .A(
        oc8051_sfr1_oc8051_ports1_n56), .B(oc8051_sfr1_oc8051_ports1_n25), 
        .S0(oc8051_sfr1_oc8051_ports1_n57), .Y(oc8051_sfr1_oc8051_ports1_n151)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u73 ( .A(p3_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n54) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u72 ( .A0(
        oc8051_sfr1_oc8051_ports1_n22), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n55)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u71 ( .A(
        oc8051_sfr1_oc8051_ports1_n54), .B(oc8051_sfr1_oc8051_ports1_n20), 
        .S0(oc8051_sfr1_oc8051_ports1_n55), .Y(oc8051_sfr1_oc8051_ports1_n152)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u70 ( .A(p3_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n52) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u69 ( .A0(
        oc8051_sfr1_oc8051_ports1_n17), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n53)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u68 ( .A(
        oc8051_sfr1_oc8051_ports1_n52), .B(oc8051_sfr1_oc8051_ports1_n15), 
        .S0(oc8051_sfr1_oc8051_ports1_n53), .Y(oc8051_sfr1_oc8051_ports1_n153)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u67 ( .A(p3_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n50) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u66 ( .A0(
        oc8051_sfr1_oc8051_ports1_n12), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n51)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u65 ( .A(
        oc8051_sfr1_oc8051_ports1_n50), .B(oc8051_sfr1_oc8051_ports1_n10), 
        .S0(oc8051_sfr1_oc8051_ports1_n51), .Y(oc8051_sfr1_oc8051_ports1_n154)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u64 ( .A(p3_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n46) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u63 ( .A0(
        oc8051_sfr1_oc8051_ports1_n5), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n47)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u62 ( .A(
        oc8051_sfr1_oc8051_ports1_n46), .B(oc8051_sfr1_oc8051_ports1_n3), .S0(
        oc8051_sfr1_oc8051_ports1_n47), .Y(oc8051_sfr1_oc8051_ports1_n155) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u61 ( .A(wr_addr[5]), .B(
        oc8051_sfr1_oc8051_ports1_n44), .C(oc8051_sfr1_oc8051_ports1_n45), .Y(
        oc8051_sfr1_oc8051_ports1_n1) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u60 ( .A(n_5_net_), .B(
        oc8051_sfr1_oc8051_ports1_n44), .C(wr_addr[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n6) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u59 ( .A(
        oc8051_sfr1_oc8051_ports1_n6), .Y(oc8051_sfr1_oc8051_ports1_n7) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u58 ( .A(
        oc8051_sfr1_oc8051_ports1_n43), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n39) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u57 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n42), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n41) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u56 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n39), 
        .B0(oc8051_sfr1_oc8051_ports1_n40), .C0(oc8051_sfr1_oc8051_ports1_n41), 
        .Y(oc8051_sfr1_oc8051_ports1_n156) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u55 ( .A(
        oc8051_sfr1_oc8051_ports1_n38), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n34) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u54 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n37), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n36) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u53 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n34), 
        .B0(oc8051_sfr1_oc8051_ports1_n35), .C0(oc8051_sfr1_oc8051_ports1_n36), 
        .Y(oc8051_sfr1_oc8051_ports1_n157) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u52 ( .A(
        oc8051_sfr1_oc8051_ports1_n33), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n29) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u51 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n32), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n31) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u50 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n29), 
        .B0(oc8051_sfr1_oc8051_ports1_n30), .C0(oc8051_sfr1_oc8051_ports1_n31), 
        .Y(oc8051_sfr1_oc8051_ports1_n158) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u49 ( .A(
        oc8051_sfr1_oc8051_ports1_n28), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n24) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u48 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n27), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n26) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u47 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n24), 
        .B0(oc8051_sfr1_oc8051_ports1_n25), .C0(oc8051_sfr1_oc8051_ports1_n26), 
        .Y(oc8051_sfr1_oc8051_ports1_n159) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u46 ( .A(
        oc8051_sfr1_oc8051_ports1_n23), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n19) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u45 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n22), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n21) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u44 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n19), 
        .B0(oc8051_sfr1_oc8051_ports1_n20), .C0(oc8051_sfr1_oc8051_ports1_n21), 
        .Y(oc8051_sfr1_oc8051_ports1_n160) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u43 ( .A(
        oc8051_sfr1_oc8051_ports1_n18), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n14) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u42 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n17), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n16) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u41 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n14), 
        .B0(oc8051_sfr1_oc8051_ports1_n15), .C0(oc8051_sfr1_oc8051_ports1_n16), 
        .Y(oc8051_sfr1_oc8051_ports1_n161) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u40 ( .A(
        oc8051_sfr1_oc8051_ports1_n13), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n9) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u39 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n12), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n11) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u38 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n9), .B0(
        oc8051_sfr1_oc8051_ports1_n10), .C0(oc8051_sfr1_oc8051_ports1_n11), 
        .Y(oc8051_sfr1_oc8051_ports1_n162) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u37 ( .A(
        oc8051_sfr1_oc8051_ports1_n7), .B(oc8051_sfr1_oc8051_ports1_n8), .Y(
        oc8051_sfr1_oc8051_ports1_n2) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u36 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n5), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n4) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u35 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n2), .B0(
        oc8051_sfr1_oc8051_ports1_n3), .C0(oc8051_sfr1_oc8051_ports1_n4), .Y(
        oc8051_sfr1_oc8051_ports1_n163) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u34 ( .A(p0_i[0]), .B(p0_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u33 ( .A(p0_i[1]), .B(p0_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u32 ( .A(p0_i[2]), .B(p0_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u31 ( .A(p0_i[3]), .B(p0_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u30 ( .A(p0_i[4]), .B(p0_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u29 ( .A(p0_i[5]), .B(p0_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u28 ( .A(p0_i[6]), .B(p0_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u27 ( .A(p0_i[7]), .B(p0_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_7_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u26 ( .A(p1_i[0]), .B(p1_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u25 ( .A(p1_i[1]), .B(p1_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u24 ( .A(p1_i[2]), .B(p1_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u23 ( .A(p1_i[3]), .B(p1_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u22 ( .A(p1_i[4]), .B(p1_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u21 ( .A(p1_i[5]), .B(p1_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u20 ( .A(p1_i[6]), .B(p1_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u19 ( .A(p1_i[7]), .B(p1_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_7_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u18 ( .A(p2_i[0]), .B(p2_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u17 ( .A(p2_i[1]), .B(p2_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u16 ( .A(p2_i[2]), .B(p2_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u15 ( .A(p2_i[3]), .B(p2_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u14 ( .A(p2_i[4]), .B(p2_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u13 ( .A(p2_i[5]), .B(p2_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u12 ( .A(p2_i[6]), .B(p2_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u11 ( .A(p2_i[7]), .B(p2_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_7_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u10 ( .A(p3_i[0]), .B(p3_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u9 ( .A(p3_i[1]), .B(p3_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u8 ( .A(p3_i[2]), .B(p3_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u7 ( .A(p3_i[3]), .B(p3_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u6 ( .A(p3_i[4]), .B(p3_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u5 ( .A(p3_i[5]), .B(p3_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u4 ( .A(p3_i[6]), .B(p3_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u3 ( .A(p3_i[7]), .B(p3_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_7_) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_ports1_u2 ( .A(wb_rst_i), .Y(
        oc8051_sfr1_oc8051_ports1_n106) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n140), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n141), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n142), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n143), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n144), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n145), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n146), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n147), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[7]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n148), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n149), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n150), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n151), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n152), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n153), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n154), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n155), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[7]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n132), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n133), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n134), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n135), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n136), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n137), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n138), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n139), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[7]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n156), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n157), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n158), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n159), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n160), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n161), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n162), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n163), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[7]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u238 ( .A(oc8051_sfr1_pcon[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n161) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u237 ( .A(oc8051_sfr1_scon_6_), .Y(
        oc8051_sfr1_oc8051_uatr1_n30) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u236 ( .A(
        oc8051_sfr1_oc8051_uatr1_n205), .Y(oc8051_sfr1_oc8051_uatr1_n165) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u235 ( .A(oc8051_sfr1_tf1), .Y(
        oc8051_sfr1_oc8051_uatr1_n166) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u234 ( .A(
        oc8051_sfr1_oc8051_uatr1_n165), .B(oc8051_sfr1_oc8051_uatr1_n166), .Y(
        oc8051_sfr1_oc8051_uatr1_n163) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u233 ( .A(
        oc8051_sfr1_oc8051_uatr1_n163), .B(oc8051_sfr1_brate2), .S0(
        oc8051_sfr1_tclk), .Y(oc8051_sfr1_oc8051_uatr1_n164) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u232 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n30), .A1(oc8051_sfr1_scon_7_), .B0(
        oc8051_sfr1_oc8051_uatr1_n164), .Y(oc8051_sfr1_oc8051_uatr1_n2) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u231 ( .A1N(
        oc8051_sfr1_oc8051_uatr1_smod_clk_tr), .A0(
        oc8051_sfr1_oc8051_uatr1_n161), .B0(oc8051_sfr1_oc8051_uatr1_n2), .Y(
        oc8051_sfr1_oc8051_uatr1_n174) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u230 ( .A(
        oc8051_sfr1_oc8051_uatr1_n163), .B(oc8051_sfr1_brate2), .S0(
        oc8051_sfr1_rclk), .Y(oc8051_sfr1_oc8051_uatr1_n162) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u229 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n30), .A1(oc8051_sfr1_scon_7_), .B0(
        oc8051_sfr1_oc8051_uatr1_n162), .Y(oc8051_sfr1_oc8051_uatr1_n91) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u228 ( .A1N(
        oc8051_sfr1_oc8051_uatr1_smod_clk_re), .A0(
        oc8051_sfr1_oc8051_uatr1_n161), .B0(oc8051_sfr1_oc8051_uatr1_n91), .Y(
        oc8051_sfr1_oc8051_uatr1_n269) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u227 ( .A(oc8051_sfr1_scon_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n117) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u226 ( .A(
        oc8051_sfr1_oc8051_uatr1_n180), .B(oc8051_sfr1_oc8051_uatr1_n117), .Y(
        oc8051_sfr1_uart_int) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u225 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_), .B(oc8051_sfr1_sbuf[7]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n181) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u224 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_), .B(oc8051_sfr1_sbuf[6]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n182) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u223 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_), .B(oc8051_sfr1_sbuf[5]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n183) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u222 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_), .B(oc8051_sfr1_sbuf[4]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n184) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u221 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_), .B(oc8051_sfr1_sbuf[3]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n185) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u220 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_), .B(oc8051_sfr1_sbuf[2]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n186) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u219 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_), .B(oc8051_sfr1_sbuf[1]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n187) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u218 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_), .B(oc8051_sfr1_sbuf[0]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n188) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u217 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_uatr1_n22) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u216 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_uatr1_n21) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u215 ( .A(
        oc8051_sfr1_oc8051_uatr1_n22), .B(oc8051_sfr1_oc8051_uatr1_n21), .Y(
        oc8051_sfr1_oc8051_uatr1_n16) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u214 ( .A(wr_addr[6]), .B(
        wr_addr[5]), .Y(oc8051_sfr1_oc8051_uatr1_n160) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u213 ( .A(wr_addr[7]), .B(n_5_net_), .C(oc8051_sfr1_oc8051_uatr1_n160), .Y(oc8051_sfr1_oc8051_uatr1_n129) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u212 ( .A(wr_addr[3]), .B(
        oc8051_sfr1_wr_bit_r), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_uatr1_n159) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u211 ( .A(
        oc8051_sfr1_oc8051_uatr1_n16), .B(oc8051_sfr1_oc8051_uatr1_n129), .C(
        wr_addr[2]), .D(oc8051_sfr1_oc8051_uatr1_n159), .Y(
        oc8051_sfr1_oc8051_uatr1_n158) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u210 ( .A(oc8051_sfr1_pcon[0]), 
        .B(wr_dat[0]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n190) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u209 ( .A(oc8051_sfr1_pcon[1]), 
        .B(wr_dat[1]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n191) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u208 ( .A(oc8051_sfr1_pcon[2]), 
        .B(wr_dat[2]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n192) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u207 ( .A(oc8051_sfr1_pcon[3]), 
        .B(wr_dat[3]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n193) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u206 ( .A(oc8051_sfr1_pcon[4]), 
        .B(wr_dat[4]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n194) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u205 ( .A(oc8051_sfr1_pcon[5]), 
        .B(wr_dat[5]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n195) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u204 ( .A(oc8051_sfr1_pcon[6]), 
        .B(wr_dat[6]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n196) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u203 ( .A(oc8051_sfr1_pcon[7]), 
        .B(wr_dat[7]), .S0(oc8051_sfr1_oc8051_uatr1_n158), .Y(
        oc8051_sfr1_oc8051_uatr1_n197) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u202 ( .A(oc8051_sfr1_scon_7_), .Y(
        oc8051_sfr1_oc8051_uatr1_n34) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u201 ( .A(
        oc8051_sfr1_oc8051_uatr1_n30), .B(oc8051_sfr1_oc8051_uatr1_n34), .Y(
        oc8051_sfr1_oc8051_uatr1_n88) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u200 ( .A(
        oc8051_sfr1_oc8051_uatr1_receive), .B(oc8051_sfr1_oc8051_uatr1_n88), 
        .C(oc8051_sfr1_oc8051_uatr1_shift_re), .Y(
        oc8051_sfr1_oc8051_uatr1_n147) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u199 ( .A(
        oc8051_sfr1_oc8051_uatr1_n147), .Y(oc8051_sfr1_oc8051_uatr1_n140) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u198 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_done), .B(oc8051_sfr1_oc8051_uatr1_n140), 
        .Y(oc8051_sfr1_oc8051_uatr1_n95) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u197 ( .A(
        oc8051_sfr1_oc8051_uatr1_n95), .Y(oc8051_sfr1_oc8051_uatr1_n101) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u196 ( .A(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .B(
        oc8051_sfr1_oc8051_uatr1_n101), .C(
        oc8051_sfr1_oc8051_uatr1_re_count_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n108) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u195 ( .A(
        oc8051_sfr1_oc8051_uatr1_n88), .Y(oc8051_sfr1_oc8051_uatr1_n77) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u194 ( .A(oc8051_sfr1_pres_ow), 
        .B(oc8051_sfr1_oc8051_uatr1_n77), .C(oc8051_sfr1_oc8051_uatr1_receive), 
        .Y(oc8051_sfr1_oc8051_uatr1_n103) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u193 ( .A(
        oc8051_sfr1_oc8051_uatr1_n103), .Y(oc8051_sfr1_oc8051_uatr1_n106) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u192 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_done), .Y(oc8051_sfr1_oc8051_uatr1_n127)
         );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u191 ( .A(
        oc8051_sfr1_oc8051_uatr1_n106), .B(oc8051_sfr1_oc8051_uatr1_n140), .C(
        oc8051_sfr1_oc8051_uatr1_n127), .Y(oc8051_sfr1_oc8051_uatr1_n137) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u190 ( .A(
        oc8051_sfr1_oc8051_uatr1_n137), .B(oc8051_sfr1_oc8051_uatr1_shift_re), 
        .C(oc8051_sfr1_scon_4_), .D(oc8051_sfr1_oc8051_uatr1_n88), .Y(
        oc8051_sfr1_oc8051_uatr1_n148) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u189 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n137), .B(oc8051_sfr1_oc8051_uatr1_n88), .Y(
        oc8051_sfr1_oc8051_uatr1_n135) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u188 ( .A(oc8051_sfr1_scon_0_), 
        .B(oc8051_sfr1_oc8051_uatr1_receive), .Y(oc8051_sfr1_oc8051_uatr1_n133) );
  AOI32_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u187 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n135), .A1(oc8051_sfr1_scon_4_), .A2(
        oc8051_sfr1_oc8051_uatr1_n133), .B0(oc8051_sfr1_oc8051_uatr1_n106), 
        .B1(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n157) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u186 ( .A(
        oc8051_sfr1_oc8051_uatr1_n108), .B(oc8051_sfr1_oc8051_uatr1_n148), .C(
        oc8051_sfr1_oc8051_uatr1_n157), .Y(oc8051_sfr1_oc8051_uatr1_n100) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u185 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_), .Y(
        oc8051_sfr1_oc8051_uatr1_n156) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u184 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_), .Y(
        oc8051_sfr1_oc8051_uatr1_n98) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u183 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n101), .A1(oc8051_sfr1_oc8051_uatr1_n106), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .Y(oc8051_sfr1_oc8051_uatr1_n104)
         );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u182 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n100), .A1(oc8051_sfr1_oc8051_uatr1_n156), 
        .B0(oc8051_sfr1_oc8051_uatr1_n98), .B1(oc8051_sfr1_oc8051_uatr1_n104), 
        .Y(oc8051_sfr1_oc8051_uatr1_n206) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u181 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_), .Y(
        oc8051_sfr1_oc8051_uatr1_n155) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u180 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_), .Y(
        oc8051_sfr1_oc8051_uatr1_n154) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u179 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n155), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .B1(oc8051_sfr1_oc8051_uatr1_n154), 
        .C0(oc8051_sfr1_oc8051_uatr1_n148), .Y(oc8051_sfr1_oc8051_uatr1_n207)
         );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u178 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n100), .A1(oc8051_sfr1_oc8051_uatr1_n155), 
        .B0(oc8051_sfr1_oc8051_uatr1_n104), .B1(oc8051_sfr1_oc8051_uatr1_n156), 
        .Y(oc8051_sfr1_oc8051_uatr1_n208) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u177 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_), .Y(
        oc8051_sfr1_oc8051_uatr1_n153) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u176 ( .A(
        oc8051_sfr1_oc8051_uatr1_n148), .Y(oc8051_sfr1_oc8051_uatr1_n134) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u175 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n135), .A1(oc8051_sfr1_oc8051_uatr1_n134), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .Y(oc8051_sfr1_oc8051_uatr1_n105)
         );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u174 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n154), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .B1(oc8051_sfr1_oc8051_uatr1_n153), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n209)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u173 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_), .Y(
        oc8051_sfr1_oc8051_uatr1_n152) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u172 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n153), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .B1(oc8051_sfr1_oc8051_uatr1_n152), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n210)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u171 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_), .Y(
        oc8051_sfr1_oc8051_uatr1_n151) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u170 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n152), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .B1(oc8051_sfr1_oc8051_uatr1_n151), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n211)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u169 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_), .Y(
        oc8051_sfr1_oc8051_uatr1_n150) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u168 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n151), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .B1(oc8051_sfr1_oc8051_uatr1_n150), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n212)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u167 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n149) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u166 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n150), 
        .B0(oc8051_sfr1_oc8051_uatr1_n100), .B1(oc8051_sfr1_oc8051_uatr1_n149), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n213)
         );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u165 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n149), 
        .B0(oc8051_sfr1_oc8051_uatr1_n202), .B1(oc8051_sfr1_oc8051_uatr1_n100), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n214)
         );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u164 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n202), .A1(oc8051_sfr1_oc8051_uatr1_n104), 
        .B0(oc8051_sfr1_oc8051_uatr1_n203), .B1(oc8051_sfr1_oc8051_uatr1_n100), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n215)
         );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u163 ( .A(
        oc8051_sfr1_oc8051_uatr1_n148), .B(oc8051_sfr1_oc8051_uatr1_n95), .Y(
        oc8051_sfr1_oc8051_uatr1_n139) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u162 ( .A(
        oc8051_sfr1_oc8051_uatr1_n140), .B(oc8051_sfr1_oc8051_uatr1_n139), .C(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n141) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u161 ( .A(
        oc8051_sfr1_oc8051_uatr1_n141), .B(
        oc8051_sfr1_oc8051_uatr1_re_count_1_), .C(
        oc8051_sfr1_oc8051_uatr1_re_count_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n145) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u160 ( .A0(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .A1(
        oc8051_sfr1_oc8051_uatr1_n147), .B0(oc8051_sfr1_oc8051_uatr1_n139), 
        .Y(oc8051_sfr1_oc8051_uatr1_n142) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u159 ( .A1N(
        oc8051_sfr1_oc8051_uatr1_re_count_1_), .A0(
        oc8051_sfr1_oc8051_uatr1_n140), .B0(oc8051_sfr1_oc8051_uatr1_n142), 
        .Y(oc8051_sfr1_oc8051_uatr1_n144) );
  OA21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u158 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n147), .A1(
        oc8051_sfr1_oc8051_uatr1_re_count_2_), .B0(
        oc8051_sfr1_oc8051_uatr1_n144), .Y(oc8051_sfr1_oc8051_uatr1_n146) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u157 ( .A(
        oc8051_sfr1_oc8051_uatr1_n145), .B(oc8051_sfr1_oc8051_uatr1_n146), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n216) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u156 ( .A(
        oc8051_sfr1_oc8051_uatr1_n141), .B(
        oc8051_sfr1_oc8051_uatr1_re_count_1_), .Y(
        oc8051_sfr1_oc8051_uatr1_n143) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u155 ( .A(
        oc8051_sfr1_oc8051_uatr1_n143), .B(oc8051_sfr1_oc8051_uatr1_n144), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n217) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u154 ( .A(
        oc8051_sfr1_oc8051_uatr1_n141), .B(oc8051_sfr1_oc8051_uatr1_n142), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_1_), .Y(
        oc8051_sfr1_oc8051_uatr1_n218) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u153 ( .A(
        oc8051_sfr1_oc8051_uatr1_n140), .B(oc8051_sfr1_oc8051_uatr1_n139), .Y(
        oc8051_sfr1_oc8051_uatr1_n138) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u152 ( .A(
        oc8051_sfr1_oc8051_uatr1_n138), .B(oc8051_sfr1_oc8051_uatr1_n139), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n219) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u151 ( .A(oc8051_sfr1_scon_4_), .Y(
        oc8051_sfr1_oc8051_uatr1_n20) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u150 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n88), .A1(oc8051_sfr1_oc8051_uatr1_n20), .A2(
        oc8051_sfr1_oc8051_uatr1_n137), .B0(oc8051_sfr1_oc8051_uatr1_n134), 
        .Y(oc8051_sfr1_oc8051_uatr1_n136) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u149 ( .A(rxd_i), .B(
        oc8051_sfr1_oc8051_uatr1_rxd_r), .S0(oc8051_sfr1_oc8051_uatr1_n136), 
        .Y(oc8051_sfr1_oc8051_uatr1_n220) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u148 ( .A(rxd_i), .Y(
        oc8051_sfr1_oc8051_uatr1_n93) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u147 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n134), .A1(oc8051_sfr1_oc8051_uatr1_n93), 
        .A2(oc8051_sfr1_oc8051_uatr1_rxd_r), .B0(oc8051_sfr1_oc8051_uatr1_n135), .Y(oc8051_sfr1_oc8051_uatr1_n130) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u146 ( .A(
        oc8051_sfr1_oc8051_uatr1_receive), .Y(oc8051_sfr1_oc8051_uatr1_n131)
         );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u145 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n133), .A1(oc8051_sfr1_scon_4_), .B0(
        oc8051_sfr1_oc8051_uatr1_n127), .C0(oc8051_sfr1_oc8051_uatr1_n134), 
        .Y(oc8051_sfr1_oc8051_uatr1_n132) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u144 ( .A(
        oc8051_sfr1_oc8051_uatr1_n130), .B(oc8051_sfr1_oc8051_uatr1_n131), 
        .S0(oc8051_sfr1_oc8051_uatr1_n132), .Y(oc8051_sfr1_oc8051_uatr1_n221)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u143 ( .A(wr_addr[3]), .B(
        oc8051_sfr1_oc8051_uatr1_n129), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_uatr1_n128) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u142 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_uatr1_n128), .Y(oc8051_sfr1_oc8051_uatr1_n36) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u141 ( .A(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_uatr1_n35) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u140 ( .AN(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_uatr1_n128), .C(oc8051_sfr1_oc8051_uatr1_n22), 
        .D(oc8051_sfr1_oc8051_uatr1_n35), .Y(oc8051_sfr1_oc8051_uatr1_n89) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u139 ( .A(
        oc8051_sfr1_oc8051_uatr1_n89), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_uatr1_n14) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u138 ( .A(
        oc8051_sfr1_oc8051_uatr1_n14), .Y(oc8051_sfr1_oc8051_uatr1_n115) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u137 ( .A(
        oc8051_sfr1_oc8051_uatr1_n198), .B(oc8051_sfr1_oc8051_uatr1_n36), .C(
        oc8051_sfr1_oc8051_uatr1_n115), .D(oc8051_sfr1_oc8051_uatr1_n127), .Y(
        oc8051_sfr1_oc8051_uatr1_n119) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u136 ( .A(
        oc8051_sfr1_oc8051_uatr1_n36), .Y(oc8051_sfr1_oc8051_uatr1_n126) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u135 ( .A(descy), .B(
        oc8051_sfr1_oc8051_uatr1_n126), .Y(oc8051_sfr1_oc8051_uatr1_n11) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u134 ( .A(
        oc8051_sfr1_oc8051_uatr1_n11), .Y(oc8051_sfr1_oc8051_uatr1_n113) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u133 ( .A0(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_), .A1(
        oc8051_sfr1_oc8051_uatr1_n119), .B0(oc8051_sfr1_oc8051_uatr1_n14), 
        .B1(wr_dat[2]), .C0(oc8051_sfr1_oc8051_uatr1_n113), .Y(
        oc8051_sfr1_oc8051_uatr1_n122) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u132 ( .A(oc8051_sfr1_scon_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n123) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u131 ( .A(
        oc8051_sfr1_oc8051_uatr1_n126), .B(oc8051_sfr1_oc8051_uatr1_n35), .Y(
        oc8051_sfr1_oc8051_uatr1_n15) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u130 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n15), .A1(wr_addr[0]), .A2(
        oc8051_sfr1_oc8051_uatr1_n22), .B0(oc8051_sfr1_oc8051_uatr1_n115), .Y(
        oc8051_sfr1_oc8051_uatr1_n125) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u129 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n119), .A1(oc8051_sfr1_oc8051_uatr1_n88), 
        .B0(oc8051_sfr1_oc8051_uatr1_n125), .Y(oc8051_sfr1_oc8051_uatr1_n124)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u128 ( .A(
        oc8051_sfr1_oc8051_uatr1_n122), .B(oc8051_sfr1_oc8051_uatr1_n123), 
        .S0(oc8051_sfr1_oc8051_uatr1_n124), .Y(oc8051_sfr1_oc8051_uatr1_n222)
         );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u127 ( .A0(wr_dat[0]), .A1(
        oc8051_sfr1_oc8051_uatr1_n14), .B0(oc8051_sfr1_oc8051_uatr1_n113), 
        .C0(oc8051_sfr1_oc8051_uatr1_n119), .Y(oc8051_sfr1_oc8051_uatr1_n116)
         );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u126 ( .A(
        oc8051_sfr1_oc8051_uatr1_n88), .B(oc8051_sfr1_oc8051_uatr1_n98), .C(
        oc8051_sfr1_scon_5_), .Y(oc8051_sfr1_oc8051_uatr1_n120) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u125 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n15), .A1(wr_addr[1]), .A2(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_uatr1_n115), .Y(oc8051_sfr1_oc8051_uatr1_n121) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u124 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n119), .A1(oc8051_sfr1_oc8051_uatr1_n120), 
        .B0(oc8051_sfr1_oc8051_uatr1_n121), .Y(oc8051_sfr1_oc8051_uatr1_n118)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u123 ( .A(
        oc8051_sfr1_oc8051_uatr1_n116), .B(oc8051_sfr1_oc8051_uatr1_n117), 
        .S0(oc8051_sfr1_oc8051_uatr1_n118), .Y(oc8051_sfr1_oc8051_uatr1_n223)
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u122 ( .A(wr_dat[1]), .B(
        oc8051_sfr1_oc8051_uatr1_n36), .S0(oc8051_sfr1_oc8051_uatr1_n115), .Y(
        oc8051_sfr1_oc8051_uatr1_n114) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u121 ( .A(
        oc8051_sfr1_oc8051_uatr1_n113), .B(oc8051_sfr1_oc8051_uatr1_n114), .Y(
        oc8051_sfr1_oc8051_uatr1_n109) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u120 ( .A(
        oc8051_sfr1_oc8051_uatr1_n198), .Y(oc8051_sfr1_oc8051_uatr1_n111) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u119 ( .A(
        oc8051_sfr1_oc8051_uatr1_n15), .B(wr_addr[1]), .C(
        oc8051_sfr1_oc8051_uatr1_n21), .Y(oc8051_sfr1_oc8051_uatr1_n112) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u118 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n36), .A1(oc8051_sfr1_oc8051_uatr1_n111), 
        .B0(oc8051_sfr1_oc8051_uatr1_n14), .C0(oc8051_sfr1_oc8051_uatr1_n112), 
        .Y(oc8051_sfr1_oc8051_uatr1_n110) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u117 ( .A(
        oc8051_sfr1_oc8051_uatr1_n109), .B(oc8051_sfr1_oc8051_uatr1_n180), 
        .S0(oc8051_sfr1_oc8051_uatr1_n110), .Y(oc8051_sfr1_oc8051_uatr1_n224)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u116 ( .A(
        oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n107) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u115 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n106), .A1(oc8051_sfr1_oc8051_uatr1_n107), 
        .B0(oc8051_sfr1_oc8051_uatr1_rx_done), .C0(
        oc8051_sfr1_oc8051_uatr1_n204), .Y(oc8051_sfr1_oc8051_uatr1_n225) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u114 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n203), .A1(oc8051_sfr1_oc8051_uatr1_n104), 
        .B0(oc8051_sfr1_oc8051_uatr1_n204), .B1(oc8051_sfr1_oc8051_uatr1_n100), 
        .C0(oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n226)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u113 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_sam_1_), .Y(oc8051_sfr1_oc8051_uatr1_n96)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u112 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_sam_0_), .Y(oc8051_sfr1_oc8051_uatr1_n92)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u111 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n96), .A1(oc8051_sfr1_oc8051_uatr1_n92), .B0(
        oc8051_sfr1_oc8051_uatr1_n95), .C0(oc8051_sfr1_oc8051_uatr1_n103), .Y(
        oc8051_sfr1_oc8051_uatr1_n102) );
  AOI32_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u110 ( .A0(
        oc8051_sfr1_oc8051_uatr1_rx_sam_0_), .A1(oc8051_sfr1_oc8051_uatr1_n101), .A2(oc8051_sfr1_oc8051_uatr1_rx_sam_1_), .B0(rxd_i), .B1(
        oc8051_sfr1_oc8051_uatr1_n102), .Y(oc8051_sfr1_oc8051_uatr1_n99) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u109 ( .A(
        oc8051_sfr1_oc8051_uatr1_n98), .B(oc8051_sfr1_oc8051_uatr1_n99), .S0(
        oc8051_sfr1_oc8051_uatr1_n100), .Y(oc8051_sfr1_oc8051_uatr1_n227) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u108 ( .A(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .B(oc8051_sfr1_oc8051_uatr1_n95), .Y(oc8051_sfr1_oc8051_uatr1_n97) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u107 ( .A(
        oc8051_sfr1_oc8051_uatr1_n96), .B(oc8051_sfr1_oc8051_uatr1_n93), .S0(
        oc8051_sfr1_oc8051_uatr1_n97), .Y(oc8051_sfr1_oc8051_uatr1_n228) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u106 ( .A(
        oc8051_sfr1_oc8051_uatr1_re_count_3_), .B(oc8051_sfr1_oc8051_uatr1_n95), .Y(oc8051_sfr1_oc8051_uatr1_n94) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u105 ( .A(
        oc8051_sfr1_oc8051_uatr1_n92), .B(oc8051_sfr1_oc8051_uatr1_n93), .S0(
        oc8051_sfr1_oc8051_uatr1_n94), .Y(oc8051_sfr1_oc8051_uatr1_n229) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u104 ( .A(
        oc8051_sfr1_oc8051_uatr1_n91), .B(oc8051_sfr1_pcon[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n90) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u103 ( .A(
        oc8051_sfr1_oc8051_uatr1_smod_clk_re), .B(oc8051_sfr1_oc8051_uatr1_n90), .Y(oc8051_sfr1_oc8051_uatr1_n230) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u102 ( .A(
        oc8051_sfr1_oc8051_uatr1_trans), .Y(oc8051_sfr1_oc8051_uatr1_n39) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u101 ( .A(
        oc8051_sfr1_oc8051_uatr1_n21), .B(oc8051_sfr1_oc8051_uatr1_n89), .Y(
        oc8051_sfr1_oc8051_uatr1_n54) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u100 ( .A(
        oc8051_sfr1_oc8051_uatr1_n39), .B(oc8051_sfr1_oc8051_uatr1_n54), .Y(
        oc8051_sfr1_oc8051_uatr1_n5) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u99 ( .A(
        oc8051_sfr1_oc8051_uatr1_n5), .B(oc8051_sfr1_oc8051_uatr1_n88), .C(
        oc8051_sfr1_oc8051_uatr1_shift_tr), .Y(oc8051_sfr1_oc8051_uatr1_n55)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u98 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_), .Y(oc8051_sfr1_oc8051_uatr1_n60) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u97 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_), .B(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_), .C(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_), .Y(oc8051_sfr1_oc8051_uatr1_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u96 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_7_), .Y(oc8051_sfr1_oc8051_uatr1_n73) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u95 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_), .Y(oc8051_sfr1_oc8051_uatr1_n75) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u94 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_6_), .Y(oc8051_sfr1_oc8051_uatr1_n71) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u93 ( .A(
        oc8051_sfr1_oc8051_uatr1_n73), .B(oc8051_sfr1_oc8051_uatr1_n75), .C(
        oc8051_sfr1_oc8051_uatr1_n71), .Y(oc8051_sfr1_oc8051_uatr1_n87) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u92 ( .A(
        oc8051_sfr1_oc8051_uatr1_n87), .B(oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_), .C(oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_), .Y(oc8051_sfr1_oc8051_uatr1_n86)
         );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u91 ( .A(
        oc8051_sfr1_oc8051_uatr1_n200), .B(oc8051_sfr1_oc8051_uatr1_n199), .C(
        oc8051_sfr1_oc8051_uatr1_n85), .D(oc8051_sfr1_oc8051_uatr1_n86), .Y(
        oc8051_sfr1_oc8051_uatr1_n41) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u90 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n55), .B(oc8051_sfr1_oc8051_uatr1_n60), .C(
        oc8051_sfr1_oc8051_uatr1_n41), .Y(oc8051_sfr1_oc8051_uatr1_n8) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u89 ( .A(
        oc8051_sfr1_oc8051_uatr1_n8), .B(oc8051_sfr1_oc8051_uatr1_n60), .C(
        oc8051_sfr1_oc8051_uatr1_trans), .Y(oc8051_sfr1_oc8051_uatr1_n82) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u88 ( .A(
        oc8051_sfr1_oc8051_uatr1_n54), .Y(oc8051_sfr1_oc8051_uatr1_n37) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u87 ( .A(
        oc8051_sfr1_oc8051_uatr1_n77), .B(oc8051_sfr1_oc8051_uatr1_n5), .C(
        oc8051_sfr1_pres_ow), .Y(oc8051_sfr1_oc8051_uatr1_n7) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u86 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .Y(oc8051_sfr1_oc8051_uatr1_n84) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u85 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_2_), .Y(oc8051_sfr1_oc8051_uatr1_n46) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u84 ( .AN(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .B(oc8051_sfr1_oc8051_uatr1_n84), .C(oc8051_sfr1_oc8051_uatr1_n201), .D(oc8051_sfr1_oc8051_uatr1_n46), .Y(
        oc8051_sfr1_oc8051_uatr1_n42) );
  OR2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u83 ( .A(
        oc8051_sfr1_oc8051_uatr1_n42), .B(oc8051_sfr1_oc8051_uatr1_n55), .Y(
        oc8051_sfr1_oc8051_uatr1_n6) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u82 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n41), .A1(oc8051_sfr1_oc8051_uatr1_n7), .B0(
        oc8051_sfr1_oc8051_uatr1_n6), .Y(oc8051_sfr1_oc8051_uatr1_n81) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u81 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n37), .A1(oc8051_sfr1_oc8051_uatr1_n39), .B0(
        oc8051_sfr1_oc8051_uatr1_n81), .Y(oc8051_sfr1_oc8051_uatr1_n83) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u80 ( .A(
        oc8051_sfr1_oc8051_uatr1_n82), .B(txd_o), .S0(
        oc8051_sfr1_oc8051_uatr1_n83), .Y(oc8051_sfr1_oc8051_uatr1_n231) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u79 ( .A(
        oc8051_sfr1_oc8051_uatr1_n81), .B(oc8051_sfr1_oc8051_uatr1_n54), .Y(
        oc8051_sfr1_oc8051_uatr1_n79) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u78 ( .A(
        oc8051_sfr1_oc8051_uatr1_n79), .Y(oc8051_sfr1_oc8051_uatr1_n38) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u77 ( .B0(
        oc8051_sfr1_oc8051_uatr1_n7), .B1(oc8051_sfr1_oc8051_uatr1_n55), .A0N(
        oc8051_sfr1_oc8051_uatr1_n38), .Y(oc8051_sfr1_oc8051_uatr1_n56) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u76 ( .A(oc8051_sfr1_scon_6_), 
        .B(oc8051_sfr1_scon_3_), .S0(oc8051_sfr1_scon_7_), .Y(
        oc8051_sfr1_oc8051_uatr1_n80) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u75 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n199), .A1(oc8051_sfr1_oc8051_uatr1_n56), 
        .B0(oc8051_sfr1_oc8051_uatr1_n37), .B1(oc8051_sfr1_oc8051_uatr1_n80), 
        .C0(oc8051_sfr1_oc8051_uatr1_n200), .C1(oc8051_sfr1_oc8051_uatr1_n38), 
        .Y(oc8051_sfr1_oc8051_uatr1_n232) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u74 ( .A(
        oc8051_sfr1_oc8051_uatr1_n54), .B(oc8051_sfr1_oc8051_uatr1_n77), .Y(
        oc8051_sfr1_oc8051_uatr1_n58) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u73 ( .A0(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_), .A1(
        oc8051_sfr1_oc8051_uatr1_n79), .B0(oc8051_sfr1_oc8051_uatr1_n54), .B1(
        wr_dat[7]), .Y(oc8051_sfr1_oc8051_uatr1_n78) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u72 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n200), .A1(oc8051_sfr1_oc8051_uatr1_n56), 
        .B0(oc8051_sfr1_oc8051_uatr1_n58), .C0(oc8051_sfr1_oc8051_uatr1_n78), 
        .Y(oc8051_sfr1_oc8051_uatr1_n233) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u71 ( .A(
        oc8051_sfr1_oc8051_uatr1_n37), .B(oc8051_sfr1_oc8051_uatr1_n77), .Y(
        oc8051_sfr1_oc8051_uatr1_n63) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u70 ( .A(
        oc8051_sfr1_oc8051_uatr1_n58), .Y(oc8051_sfr1_oc8051_uatr1_n64) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u69 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n63), .A1(wr_dat[6]), .B0(
        oc8051_sfr1_oc8051_uatr1_n64), .B1(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n76) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u68 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n75), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n73), .C0(
        oc8051_sfr1_oc8051_uatr1_n76), .Y(oc8051_sfr1_oc8051_uatr1_n234) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u67 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n63), .A1(wr_dat[5]), .B0(
        oc8051_sfr1_oc8051_uatr1_n64), .B1(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_uatr1_n74) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u66 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n73), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n71), .C0(
        oc8051_sfr1_oc8051_uatr1_n74), .Y(oc8051_sfr1_oc8051_uatr1_n235) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u65 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_), .Y(oc8051_sfr1_oc8051_uatr1_n69) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u64 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n63), .A1(wr_dat[4]), .B0(
        oc8051_sfr1_oc8051_uatr1_n64), .B1(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_uatr1_n72) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u63 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n71), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n69), .C0(
        oc8051_sfr1_oc8051_uatr1_n72), .Y(oc8051_sfr1_oc8051_uatr1_n236) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u62 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_), .Y(oc8051_sfr1_oc8051_uatr1_n67) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u61 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n63), .A1(wr_dat[3]), .B0(
        oc8051_sfr1_oc8051_uatr1_n64), .B1(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_uatr1_n70) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u60 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n69), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n67), .C0(
        oc8051_sfr1_oc8051_uatr1_n70), .Y(oc8051_sfr1_oc8051_uatr1_n237) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u59 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_), .Y(oc8051_sfr1_oc8051_uatr1_n65) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u58 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_uatr1_n63), .B0(oc8051_sfr1_oc8051_uatr1_n64), .B1(
        wr_dat[3]), .Y(oc8051_sfr1_oc8051_uatr1_n68) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u57 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n67), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n65), .C0(
        oc8051_sfr1_oc8051_uatr1_n68), .Y(oc8051_sfr1_oc8051_uatr1_n238) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u56 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_), .Y(oc8051_sfr1_oc8051_uatr1_n61) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u55 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_uatr1_n63), .B0(wr_dat[2]), .B1(
        oc8051_sfr1_oc8051_uatr1_n64), .Y(oc8051_sfr1_oc8051_uatr1_n66) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u54 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n65), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n61), .C0(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n239) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u53 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_), .Y(oc8051_sfr1_oc8051_uatr1_n57) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u52 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n63), .A1(wr_dat[0]), .B0(wr_dat[1]), .B1(
        oc8051_sfr1_oc8051_uatr1_n64), .Y(oc8051_sfr1_oc8051_uatr1_n62) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u51 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n61), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .B1(oc8051_sfr1_oc8051_uatr1_n57), .C0(
        oc8051_sfr1_oc8051_uatr1_n62), .Y(oc8051_sfr1_oc8051_uatr1_n240) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u50 ( .A(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_uatr1_n59) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u49 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n56), .A1(oc8051_sfr1_oc8051_uatr1_n57), .B0(
        oc8051_sfr1_oc8051_uatr1_n58), .B1(oc8051_sfr1_oc8051_uatr1_n59), .C0(
        oc8051_sfr1_oc8051_uatr1_n38), .C1(oc8051_sfr1_oc8051_uatr1_n60), .Y(
        oc8051_sfr1_oc8051_uatr1_n241) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u48 ( .A(
        oc8051_sfr1_oc8051_uatr1_n37), .B(oc8051_sfr1_oc8051_uatr1_n55), .Y(
        oc8051_sfr1_oc8051_uatr1_n49) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u47 ( .A(
        oc8051_sfr1_oc8051_uatr1_n49), .B(oc8051_sfr1_oc8051_uatr1_n37), .C(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .Y(oc8051_sfr1_oc8051_uatr1_n50) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u46 ( .A(
        oc8051_sfr1_oc8051_uatr1_n50), .Y(oc8051_sfr1_oc8051_uatr1_n45) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u45 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .B(oc8051_sfr1_oc8051_uatr1_n45), .Y(oc8051_sfr1_oc8051_uatr1_n52) );
  OA21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u44 ( .A0(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .A1(
        oc8051_sfr1_oc8051_uatr1_n54), .B0(oc8051_sfr1_oc8051_uatr1_n49), .Y(
        oc8051_sfr1_oc8051_uatr1_n51) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u43 ( .A0(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .A1(
        oc8051_sfr1_oc8051_uatr1_n54), .B0(oc8051_sfr1_oc8051_uatr1_n51), .Y(
        oc8051_sfr1_oc8051_uatr1_n47) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u42 ( .A(
        oc8051_sfr1_oc8051_uatr1_n47), .Y(oc8051_sfr1_oc8051_uatr1_n53) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u41 ( .A(
        oc8051_sfr1_oc8051_uatr1_n52), .B(oc8051_sfr1_oc8051_uatr1_n53), .S0(
        oc8051_sfr1_oc8051_uatr1_tr_count_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n242) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u40 ( .A(
        oc8051_sfr1_oc8051_uatr1_n50), .B(oc8051_sfr1_oc8051_uatr1_n51), .S0(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .Y(
        oc8051_sfr1_oc8051_uatr1_n243) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u39 ( .A(
        oc8051_sfr1_oc8051_uatr1_n49), .B(oc8051_sfr1_oc8051_uatr1_n37), .Y(
        oc8051_sfr1_oc8051_uatr1_n48) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u38 ( .A(
        oc8051_sfr1_oc8051_uatr1_n48), .B(oc8051_sfr1_oc8051_uatr1_n49), .S0(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n244) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u37 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n37), .A1(oc8051_sfr1_oc8051_uatr1_n46), .B0(
        oc8051_sfr1_oc8051_uatr1_n47), .Y(oc8051_sfr1_oc8051_uatr1_n43) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u36 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .B(oc8051_sfr1_oc8051_uatr1_n45), .C(oc8051_sfr1_oc8051_uatr1_tr_count_2_), .Y(oc8051_sfr1_oc8051_uatr1_n44)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u35 ( .A(
        oc8051_sfr1_oc8051_uatr1_n43), .B(oc8051_sfr1_oc8051_uatr1_n44), .S0(
        oc8051_sfr1_oc8051_uatr1_n201), .Y(oc8051_sfr1_oc8051_uatr1_n245) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u34 ( .A(
        oc8051_sfr1_oc8051_uatr1_n42), .B(oc8051_sfr1_oc8051_uatr1_n8), .Y(
        oc8051_sfr1_oc8051_uatr1_n40) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u33 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n41), .B(oc8051_sfr1_oc8051_uatr1_n7), .Y(
        oc8051_sfr1_oc8051_uatr1_n9) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u32 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n39), .A1(oc8051_sfr1_oc8051_uatr1_n40), .A2(
        oc8051_sfr1_oc8051_uatr1_n9), .B0(oc8051_sfr1_oc8051_uatr1_n37), .Y(
        oc8051_sfr1_oc8051_uatr1_n246) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u31 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n34), .A1(oc8051_sfr1_oc8051_uatr1_n37), .B0(
        oc8051_sfr1_oc8051_uatr1_n199), .B1(oc8051_sfr1_oc8051_uatr1_n38), .Y(
        oc8051_sfr1_oc8051_uatr1_n247) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u30 ( .A(
        oc8051_sfr1_oc8051_uatr1_n35), .B(oc8051_sfr1_oc8051_uatr1_n36), .Y(
        oc8051_sfr1_oc8051_uatr1_n23) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u29 ( .A(
        oc8051_sfr1_oc8051_uatr1_n23), .B(oc8051_sfr1_oc8051_uatr1_n16), .Y(
        oc8051_sfr1_oc8051_uatr1_n31) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u28 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n31), .B(oc8051_sfr1_oc8051_uatr1_n34), .Y(
        oc8051_sfr1_oc8051_uatr1_n33) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u27 ( .A(
        oc8051_sfr1_oc8051_uatr1_n33), .B(wr_dat[7]), .S0(
        oc8051_sfr1_oc8051_uatr1_n14), .Y(oc8051_sfr1_oc8051_uatr1_n32) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u26 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n11), .A1(oc8051_sfr1_oc8051_uatr1_n31), .B0(
        oc8051_sfr1_oc8051_uatr1_n32), .Y(oc8051_sfr1_oc8051_uatr1_n248) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u25 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_uatr1_n21), .C(oc8051_sfr1_oc8051_uatr1_n23), .Y(
        oc8051_sfr1_oc8051_uatr1_n27) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u24 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n27), .B(oc8051_sfr1_oc8051_uatr1_n30), .Y(
        oc8051_sfr1_oc8051_uatr1_n29) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u23 ( .A(
        oc8051_sfr1_oc8051_uatr1_n29), .B(wr_dat[6]), .S0(
        oc8051_sfr1_oc8051_uatr1_n14), .Y(oc8051_sfr1_oc8051_uatr1_n28) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u22 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n11), .A1(oc8051_sfr1_oc8051_uatr1_n27), .B0(
        oc8051_sfr1_oc8051_uatr1_n28), .Y(oc8051_sfr1_oc8051_uatr1_n249) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u21 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_uatr1_n22), .C(oc8051_sfr1_oc8051_uatr1_n23), .Y(
        oc8051_sfr1_oc8051_uatr1_n24) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u20 ( .A(
        oc8051_sfr1_oc8051_uatr1_n24), .B(oc8051_sfr1_scon_5_), .Y(
        oc8051_sfr1_oc8051_uatr1_n26) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u19 ( .A(
        oc8051_sfr1_oc8051_uatr1_n26), .B(wr_dat[5]), .S0(
        oc8051_sfr1_oc8051_uatr1_n14), .Y(oc8051_sfr1_oc8051_uatr1_n25) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u18 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n11), .A1(oc8051_sfr1_oc8051_uatr1_n24), .B0(
        oc8051_sfr1_oc8051_uatr1_n25), .Y(oc8051_sfr1_oc8051_uatr1_n250) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u17 ( .A(
        oc8051_sfr1_oc8051_uatr1_n21), .B(oc8051_sfr1_oc8051_uatr1_n22), .C(
        oc8051_sfr1_oc8051_uatr1_n23), .Y(oc8051_sfr1_oc8051_uatr1_n17) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u16 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n17), .B(oc8051_sfr1_oc8051_uatr1_n20), .Y(
        oc8051_sfr1_oc8051_uatr1_n19) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u15 ( .A(
        oc8051_sfr1_oc8051_uatr1_n19), .B(wr_dat[4]), .S0(
        oc8051_sfr1_oc8051_uatr1_n14), .Y(oc8051_sfr1_oc8051_uatr1_n18) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u14 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n11), .A1(oc8051_sfr1_oc8051_uatr1_n17), .B0(
        oc8051_sfr1_oc8051_uatr1_n18), .Y(oc8051_sfr1_oc8051_uatr1_n251) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u13 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n15), .B(oc8051_sfr1_oc8051_uatr1_n16), .Y(
        oc8051_sfr1_oc8051_uatr1_n10) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u12 ( .A(
        oc8051_sfr1_oc8051_uatr1_n10), .B(oc8051_sfr1_scon_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n13) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u11 ( .A(
        oc8051_sfr1_oc8051_uatr1_n13), .B(wr_dat[3]), .S0(
        oc8051_sfr1_oc8051_uatr1_n14), .Y(oc8051_sfr1_oc8051_uatr1_n12) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u10 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n10), .A1(oc8051_sfr1_oc8051_uatr1_n11), .B0(
        oc8051_sfr1_oc8051_uatr1_n12), .Y(oc8051_sfr1_oc8051_uatr1_n252) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u9 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n8), .B(oc8051_sfr1_oc8051_uatr1_n9), .Y(
        oc8051_sfr1_oc8051_uatr1_n3) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u8 ( .A(
        oc8051_sfr1_oc8051_uatr1_n5), .B(oc8051_sfr1_oc8051_uatr1_n6), .C(
        oc8051_sfr1_oc8051_uatr1_n7), .Y(oc8051_sfr1_oc8051_uatr1_n4) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u7 ( .A(
        oc8051_sfr1_oc8051_uatr1_n3), .B(oc8051_sfr1_oc8051_uatr1_n198), .S0(
        oc8051_sfr1_oc8051_uatr1_n4), .Y(oc8051_sfr1_oc8051_uatr1_n253) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u6 ( .A(
        oc8051_sfr1_oc8051_uatr1_n2), .B(oc8051_sfr1_pcon[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n1) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u5 ( .A(
        oc8051_sfr1_oc8051_uatr1_smod_clk_tr), .B(oc8051_sfr1_oc8051_uatr1_n1), 
        .Y(oc8051_sfr1_oc8051_uatr1_n254) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u4 ( .A(wb_rst_i), .Y(
        oc8051_sfr1_oc8051_uatr1_n168) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u3 ( .A(
        oc8051_sfr1_oc8051_uatr1_n180), .Y(oc8051_sfr1_scon_1_) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n224), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n180) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tx_done_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n253), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n198) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_9_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n232), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n200) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_10_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n247), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n199) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n245), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n201) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rx_done_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n225), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_uatr1_n168), .Q(oc8051_sfr1_oc8051_uatr1_rx_done)
         );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n215), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n203) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n214), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n202) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n226), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n204) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_t1_ow_buf_reg ( .D(
        oc8051_sfr1_tf1), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n205) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n248), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n251), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n243), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n219), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n197), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n244), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n218), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n249), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n223), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_receive_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n221), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_receive) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n252), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n250), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n242), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_tr_count_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n216), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n217), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n222), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_smod_clk_tr_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n254), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_smod_clk_tr) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_smod_clk_re_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n230), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_smod_clk_re) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rx_sam_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n228), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_rx_sam_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_trans_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n246), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_trans) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_11_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n227), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n239), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n237), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_8_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n233), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rx_sam_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n229), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_rx_sam_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n240), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_shift_re_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n269), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_shift_re) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n238), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n236), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n213), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n212), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n211), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n210), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n209), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_8_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n207), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_9_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n208), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_10_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n206), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n181), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n182), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n183), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n184), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n185), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n186), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n187), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n188), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n190), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n191), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n192), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n193), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n194), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n195), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n196), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n241), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n235), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n234), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_shift_tr_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n174), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_shift_tr) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rxd_r_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n220), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_uatr1_n168), .Q(oc8051_sfr1_oc8051_uatr1_rxd_r) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_txd_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n231), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_uatr1_n168), .Q(txd_o) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u245 ( .A(oc8051_sfr1_oc8051_int1_n8), .Y(int_src[5]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u244 ( .A(oc8051_sfr1_oc8051_int1_n7), .Y(int_src[4]) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u243 ( .A(int_src[5]), .B(
        int_src[4]), .Y(oc8051_sfr1_oc8051_int1_n204) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u242 ( .A(
        oc8051_sfr1_oc8051_int1_n4), .B(oc8051_sfr1_oc8051_int1_n5), .C(
        oc8051_sfr1_oc8051_int1_n204), .D(oc8051_sfr1_oc8051_int1_n6), .Y(intr) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u241 ( .A(reti), .B(
        oc8051_sfr1_oc8051_int1_int_proc), .Y(oc8051_sfr1_oc8051_int1_n115) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u240 ( .A(oc8051_sfr1_ie_0_), .B(
        oc8051_sfr1_ip_0_), .C(oc8051_sfr1_tcon_1_), .Y(
        oc8051_sfr1_oc8051_int1_n179) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u239 ( .A(oc8051_sfr1_tcon_5_), 
        .B(oc8051_sfr1_ie_1_), .Y(oc8051_sfr1_oc8051_int1_n176) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u238 ( .A(
        oc8051_sfr1_oc8051_int1_n176), .Y(oc8051_sfr1_oc8051_int1_n183) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u237 ( .A(
        oc8051_sfr1_oc8051_int1_n183), .B(oc8051_sfr1_ip_1_), .Y(
        oc8051_sfr1_oc8051_int1_n178) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u236 ( .A(oc8051_sfr1_ie_2_), .B(
        oc8051_sfr1_ip_2_), .C(oc8051_sfr1_tcon_3_), .Y(
        oc8051_sfr1_oc8051_int1_n203) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u235 ( .A(
        oc8051_sfr1_oc8051_int1_n179), .B(oc8051_sfr1_oc8051_int1_n178), .C(
        oc8051_sfr1_oc8051_int1_n203), .Y(oc8051_sfr1_oc8051_int1_n195) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u234 ( .A(oc8051_sfr1_tcon_7_), 
        .B(oc8051_sfr1_ie_3_), .Y(oc8051_sfr1_oc8051_int1_n190) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u233 ( .A(oc8051_sfr1_ip_3_), .Y(
        oc8051_sfr1_oc8051_int1_n30) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u232 ( .A(
        oc8051_sfr1_oc8051_int1_n190), .B(oc8051_sfr1_oc8051_int1_n30), .Y(
        oc8051_sfr1_oc8051_int1_n196) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u231 ( .AN(
        oc8051_sfr1_oc8051_int1_n195), .B(oc8051_sfr1_oc8051_int1_n196), .Y(
        oc8051_sfr1_oc8051_int1_n189) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u230 ( .A(oc8051_sfr1_tc2_int), .Y(
        oc8051_sfr1_oc8051_int1_n192) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u229 ( .A(oc8051_sfr1_ie_5_), .Y(
        oc8051_sfr1_oc8051_int1_n61) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u228 ( .A(oc8051_sfr1_ie_4_), .B(
        oc8051_sfr1_ip_4_), .C(oc8051_sfr1_uart_int), .Y(
        oc8051_sfr1_oc8051_int1_n188) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u227 ( .A0(
        oc8051_sfr1_oc8051_int1_n192), .A1(oc8051_sfr1_oc8051_int1_n11), .A2(
        oc8051_sfr1_oc8051_int1_n61), .B0(oc8051_sfr1_oc8051_int1_n188), .Y(
        oc8051_sfr1_oc8051_int1_n200) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u226 ( .A(oc8051_sfr1_ie_7_), .Y(
        oc8051_sfr1_oc8051_int1_n50) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u225 ( .A(
        oc8051_sfr1_oc8051_int1_int_lev_1__0_), .Y(
        oc8051_sfr1_oc8051_int1_n151) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u224 ( .A(
        oc8051_sfr1_oc8051_int1_int_lev_0__0_), .Y(
        oc8051_sfr1_oc8051_int1_n148) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u223 ( .A(
        oc8051_sfr1_oc8051_int1_n151), .B(oc8051_sfr1_oc8051_int1_n148), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n202)
         );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u222 ( .A0(
        oc8051_sfr1_oc8051_int1_n50), .A1(oc8051_sfr1_oc8051_int1_n202), .B0(
        oc8051_sfr1_oc8051_int1_int_proc), .Y(oc8051_sfr1_oc8051_int1_n201) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u221 ( .A1N(
        oc8051_sfr1_oc8051_int1_n189), .A0(oc8051_sfr1_oc8051_int1_n200), .B0(
        oc8051_sfr1_oc8051_int1_n201), .Y(oc8051_sfr1_oc8051_int1_n197) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u220 ( .A(
        oc8051_sfr1_oc8051_int1_n115), .B(oc8051_sfr1_oc8051_int1_n197), .Y(
        oc8051_sfr1_oc8051_int1_n112) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u219 ( .A(
        oc8051_sfr1_oc8051_int1_n112), .Y(oc8051_sfr1_oc8051_int1_n146) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u218 ( .A(
        oc8051_sfr1_oc8051_int1_n190), .Y(oc8051_sfr1_oc8051_int1_n199) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u217 ( .A(oc8051_sfr1_ie_2_), .Y(
        oc8051_sfr1_oc8051_int1_n70) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u216 ( .A(oc8051_sfr1_tcon_3_), .Y(
        oc8051_sfr1_oc8051_int1_n139) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u215 ( .A(oc8051_sfr1_tcon_1_), .Y(
        oc8051_sfr1_oc8051_int1_n130) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u214 ( .A(oc8051_sfr1_ie_0_), .Y(
        oc8051_sfr1_oc8051_int1_n77) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u213 ( .A(
        oc8051_sfr1_oc8051_int1_n130), .B(oc8051_sfr1_oc8051_int1_n77), .Y(
        oc8051_sfr1_oc8051_int1_n175) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u212 ( .A(
        oc8051_sfr1_oc8051_int1_n175), .Y(oc8051_sfr1_oc8051_int1_n180) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u211 ( .A0(
        oc8051_sfr1_oc8051_int1_n70), .A1(oc8051_sfr1_oc8051_int1_n139), .B0(
        oc8051_sfr1_oc8051_int1_n180), .C0(oc8051_sfr1_oc8051_int1_n176), .Y(
        oc8051_sfr1_oc8051_int1_n186) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u210 ( .A0(oc8051_sfr1_ie_4_), 
        .A1(oc8051_sfr1_uart_int), .B0(oc8051_sfr1_oc8051_int1_n199), .C0(
        oc8051_sfr1_oc8051_int1_n186), .Y(oc8051_sfr1_oc8051_int1_n193) );
  OA21A1OI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u209 ( .A0(
        oc8051_sfr1_oc8051_int1_n61), .A1(oc8051_sfr1_oc8051_int1_n192), .B0(
        oc8051_sfr1_oc8051_int1_n193), .C0(oc8051_sfr1_oc8051_int1_int_proc), 
        .Y(oc8051_sfr1_oc8051_int1_n198) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u208 ( .A(
        oc8051_sfr1_oc8051_int1_n146), .B(oc8051_sfr1_ie_7_), .C(
        oc8051_sfr1_oc8051_int1_n198), .Y(oc8051_sfr1_oc8051_int1_n174) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u207 ( .A(
        oc8051_sfr1_oc8051_int1_n115), .Y(oc8051_sfr1_oc8051_int1_n116) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u206 ( .A(
        oc8051_sfr1_oc8051_int1_n197), .B(oc8051_sfr1_oc8051_int1_n116), .Y(
        oc8051_sfr1_oc8051_int1_n150) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u205 ( .A(
        oc8051_sfr1_oc8051_int1_n150), .B(oc8051_sfr1_oc8051_int1_n195), .C(
        oc8051_sfr1_oc8051_int1_n196), .Y(oc8051_sfr1_oc8051_int1_n194) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u204 ( .A0(
        oc8051_sfr1_oc8051_int1_n174), .A1(oc8051_sfr1_oc8051_int1_n190), .A2(
        oc8051_sfr1_oc8051_int1_n186), .B0(oc8051_sfr1_oc8051_int1_n194), .Y(
        oc8051_sfr1_oc8051_int1_n156) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u203 ( .A(
        oc8051_sfr1_oc8051_int1_n156), .Y(oc8051_sfr1_oc8051_int1_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u202 ( .A(
        oc8051_sfr1_oc8051_int1_n174), .Y(oc8051_sfr1_oc8051_int1_n147) );
  AOI32_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u201 ( .A0(
        oc8051_sfr1_oc8051_int1_n189), .A1(oc8051_sfr1_oc8051_int1_n188), .A2(
        oc8051_sfr1_oc8051_int1_n150), .B0(oc8051_sfr1_oc8051_int1_n147), .B1(
        oc8051_sfr1_oc8051_int1_n193), .Y(oc8051_sfr1_oc8051_int1_n191) );
  OR3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u200 ( .A(
        oc8051_sfr1_oc8051_int1_n191), .B(oc8051_sfr1_oc8051_int1_n61), .C(
        oc8051_sfr1_oc8051_int1_n192), .Y(oc8051_sfr1_oc8051_int1_n154) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u199 ( .A(oc8051_sfr1_ie_4_), .B(
        oc8051_sfr1_oc8051_int1_n190), .C(oc8051_sfr1_uart_int), .Y(
        oc8051_sfr1_oc8051_int1_n185) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u198 ( .AN(
        oc8051_sfr1_oc8051_int1_n188), .B(oc8051_sfr1_oc8051_int1_n150), .C(
        oc8051_sfr1_oc8051_int1_n189), .Y(oc8051_sfr1_oc8051_int1_n187) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u197 ( .A0(
        oc8051_sfr1_oc8051_int1_n185), .A1(oc8051_sfr1_oc8051_int1_n186), .A2(
        oc8051_sfr1_oc8051_int1_n174), .B0(oc8051_sfr1_oc8051_int1_n187), .Y(
        oc8051_sfr1_oc8051_int1_n171) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u196 ( .A(
        oc8051_sfr1_oc8051_int1_n171), .Y(oc8051_sfr1_oc8051_int1_n160) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u195 ( .A(
        oc8051_sfr1_oc8051_int1_n159), .B(oc8051_sfr1_oc8051_int1_n154), .C(
        oc8051_sfr1_oc8051_int1_n160), .Y(oc8051_sfr1_oc8051_int1_n167) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u194 ( .A(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n144)
         );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u193 ( .A(
        oc8051_sfr1_oc8051_int1_n144), .B(oc8051_sfr1_oc8051_int1_int_dept_1_), 
        .Y(oc8051_sfr1_oc8051_int1_n114) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u192 ( .A(
        oc8051_sfr1_oc8051_int1_n150), .Y(oc8051_sfr1_oc8051_int1_n181) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u191 ( .A(
        oc8051_sfr1_oc8051_int1_n150), .B(oc8051_sfr1_ip_2_), .C(
        oc8051_sfr1_oc8051_int1_n179), .D(oc8051_sfr1_oc8051_int1_n178), .Y(
        oc8051_sfr1_oc8051_int1_n184) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u190 ( .A0(
        oc8051_sfr1_oc8051_int1_n174), .A1(oc8051_sfr1_oc8051_int1_n183), .A2(
        oc8051_sfr1_oc8051_int1_n175), .B0(oc8051_sfr1_oc8051_int1_n184), .Y(
        oc8051_sfr1_oc8051_int1_n182) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u189 ( .A(oc8051_sfr1_ie_2_), .B(
        oc8051_sfr1_oc8051_int1_n182), .C(oc8051_sfr1_tcon_3_), .Y(
        oc8051_sfr1_oc8051_int1_n158) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u188 ( .A0(
        oc8051_sfr1_oc8051_int1_n174), .A1(oc8051_sfr1_oc8051_int1_n180), .B0(
        oc8051_sfr1_oc8051_int1_n181), .B1(oc8051_sfr1_oc8051_int1_n179), .C0(
        oc8051_sfr1_oc8051_int1_n158), .Y(oc8051_sfr1_oc8051_int1_n170) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u187 ( .AN(
        oc8051_sfr1_oc8051_int1_n178), .B(oc8051_sfr1_oc8051_int1_n150), .C(
        oc8051_sfr1_oc8051_int1_n179), .Y(oc8051_sfr1_oc8051_int1_n177) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u186 ( .A0(
        oc8051_sfr1_oc8051_int1_n174), .A1(oc8051_sfr1_oc8051_int1_n175), .A2(
        oc8051_sfr1_oc8051_int1_n176), .B0(oc8051_sfr1_oc8051_int1_n177), .Y(
        oc8051_sfr1_oc8051_int1_n157) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u185 ( .A(
        oc8051_sfr1_oc8051_int1_n157), .Y(oc8051_sfr1_oc8051_int1_n173) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u184 ( .AN(
        oc8051_sfr1_oc8051_int1_n170), .B(oc8051_sfr1_oc8051_int1_n173), .C(
        oc8051_sfr1_oc8051_int1_n167), .Y(oc8051_sfr1_oc8051_int1_n161) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u183 ( .A(
        oc8051_sfr1_oc8051_int1_n114), .B(oc8051_sfr1_oc8051_int1_n161), .Y(
        oc8051_sfr1_oc8051_int1_n169) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u182 ( .A(
        oc8051_sfr1_oc8051_int1_n10), .B(oc8051_sfr1_oc8051_int1_n167), .S0(
        oc8051_sfr1_oc8051_int1_n169), .Y(oc8051_sfr1_oc8051_int1_n226) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u181 ( .A(
        oc8051_sfr1_oc8051_int1_isrc_1__1_), .Y(oc8051_sfr1_oc8051_int1_n172)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u180 ( .A(
        oc8051_sfr1_oc8051_int1_n158), .B(oc8051_sfr1_oc8051_int1_n154), .C(
        oc8051_sfr1_oc8051_int1_n173), .Y(oc8051_sfr1_oc8051_int1_n166) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u179 ( .A(
        oc8051_sfr1_oc8051_int1_n172), .B(oc8051_sfr1_oc8051_int1_n166), .S0(
        oc8051_sfr1_oc8051_int1_n169), .Y(oc8051_sfr1_oc8051_int1_n227) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u178 ( .A(
        oc8051_sfr1_oc8051_int1_isrc_1__0_), .Y(oc8051_sfr1_oc8051_int1_n168)
         );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u177 ( .A(
        oc8051_sfr1_oc8051_int1_n170), .B(oc8051_sfr1_oc8051_int1_n171), .Y(
        oc8051_sfr1_oc8051_int1_n163) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u176 ( .A(
        oc8051_sfr1_oc8051_int1_n168), .B(oc8051_sfr1_oc8051_int1_n163), .S0(
        oc8051_sfr1_oc8051_int1_n169), .Y(oc8051_sfr1_oc8051_int1_n228) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u175 ( .A(
        oc8051_sfr1_oc8051_int1_int_dept_1_), .B(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n113)
         );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u174 ( .A(
        oc8051_sfr1_oc8051_int1_n113), .B(oc8051_sfr1_oc8051_int1_n161), .Y(
        oc8051_sfr1_oc8051_int1_n164) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u173 ( .A(
        oc8051_sfr1_oc8051_int1_n9), .B(oc8051_sfr1_oc8051_int1_n167), .S0(
        oc8051_sfr1_oc8051_int1_n164), .Y(oc8051_sfr1_oc8051_int1_n229) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u172 ( .A(
        oc8051_sfr1_oc8051_int1_isrc_0__1_), .Y(oc8051_sfr1_oc8051_int1_n165)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u171 ( .A(
        oc8051_sfr1_oc8051_int1_n165), .B(oc8051_sfr1_oc8051_int1_n166), .S0(
        oc8051_sfr1_oc8051_int1_n164), .Y(oc8051_sfr1_oc8051_int1_n230) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u170 ( .A(
        oc8051_sfr1_oc8051_int1_isrc_0__0_), .Y(oc8051_sfr1_oc8051_int1_n162)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u169 ( .A(
        oc8051_sfr1_oc8051_int1_n162), .B(oc8051_sfr1_oc8051_int1_n163), .S0(
        oc8051_sfr1_oc8051_int1_n164), .Y(oc8051_sfr1_oc8051_int1_n231) );
  OR2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u168 ( .A(
        oc8051_sfr1_oc8051_int1_n161), .B(oc8051_sfr1_oc8051_int1_n146), .Y(
        oc8051_sfr1_oc8051_int1_n153) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u167 ( .A0(
        oc8051_sfr1_oc8051_int1_n8), .A1(oc8051_sfr1_oc8051_int1_n153), .B0(
        oc8051_sfr1_oc8051_int1_n154), .C0(oc8051_sfr1_oc8051_int1_n160), .Y(
        oc8051_sfr1_oc8051_int1_n232) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u166 ( .A0(
        oc8051_sfr1_oc8051_int1_n7), .A1(oc8051_sfr1_oc8051_int1_n153), .B0(
        oc8051_sfr1_oc8051_int1_n158), .C0(oc8051_sfr1_oc8051_int1_n159), .Y(
        oc8051_sfr1_oc8051_int1_n233) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u165 ( .A(
        oc8051_sfr1_oc8051_int1_n156), .B(oc8051_sfr1_oc8051_int1_n157), .Y(
        oc8051_sfr1_oc8051_int1_n155) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u164 ( .A0(
        oc8051_sfr1_oc8051_int1_n6), .A1(oc8051_sfr1_oc8051_int1_n153), .B0(
        oc8051_sfr1_oc8051_int1_n154), .C0(oc8051_sfr1_oc8051_int1_n155), .Y(
        oc8051_sfr1_oc8051_int1_n234) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u163 ( .A(
        oc8051_sfr1_oc8051_int1_n150), .B(oc8051_sfr1_oc8051_int1_n147), .Y(
        oc8051_sfr1_oc8051_int1_n117) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u162 ( .A0(
        oc8051_sfr1_oc8051_int1_n5), .A1(oc8051_sfr1_oc8051_int1_n153), .B0(
        oc8051_sfr1_oc8051_int1_n117), .Y(oc8051_sfr1_oc8051_int1_n235) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u161 ( .A0(
        oc8051_sfr1_oc8051_int1_n4), .A1(oc8051_sfr1_oc8051_int1_n153), .B0(
        oc8051_sfr1_oc8051_int1_n117), .Y(oc8051_sfr1_oc8051_int1_n236) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u160 ( .A(
        oc8051_sfr1_oc8051_int1_n150), .B(oc8051_sfr1_oc8051_int1_n114), .Y(
        oc8051_sfr1_oc8051_int1_n152) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u159 ( .A0(
        oc8051_sfr1_oc8051_int1_n147), .A1(oc8051_sfr1_oc8051_int1_n114), .B0(
        oc8051_sfr1_oc8051_int1_n151), .C0(oc8051_sfr1_oc8051_int1_n152), .Y(
        oc8051_sfr1_oc8051_int1_n237) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u158 ( .A(
        oc8051_sfr1_oc8051_int1_n150), .B(oc8051_sfr1_oc8051_int1_n113), .Y(
        oc8051_sfr1_oc8051_int1_n149) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u157 ( .A0(
        oc8051_sfr1_oc8051_int1_n147), .A1(oc8051_sfr1_oc8051_int1_n113), .B0(
        oc8051_sfr1_oc8051_int1_n148), .C0(oc8051_sfr1_oc8051_int1_n149), .Y(
        oc8051_sfr1_oc8051_int1_n238) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u156 ( .A(
        oc8051_sfr1_oc8051_int1_n146), .B(oc8051_sfr1_oc8051_int1_n144), .Y(
        oc8051_sfr1_oc8051_int1_n145) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u155 ( .A(
        oc8051_sfr1_oc8051_int1_n117), .B(oc8051_sfr1_oc8051_int1_n115), .Y(
        oc8051_sfr1_oc8051_int1_n108) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u154 ( .A(
        oc8051_sfr1_oc8051_int1_n144), .B(oc8051_sfr1_oc8051_int1_n145), .S0(
        oc8051_sfr1_oc8051_int1_n108), .Y(oc8051_sfr1_oc8051_int1_n239) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u153 ( .A(wr_addr[4]), .B(
        wr_addr[6]), .C(wr_addr[5]), .Y(oc8051_sfr1_oc8051_int1_n143) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u152 ( .A(wr_addr[7]), .B(n_5_net_), 
        .C(wr_addr[3]), .D(oc8051_sfr1_oc8051_int1_n143), .Y(
        oc8051_sfr1_oc8051_int1_n142) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u151 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n41) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u150 ( .A(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_int1_n46) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u149 ( .A(wr_addr[2]), .B(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_int1_n39) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u148 ( .A(
        oc8051_sfr1_oc8051_int1_n41), .B(oc8051_sfr1_oc8051_int1_n46), .C(
        oc8051_sfr1_oc8051_int1_n39), .Y(oc8051_sfr1_oc8051_int1_n79) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u147 ( .A(
        oc8051_sfr1_oc8051_int1_n142), .B(oc8051_sfr1_oc8051_int1_n79), .Y(
        oc8051_sfr1_oc8051_int1_n85) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u146 ( .A1N(
        oc8051_sfr1_oc8051_int1_ie1_buff), .A0(oc8051_sfr1_tcon_2_), .B0(
        int1_i), .Y(oc8051_sfr1_oc8051_int1_n141) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u145 ( .AN(
        oc8051_sfr1_oc8051_int1_n142), .B(oc8051_sfr1_oc8051_int1_n46), .Y(
        oc8051_sfr1_oc8051_int1_n98) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u144 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_int1_n100) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u143 ( .A(
        oc8051_sfr1_oc8051_int1_n100), .B(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_int1_n32) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u142 ( .A(
        oc8051_sfr1_oc8051_int1_n98), .B(oc8051_sfr1_oc8051_int1_n32), .Y(
        oc8051_sfr1_oc8051_int1_n89) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u141 ( .AN(
        oc8051_sfr1_oc8051_int1_n89), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n140) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u140 ( .A(descy), .B(
        oc8051_sfr1_oc8051_int1_n141), .S0(oc8051_sfr1_oc8051_int1_n140), .Y(
        oc8051_sfr1_oc8051_int1_n134) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u139 ( .A(
        oc8051_sfr1_oc8051_int1_n10), .B(oc8051_sfr1_oc8051_int1_n9), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n106)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u138 ( .A(
        oc8051_sfr1_oc8051_int1_int_proc), .Y(oc8051_sfr1_oc8051_int1_n104) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u137 ( .A(int_ack), .Y(
        oc8051_sfr1_oc8051_int1_n103) );
  OR3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u136 ( .A(
        oc8051_sfr1_oc8051_int1_n106), .B(oc8051_sfr1_oc8051_int1_n104), .C(
        oc8051_sfr1_oc8051_int1_n103), .Y(oc8051_sfr1_oc8051_int1_n123) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u135 ( .A(
        oc8051_sfr1_oc8051_int1_isrc_1__1_), .B(
        oc8051_sfr1_oc8051_int1_isrc_0__1_), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n107)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u134 ( .A(
        oc8051_sfr1_oc8051_int1_isrc_1__0_), .B(
        oc8051_sfr1_oc8051_int1_isrc_0__0_), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n105)
         );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u133 ( .A0(
        oc8051_sfr1_oc8051_int1_n123), .A1(oc8051_sfr1_oc8051_int1_n107), .A2(
        oc8051_sfr1_oc8051_int1_n105), .B0(oc8051_sfr1_oc8051_int1_n140), .Y(
        oc8051_sfr1_oc8051_int1_n137) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u132 ( .A(oc8051_sfr1_tcon_2_), .Y(
        oc8051_sfr1_oc8051_int1_n138) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u131 ( .A(
        oc8051_sfr1_oc8051_int1_n137), .B(oc8051_sfr1_oc8051_int1_n138), .C(
        oc8051_sfr1_oc8051_int1_n139), .Y(oc8051_sfr1_oc8051_int1_n136) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u130 ( .A(
        oc8051_sfr1_oc8051_int1_n136), .B(wr_dat[3]), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n135) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u129 ( .A0(
        oc8051_sfr1_oc8051_int1_n85), .A1(oc8051_sfr1_oc8051_int1_n134), .B0(
        oc8051_sfr1_oc8051_int1_n135), .Y(oc8051_sfr1_oc8051_int1_n240) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u128 ( .A1N(
        oc8051_sfr1_oc8051_int1_ie0_buff), .A0(oc8051_sfr1_tcon_0_), .B0(
        int0_i), .Y(oc8051_sfr1_oc8051_int1_n133) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u127 ( .A(
        oc8051_sfr1_oc8051_int1_n98), .B(oc8051_sfr1_oc8051_int1_n39), .Y(
        oc8051_sfr1_oc8051_int1_n92) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u126 ( .AN(
        oc8051_sfr1_oc8051_int1_n92), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n132) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u125 ( .A(descy), .B(
        oc8051_sfr1_oc8051_int1_n133), .S0(oc8051_sfr1_oc8051_int1_n132), .Y(
        oc8051_sfr1_oc8051_int1_n125) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u124 ( .A(
        oc8051_sfr1_oc8051_int1_n107), .Y(oc8051_sfr1_oc8051_int1_n131) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u123 ( .A0(
        oc8051_sfr1_oc8051_int1_n123), .A1(oc8051_sfr1_oc8051_int1_n105), .A2(
        oc8051_sfr1_oc8051_int1_n131), .B0(oc8051_sfr1_oc8051_int1_n132), .Y(
        oc8051_sfr1_oc8051_int1_n128) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u122 ( .A(oc8051_sfr1_tcon_0_), .Y(
        oc8051_sfr1_oc8051_int1_n129) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u121 ( .A(
        oc8051_sfr1_oc8051_int1_n128), .B(oc8051_sfr1_oc8051_int1_n129), .C(
        oc8051_sfr1_oc8051_int1_n130), .Y(oc8051_sfr1_oc8051_int1_n127) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u120 ( .A(
        oc8051_sfr1_oc8051_int1_n127), .B(wr_dat[1]), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n126) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u119 ( .A0(
        oc8051_sfr1_oc8051_int1_n85), .A1(oc8051_sfr1_oc8051_int1_n125), .B0(
        oc8051_sfr1_oc8051_int1_n126), .Y(oc8051_sfr1_oc8051_int1_n241) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u118 ( .A(
        oc8051_sfr1_oc8051_int1_n105), .Y(oc8051_sfr1_oc8051_int1_n124) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u117 ( .A0(
        oc8051_sfr1_oc8051_int1_n123), .A1(oc8051_sfr1_oc8051_int1_n107), .A2(
        oc8051_sfr1_oc8051_int1_n124), .B0(oc8051_sfr1_tcon_5_), .Y(
        oc8051_sfr1_oc8051_int1_n122) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u116 ( .A1N(oc8051_sfr1_tf0), 
        .A0(oc8051_sfr1_oc8051_int1_tf0_buff), .B0(
        oc8051_sfr1_oc8051_int1_n122), .Y(oc8051_sfr1_oc8051_int1_n120) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u115 ( .A(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_int1_n99) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u114 ( .A(
        oc8051_sfr1_oc8051_int1_n99), .B(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_int1_n24) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u113 ( .A(
        oc8051_sfr1_oc8051_int1_n98), .B(oc8051_sfr1_oc8051_int1_n24), .Y(
        oc8051_sfr1_oc8051_int1_n86) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u112 ( .A(
        oc8051_sfr1_oc8051_int1_n41), .B(oc8051_sfr1_oc8051_int1_n86), .Y(
        oc8051_sfr1_oc8051_int1_n121) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u111 ( .A(
        oc8051_sfr1_oc8051_int1_n120), .B(descy), .S0(
        oc8051_sfr1_oc8051_int1_n121), .Y(oc8051_sfr1_oc8051_int1_n118) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u110 ( .A(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_int1_n119) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u109 ( .A(
        oc8051_sfr1_oc8051_int1_n118), .B(oc8051_sfr1_oc8051_int1_n119), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n242) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u108 ( .A0(
        oc8051_sfr1_oc8051_int1_n114), .A1(oc8051_sfr1_oc8051_int1_n116), .B0(
        oc8051_sfr1_oc8051_int1_n104), .C0(oc8051_sfr1_oc8051_int1_n117), .Y(
        oc8051_sfr1_oc8051_int1_n243) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u107 ( .A(
        oc8051_sfr1_oc8051_int1_n115), .B(oc8051_sfr1_oc8051_int1_int_dept_0_), 
        .Y(oc8051_sfr1_oc8051_int1_n110) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u106 ( .A(
        oc8051_sfr1_oc8051_int1_n113), .B(oc8051_sfr1_oc8051_int1_n114), .S0(
        oc8051_sfr1_oc8051_int1_n115), .Y(oc8051_sfr1_oc8051_int1_n111) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u105 ( .A0(
        oc8051_sfr1_oc8051_int1_n110), .A1(oc8051_sfr1_oc8051_int1_int_dept_1_), .B0(oc8051_sfr1_oc8051_int1_n111), .C0(oc8051_sfr1_oc8051_int1_n112), .Y(
        oc8051_sfr1_oc8051_int1_n109) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u104 ( .A1N(
        oc8051_sfr1_oc8051_int1_int_dept_1_), .A0(oc8051_sfr1_oc8051_int1_n108), .B0(oc8051_sfr1_oc8051_int1_n109), .Y(oc8051_sfr1_oc8051_int1_n244) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u103 ( .A(
        oc8051_sfr1_oc8051_int1_n105), .B(oc8051_sfr1_oc8051_int1_n106), .C(
        oc8051_sfr1_oc8051_int1_n107), .Y(oc8051_sfr1_oc8051_int1_n102) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u102 ( .A0(
        oc8051_sfr1_oc8051_int1_n102), .A1(oc8051_sfr1_oc8051_int1_n103), .A2(
        oc8051_sfr1_oc8051_int1_n104), .B0(oc8051_sfr1_tcon_7_), .Y(
        oc8051_sfr1_oc8051_int1_n101) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u101 ( .A1N(oc8051_sfr1_tf1), 
        .A0(oc8051_sfr1_oc8051_int1_tf1_buff), .B0(
        oc8051_sfr1_oc8051_int1_n101), .Y(oc8051_sfr1_oc8051_int1_n96) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u100 ( .A(
        oc8051_sfr1_oc8051_int1_n99), .B(oc8051_sfr1_oc8051_int1_n100), .Y(
        oc8051_sfr1_oc8051_int1_n13) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u99 ( .A(
        oc8051_sfr1_oc8051_int1_n98), .B(oc8051_sfr1_oc8051_int1_n13), .Y(
        oc8051_sfr1_oc8051_int1_n82) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u98 ( .A(
        oc8051_sfr1_oc8051_int1_n41), .B(oc8051_sfr1_oc8051_int1_n82), .Y(
        oc8051_sfr1_oc8051_int1_n97) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u97 ( .A(
        oc8051_sfr1_oc8051_int1_n96), .B(descy), .S0(
        oc8051_sfr1_oc8051_int1_n97), .Y(oc8051_sfr1_oc8051_int1_n95) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u96 ( .A(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_int1_n16) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u95 ( .A(
        oc8051_sfr1_oc8051_int1_n95), .B(oc8051_sfr1_oc8051_int1_n16), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n245) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u94 ( .A(descy), .Y(
        oc8051_sfr1_oc8051_int1_n81) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u93 ( .A(
        oc8051_sfr1_oc8051_int1_n92), .B(oc8051_sfr1_tcon_0_), .Y(
        oc8051_sfr1_oc8051_int1_n94) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u92 ( .A(
        oc8051_sfr1_oc8051_int1_n94), .B(wr_dat[0]), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n93) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u91 ( .A0(
        oc8051_sfr1_oc8051_int1_n81), .A1(oc8051_sfr1_oc8051_int1_n92), .B0(
        oc8051_sfr1_oc8051_int1_n93), .Y(oc8051_sfr1_oc8051_int1_n246) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u90 ( .A(
        oc8051_sfr1_oc8051_int1_n89), .B(oc8051_sfr1_tcon_2_), .Y(
        oc8051_sfr1_oc8051_int1_n91) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u89 ( .A(
        oc8051_sfr1_oc8051_int1_n91), .B(wr_dat[2]), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n90) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u88 ( .A0(
        oc8051_sfr1_oc8051_int1_n81), .A1(oc8051_sfr1_oc8051_int1_n89), .B0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n247) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u87 ( .A(oc8051_sfr1_tr0), .B(
        oc8051_sfr1_oc8051_int1_n86), .Y(oc8051_sfr1_oc8051_int1_n88) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u86 ( .A(
        oc8051_sfr1_oc8051_int1_n88), .B(wr_dat[4]), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n87) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u85 ( .A0(
        oc8051_sfr1_oc8051_int1_n81), .A1(oc8051_sfr1_oc8051_int1_n86), .B0(
        oc8051_sfr1_oc8051_int1_n87), .Y(oc8051_sfr1_oc8051_int1_n248) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u84 ( .A(oc8051_sfr1_tr1), .B(
        oc8051_sfr1_oc8051_int1_n82), .Y(oc8051_sfr1_oc8051_int1_n84) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u83 ( .A(
        oc8051_sfr1_oc8051_int1_n84), .B(wr_dat[6]), .S0(
        oc8051_sfr1_oc8051_int1_n85), .Y(oc8051_sfr1_oc8051_int1_n83) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u82 ( .A0(
        oc8051_sfr1_oc8051_int1_n81), .A1(oc8051_sfr1_oc8051_int1_n82), .B0(
        oc8051_sfr1_oc8051_int1_n83), .Y(oc8051_sfr1_oc8051_int1_n249) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u81 ( .A(wr_addr[6]), .Y(
        oc8051_sfr1_oc8051_int1_n80) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u80 ( .A(
        oc8051_sfr1_oc8051_int1_n80), .B(wr_addr[7]), .C(wr_addr[5]), .D(
        n_5_net_), .Y(oc8051_sfr1_oc8051_int1_n47) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u79 ( .AN(wr_addr[4]), .B(
        oc8051_sfr1_oc8051_int1_n79), .C(wr_addr[3]), .D(
        oc8051_sfr1_oc8051_int1_n47), .Y(oc8051_sfr1_oc8051_int1_n58) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u78 ( .A(oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n53) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u77 ( .A(wr_addr[3]), .B(
        oc8051_sfr1_oc8051_int1_n47), .C(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_int1_n45) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u76 ( .AN(
        oc8051_sfr1_oc8051_int1_n45), .B(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_int1_n75) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u75 ( .A(
        oc8051_sfr1_oc8051_int1_n75), .B(descy), .Y(
        oc8051_sfr1_oc8051_int1_n59) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u74 ( .A(oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n54) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u73 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[0]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n76) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u72 ( .AN(
        oc8051_sfr1_oc8051_int1_n75), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n57) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u71 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n39), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n78) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u70 ( .A(
        oc8051_sfr1_oc8051_int1_n76), .B(oc8051_sfr1_oc8051_int1_n77), .S0(
        oc8051_sfr1_oc8051_int1_n78), .Y(oc8051_sfr1_oc8051_int1_n250) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u69 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[1]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n72) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u68 ( .A(oc8051_sfr1_ie_1_), .Y(
        oc8051_sfr1_oc8051_int1_n73) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u67 ( .AN(
        oc8051_sfr1_oc8051_int1_n75), .B(oc8051_sfr1_oc8051_int1_n41), .Y(
        oc8051_sfr1_oc8051_int1_n52) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u66 ( .A0(
        oc8051_sfr1_oc8051_int1_n52), .A1(oc8051_sfr1_oc8051_int1_n39), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n74) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u65 ( .A(
        oc8051_sfr1_oc8051_int1_n72), .B(oc8051_sfr1_oc8051_int1_n73), .S0(
        oc8051_sfr1_oc8051_int1_n74), .Y(oc8051_sfr1_oc8051_int1_n251) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u64 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[2]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n69) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u63 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n32), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n71) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u62 ( .A(
        oc8051_sfr1_oc8051_int1_n69), .B(oc8051_sfr1_oc8051_int1_n70), .S0(
        oc8051_sfr1_oc8051_int1_n71), .Y(oc8051_sfr1_oc8051_int1_n252) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u61 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[3]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n66) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u60 ( .A(oc8051_sfr1_ie_3_), .Y(
        oc8051_sfr1_oc8051_int1_n67) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u59 ( .A0(
        oc8051_sfr1_oc8051_int1_n52), .A1(oc8051_sfr1_oc8051_int1_n32), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n68) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u58 ( .A(
        oc8051_sfr1_oc8051_int1_n66), .B(oc8051_sfr1_oc8051_int1_n67), .S0(
        oc8051_sfr1_oc8051_int1_n68), .Y(oc8051_sfr1_oc8051_int1_n253) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u57 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[4]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n63) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u56 ( .A(oc8051_sfr1_ie_4_), .Y(
        oc8051_sfr1_oc8051_int1_n64) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u55 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n24), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n65) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u54 ( .A(
        oc8051_sfr1_oc8051_int1_n63), .B(oc8051_sfr1_oc8051_int1_n64), .S0(
        oc8051_sfr1_oc8051_int1_n65), .Y(oc8051_sfr1_oc8051_int1_n254) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u53 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[5]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n60) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u52 ( .A0(
        oc8051_sfr1_oc8051_int1_n52), .A1(oc8051_sfr1_oc8051_int1_n24), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n62) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u51 ( .A(
        oc8051_sfr1_oc8051_int1_n60), .B(oc8051_sfr1_oc8051_int1_n61), .S0(
        oc8051_sfr1_oc8051_int1_n62), .Y(oc8051_sfr1_oc8051_int1_n255) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u50 ( .A(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_int1_n21) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u49 ( .A0(
        oc8051_sfr1_oc8051_int1_n21), .A1(oc8051_sfr1_oc8051_int1_n58), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n55) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u48 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n13), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n56) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u47 ( .A(
        oc8051_sfr1_oc8051_int1_n55), .B(oc8051_sfr1_ie_6_), .S0(
        oc8051_sfr1_oc8051_int1_n56), .Y(oc8051_sfr1_oc8051_int1_n256) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u46 ( .A0(
        oc8051_sfr1_oc8051_int1_n53), .A1(wr_dat[7]), .B0(
        oc8051_sfr1_oc8051_int1_n54), .Y(oc8051_sfr1_oc8051_int1_n49) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u45 ( .A0(
        oc8051_sfr1_oc8051_int1_n52), .A1(oc8051_sfr1_oc8051_int1_n13), .B0(
        oc8051_sfr1_oc8051_int1_n53), .Y(oc8051_sfr1_oc8051_int1_n51) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u44 ( .A(
        oc8051_sfr1_oc8051_int1_n49), .B(oc8051_sfr1_oc8051_int1_n50), .S0(
        oc8051_sfr1_oc8051_int1_n51), .Y(oc8051_sfr1_oc8051_int1_n257) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u43 ( .A(
        oc8051_sfr1_oc8051_int1_n13), .B(wr_addr[4]), .C(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n48) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u42 ( .AN(wr_addr[3]), .B(
        oc8051_sfr1_oc8051_int1_n46), .C(oc8051_sfr1_oc8051_int1_n47), .D(
        oc8051_sfr1_oc8051_int1_n48), .Y(oc8051_sfr1_oc8051_int1_n15) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u41 ( .A(oc8051_sfr1_oc8051_int1_n15), .Y(oc8051_sfr1_oc8051_int1_n14) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u40 ( .A(
        oc8051_sfr1_oc8051_int1_n45), .B(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_int1_n40) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u39 ( .A(descy), .B(
        oc8051_sfr1_oc8051_int1_n40), .Y(oc8051_sfr1_oc8051_int1_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u38 ( .A(oc8051_sfr1_oc8051_int1_n17), .Y(oc8051_sfr1_oc8051_int1_n25) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u37 ( .A0(wr_dat[0]), .A1(
        oc8051_sfr1_oc8051_int1_n14), .B0(oc8051_sfr1_oc8051_int1_n25), .Y(
        oc8051_sfr1_oc8051_int1_n42) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u36 ( .A(oc8051_sfr1_ip_0_), .Y(
        oc8051_sfr1_oc8051_int1_n43) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u35 ( .AN(
        oc8051_sfr1_oc8051_int1_n40), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n20) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u34 ( .A0(
        oc8051_sfr1_oc8051_int1_n39), .A1(oc8051_sfr1_oc8051_int1_n20), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n44) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u33 ( .A(
        oc8051_sfr1_oc8051_int1_n42), .B(oc8051_sfr1_oc8051_int1_n43), .S0(
        oc8051_sfr1_oc8051_int1_n44), .Y(oc8051_sfr1_oc8051_int1_n258) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u32 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_int1_n14), .B0(oc8051_sfr1_oc8051_int1_n25), .Y(
        oc8051_sfr1_oc8051_int1_n36) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u31 ( .A(oc8051_sfr1_ip_1_), .Y(
        oc8051_sfr1_oc8051_int1_n37) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u30 ( .AN(
        oc8051_sfr1_oc8051_int1_n40), .B(oc8051_sfr1_oc8051_int1_n41), .Y(
        oc8051_sfr1_oc8051_int1_n12) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u29 ( .A0(
        oc8051_sfr1_oc8051_int1_n39), .A1(oc8051_sfr1_oc8051_int1_n12), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n38) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u28 ( .A(
        oc8051_sfr1_oc8051_int1_n36), .B(oc8051_sfr1_oc8051_int1_n37), .S0(
        oc8051_sfr1_oc8051_int1_n38), .Y(oc8051_sfr1_oc8051_int1_n259) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u27 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_int1_n14), .B0(oc8051_sfr1_oc8051_int1_n25), .Y(
        oc8051_sfr1_oc8051_int1_n33) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u26 ( .A(oc8051_sfr1_ip_2_), .Y(
        oc8051_sfr1_oc8051_int1_n34) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u25 ( .A0(
        oc8051_sfr1_oc8051_int1_n32), .A1(oc8051_sfr1_oc8051_int1_n20), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n35) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u24 ( .A(
        oc8051_sfr1_oc8051_int1_n33), .B(oc8051_sfr1_oc8051_int1_n34), .S0(
        oc8051_sfr1_oc8051_int1_n35), .Y(oc8051_sfr1_oc8051_int1_n260) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u23 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_int1_n14), .B0(oc8051_sfr1_oc8051_int1_n25), .Y(
        oc8051_sfr1_oc8051_int1_n29) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u22 ( .A0(
        oc8051_sfr1_oc8051_int1_n32), .A1(oc8051_sfr1_oc8051_int1_n12), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n31) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u21 ( .A(
        oc8051_sfr1_oc8051_int1_n29), .B(oc8051_sfr1_oc8051_int1_n30), .S0(
        oc8051_sfr1_oc8051_int1_n31), .Y(oc8051_sfr1_oc8051_int1_n261) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u20 ( .A0(wr_dat[4]), .A1(
        oc8051_sfr1_oc8051_int1_n14), .B0(oc8051_sfr1_oc8051_int1_n25), .Y(
        oc8051_sfr1_oc8051_int1_n26) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u19 ( .A(oc8051_sfr1_ip_4_), .Y(
        oc8051_sfr1_oc8051_int1_n27) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u18 ( .A0(
        oc8051_sfr1_oc8051_int1_n24), .A1(oc8051_sfr1_oc8051_int1_n20), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n28) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u17 ( .A(
        oc8051_sfr1_oc8051_int1_n26), .B(oc8051_sfr1_oc8051_int1_n27), .S0(
        oc8051_sfr1_oc8051_int1_n28), .Y(oc8051_sfr1_oc8051_int1_n262) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u16 ( .A0(wr_dat[5]), .A1(
        oc8051_sfr1_oc8051_int1_n14), .B0(oc8051_sfr1_oc8051_int1_n25), .Y(
        oc8051_sfr1_oc8051_int1_n22) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u15 ( .A0(
        oc8051_sfr1_oc8051_int1_n24), .A1(oc8051_sfr1_oc8051_int1_n12), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n23) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u14 ( .A(
        oc8051_sfr1_oc8051_int1_n22), .B(oc8051_sfr1_oc8051_int1_n11), .S0(
        oc8051_sfr1_oc8051_int1_n23), .Y(oc8051_sfr1_oc8051_int1_n263) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u13 ( .A0(
        oc8051_sfr1_oc8051_int1_n15), .A1(oc8051_sfr1_oc8051_int1_n21), .B0(
        oc8051_sfr1_oc8051_int1_n17), .Y(oc8051_sfr1_oc8051_int1_n18) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u12 ( .A0(
        oc8051_sfr1_oc8051_int1_n20), .A1(oc8051_sfr1_oc8051_int1_n13), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n19) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u11 ( .A(
        oc8051_sfr1_oc8051_int1_n18), .B(oc8051_sfr1_ip_6_), .S0(
        oc8051_sfr1_oc8051_int1_n19), .Y(oc8051_sfr1_oc8051_int1_n264) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u10 ( .A0(
        oc8051_sfr1_oc8051_int1_n15), .A1(oc8051_sfr1_oc8051_int1_n16), .B0(
        oc8051_sfr1_oc8051_int1_n17), .Y(oc8051_sfr1_oc8051_int1_n2) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u9 ( .A0(
        oc8051_sfr1_oc8051_int1_n12), .A1(oc8051_sfr1_oc8051_int1_n13), .B0(
        oc8051_sfr1_oc8051_int1_n14), .Y(oc8051_sfr1_oc8051_int1_n3) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u8 ( .A(oc8051_sfr1_oc8051_int1_n2), 
        .B(oc8051_sfr1_ip_7_), .S0(oc8051_sfr1_oc8051_int1_n3), .Y(
        oc8051_sfr1_oc8051_int1_n265) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u7 ( .A(oc8051_sfr1_oc8051_int1_n4), 
        .Y(int_src[0]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u6 ( .A(oc8051_sfr1_oc8051_int1_n5), 
        .Y(int_src[1]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u5 ( .A(oc8051_sfr1_oc8051_int1_n6), 
        .Y(int_src[3]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u4 ( .A(oc8051_sfr1_oc8051_int1_n11), 
        .Y(oc8051_sfr1_ip_5_) );
  TIELO_X1M_A12TS oc8051_sfr1_oc8051_int1_u3 ( .Y(
        oc8051_sfr1_oc8051_int1_int_vec_2_) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_5_ ( .D(
        oc8051_sfr1_oc8051_int1_n263), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n11) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n236), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n4) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n234), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n6) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n235), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n5) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_0__2_ ( .D(
        oc8051_sfr1_oc8051_int1_n229), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n9) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_1__2_ ( .D(
        oc8051_sfr1_oc8051_int1_n226), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n10) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_4_ ( .D(
        oc8051_sfr1_oc8051_int1_n233), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n7) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_5_ ( .D(
        oc8051_sfr1_oc8051_int1_n232), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n8) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_dept_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n239), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_dept_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_4_ ( .D(
        oc8051_sfr1_oc8051_int1_n254), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_2_ ( .D(
        oc8051_sfr1_oc8051_int1_n252), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_ie1_reg ( .D(
        oc8051_sfr1_oc8051_int1_n240), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_2_ ( .D(
        oc8051_sfr1_oc8051_int1_n260), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n247), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n246), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n249), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tr1) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_ie0_reg ( .D(
        oc8051_sfr1_oc8051_int1_n241), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n250), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n259), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n258), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_4_ ( .D(
        oc8051_sfr1_oc8051_int1_n262), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n251), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n253), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_7_ ( .D(
        oc8051_sfr1_oc8051_int1_n257), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_proc_reg ( .D(
        oc8051_sfr1_oc8051_int1_n243), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_proc) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_tf0_reg ( .D(
        oc8051_sfr1_oc8051_int1_n242), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_tf1_reg ( .D(
        oc8051_sfr1_oc8051_int1_n245), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_dept_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n244), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_dept_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_2_ ( .D(
        oc8051_sfr1_oc8051_int1_n248), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tr0) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_5_ ( .D(
        oc8051_sfr1_oc8051_int1_n255), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n261), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_6_ ( .D(
        oc8051_sfr1_oc8051_int1_n264), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_6_ ( .D(
        oc8051_sfr1_oc8051_int1_n256), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_7_ ( .D(
        oc8051_sfr1_oc8051_int1_n265), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_0__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n231), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_isrc_0__0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_0__1_ ( .D(
        oc8051_sfr1_oc8051_int1_n230), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_isrc_0__1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_1__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n228), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_isrc_1__0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_1__1_ ( .D(
        oc8051_sfr1_oc8051_int1_n227), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_isrc_1__1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_lev_reg_0__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n238), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_lev_0__0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_lev_reg_1__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n237), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_lev_1__0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tf1_buff_reg ( .D(oc8051_sfr1_tf1), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_tf1_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tf0_buff_reg ( .D(oc8051_sfr1_tf0), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_tf0_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie1_buff_reg ( .D(int1_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_ie1_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie0_buff_reg ( .D(int0_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_ie0_buff) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u245 ( .A(oc8051_sfr1_tmod[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u244 ( .A(oc8051_sfr1_tmod[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n79) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u243 ( .A(
        oc8051_sfr1_oc8051_tc1_n159), .B(oc8051_sfr1_oc8051_tc1_n79), .Y(
        oc8051_sfr1_oc8051_tc1_n20) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u242 ( .A(oc8051_sfr1_pres_ow), .B(
        oc8051_sfr1_oc8051_tc1_n20), .C(oc8051_sfr1_tr1), .Y(
        oc8051_sfr1_oc8051_tc1_n16) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u241 ( .A(oc8051_sfr1_tmod[0]), .B(
        oc8051_sfr1_tmod[1]), .Y(oc8051_sfr1_oc8051_tc1_n28) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u240 ( .A(oc8051_sfr1_tmod[3]), .B(
        int0_i), .Y(oc8051_sfr1_oc8051_tc1_n162) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u239 ( .A(oc8051_sfr1_pres_ow), .Y(
        oc8051_sfr1_oc8051_tc1_n154) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u238 ( .AN(t0_i), .B(
        oc8051_sfr1_oc8051_tc1_t0_buff), .Y(oc8051_sfr1_oc8051_tc1_n164) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u237 ( .A(
        oc8051_sfr1_oc8051_tc1_n154), .B(oc8051_sfr1_oc8051_tc1_n164), .S0(
        oc8051_sfr1_tmod[2]), .Y(oc8051_sfr1_oc8051_tc1_n163) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u236 ( .A(oc8051_sfr1_tr0), .B(
        oc8051_sfr1_oc8051_tc1_n162), .C(oc8051_sfr1_oc8051_tc1_n163), .Y(
        oc8051_sfr1_oc8051_tc1_n75) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u235 ( .A(oc8051_sfr1_oc8051_tc1_n75), 
        .Y(oc8051_sfr1_oc8051_tc1_n69) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u234 ( .A(
        oc8051_sfr1_oc8051_tc1_n28), .B(oc8051_sfr1_oc8051_tc1_n69), .Y(
        oc8051_sfr1_oc8051_tc1_n161) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u233 ( .A(
        oc8051_sfr1_oc8051_tc1_n159), .B(oc8051_sfr1_tmod[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n27) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u232 ( .A(
        oc8051_sfr1_oc8051_tc1_n27), .B(oc8051_sfr1_oc8051_tc1_n69), .Y(
        oc8051_sfr1_oc8051_tc1_n66) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u231 ( .A(
        oc8051_sfr1_oc8051_tc1_n161), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_n42) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u230 ( .A(oc8051_sfr1_tl0[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n43) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u229 ( .A0(
        oc8051_sfr1_oc8051_tc1_n223), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n43), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_0) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u228 ( .A(oc8051_sfr1_tl0[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n49) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u227 ( .A0(
        oc8051_sfr1_oc8051_tc1_n222), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n49), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_1) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u226 ( .A0(
        oc8051_sfr1_oc8051_tc1_n218), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n221), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_10) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u225 ( .A0(
        oc8051_sfr1_oc8051_tc1_n217), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n220), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_11) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u224 ( .A0(
        oc8051_sfr1_oc8051_tc1_n216), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n219), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_12) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u223 ( .A(
        oc8051_sfr1_oc8051_tc1_n218), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_13) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u222 ( .A(
        oc8051_sfr1_oc8051_tc1_n217), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_14) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u221 ( .A(
        oc8051_sfr1_oc8051_tc1_n216), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_15) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u220 ( .A(oc8051_sfr1_tl0[2]), .Y(
        oc8051_sfr1_oc8051_tc1_n52) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u219 ( .A0(
        oc8051_sfr1_oc8051_tc1_n221), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n52), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_2) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u218 ( .A(oc8051_sfr1_tl0[3]), .Y(
        oc8051_sfr1_oc8051_tc1_n55) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u217 ( .A0(
        oc8051_sfr1_oc8051_tc1_n220), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n55), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_3) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u216 ( .A(oc8051_sfr1_tl0[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n58) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u215 ( .A0(
        oc8051_sfr1_oc8051_tc1_n219), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n58), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_4) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u214 ( .A(oc8051_sfr1_tl0[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n61) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u213 ( .A0(
        oc8051_sfr1_oc8051_tc1_n223), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n61), .B1(oc8051_sfr1_oc8051_tc1_n66), .C0(
        oc8051_sfr1_oc8051_tc1_n218), .C1(oc8051_sfr1_oc8051_tc1_n16), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_5) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u212 ( .A(oc8051_sfr1_tl0[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n64) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u211 ( .A0(
        oc8051_sfr1_oc8051_tc1_n222), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n64), .B1(oc8051_sfr1_oc8051_tc1_n66), .C0(
        oc8051_sfr1_oc8051_tc1_n217), .C1(oc8051_sfr1_oc8051_tc1_n16), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_6) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u210 ( .A(oc8051_sfr1_tl0[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n1) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u209 ( .A0(
        oc8051_sfr1_oc8051_tc1_n221), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n1), .B1(oc8051_sfr1_oc8051_tc1_n66), .C0(
        oc8051_sfr1_oc8051_tc1_n216), .C1(oc8051_sfr1_oc8051_tc1_n16), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_7) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u208 ( .A0(
        oc8051_sfr1_oc8051_tc1_n220), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n223), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_8) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u207 ( .A0(
        oc8051_sfr1_oc8051_tc1_n219), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n222), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_9) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u206 ( .A(oc8051_sfr1_th1[5]), .B(
        oc8051_sfr1_th1[2]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_10) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u205 ( .A(oc8051_sfr1_th1[6]), .B(
        oc8051_sfr1_th1[3]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_11) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u204 ( .A(oc8051_sfr1_th1[7]), .B(
        oc8051_sfr1_th1[4]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_12) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u203 ( .A(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n120) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u202 ( .A(oc8051_sfr1_th1[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n140) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u201 ( .A(
        oc8051_sfr1_oc8051_tc1_n120), .B(oc8051_sfr1_oc8051_tc1_n140), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_13) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u200 ( .A(oc8051_sfr1_th1[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n113) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u199 ( .A(
        oc8051_sfr1_oc8051_tc1_n120), .B(oc8051_sfr1_oc8051_tc1_n113), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_14) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u198 ( .A(oc8051_sfr1_th1[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n87) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u197 ( .A(oc8051_sfr1_oc8051_tc1_n87), .B(oc8051_sfr1_oc8051_tc1_n120), .Y(oc8051_sfr1_oc8051_tc1_u3_u8_z_15) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u196 ( .A(oc8051_sfr1_th1[0]), .B(
        oc8051_sfr1_tl1[5]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_5) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u195 ( .A(oc8051_sfr1_th1[1]), .B(
        oc8051_sfr1_tl1[6]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_6) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u194 ( .A(oc8051_sfr1_th1[2]), .B(
        oc8051_sfr1_tl1[7]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_7) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u193 ( .A(oc8051_sfr1_th1[3]), .B(
        oc8051_sfr1_th1[0]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_8) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u192 ( .A(oc8051_sfr1_th1[4]), .B(
        oc8051_sfr1_th1[1]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_9) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u191 ( .A(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n26) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u190 ( .AN(n_5_net_), .B(
        oc8051_sfr1_wr_bit_r), .Y(oc8051_sfr1_oc8051_tc1_n157) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u189 ( .A(wr_addr[4]), .B(wr_addr[6]), .C(wr_addr[5]), .Y(oc8051_sfr1_oc8051_tc1_n160) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u188 ( .A(wr_addr[7]), .B(wr_addr[3]), .C(oc8051_sfr1_oc8051_tc1_n160), .Y(oc8051_sfr1_oc8051_tc1_n156) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u187 ( .AN(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_tc1_n157), .C(oc8051_sfr1_oc8051_tc1_n156), .Y(
        oc8051_sfr1_oc8051_tc1_n80) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u186 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n83) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u185 ( .A(oc8051_sfr1_oc8051_tc1_n80), .B(wr_addr[1]), .C(oc8051_sfr1_oc8051_tc1_n83), .Y(
        oc8051_sfr1_oc8051_tc1_n158) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u184 ( .A(
        oc8051_sfr1_oc8051_tc1_n159), .B(oc8051_sfr1_oc8051_tc1_n26), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n224) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u183 ( .A(wr_dat[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n30) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u182 ( .A(
        oc8051_sfr1_oc8051_tc1_n79), .B(oc8051_sfr1_oc8051_tc1_n30), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n225) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u181 ( .A(oc8051_sfr1_tmod[2]), .B(
        wr_dat[2]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n226) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u180 ( .A(oc8051_sfr1_tmod[3]), .B(
        wr_dat[3]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n227) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u179 ( .A(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n36) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u178 ( .A(
        oc8051_sfr1_oc8051_tc1_n120), .B(oc8051_sfr1_oc8051_tc1_n36), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n228) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u177 ( .A(oc8051_sfr1_tmod[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n92) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u176 ( .A(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n38) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u175 ( .A(
        oc8051_sfr1_oc8051_tc1_n92), .B(oc8051_sfr1_oc8051_tc1_n38), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n229) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u174 ( .A(oc8051_sfr1_tmod[6]), .B(
        wr_dat[6]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n230) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u173 ( .A(oc8051_sfr1_tmod[7]), .B(
        wr_dat[7]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n231) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u172 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n81) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u171 ( .A(oc8051_sfr1_oc8051_tc1_n81), .B(oc8051_sfr1_oc8051_tc1_n80), .C(oc8051_sfr1_oc8051_tc1_n83), .Y(
        oc8051_sfr1_oc8051_tc1_n90) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u170 ( .A(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_tc1_n156), .C(oc8051_sfr1_oc8051_tc1_n157), .D(
        oc8051_sfr1_oc8051_tc1_n81), .Y(oc8051_sfr1_oc8051_tc1_n82) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u169 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_tc1_n82), .Y(oc8051_sfr1_oc8051_tc1_n114) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u168 ( .A(oc8051_sfr1_oc8051_tc1_n114), .Y(oc8051_sfr1_oc8051_tc1_n99) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u167 ( .A(oc8051_sfr1_oc8051_tc1_n90), .B(oc8051_sfr1_oc8051_tc1_n99), .Y(oc8051_sfr1_oc8051_tc1_n119) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u166 ( .A(oc8051_sfr1_oc8051_tc1_n90), 
        .Y(oc8051_sfr1_oc8051_tc1_n125) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u165 ( .AN(t1_i), .B(
        oc8051_sfr1_oc8051_tc1_t1_buff), .Y(oc8051_sfr1_oc8051_tc1_n155) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u164 ( .A(
        oc8051_sfr1_oc8051_tc1_n154), .B(oc8051_sfr1_oc8051_tc1_n155), .S0(
        oc8051_sfr1_tmod[6]), .Y(oc8051_sfr1_oc8051_tc1_n152) );
  AOI21B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u163 ( .A0(oc8051_sfr1_tmod[7]), 
        .A1(int1_i), .B0N(oc8051_sfr1_tr1), .Y(oc8051_sfr1_oc8051_tc1_n153) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u162 ( .A(
        oc8051_sfr1_oc8051_tc1_n152), .B(oc8051_sfr1_oc8051_tc1_n119), .C(
        oc8051_sfr1_oc8051_tc1_n153), .Y(oc8051_sfr1_oc8051_tc1_n122) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u161 ( .A(
        oc8051_sfr1_oc8051_tc1_n125), .B(oc8051_sfr1_oc8051_tc1_n122), .Y(
        oc8051_sfr1_oc8051_tc1_n124) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u160 ( .A(
        oc8051_sfr1_oc8051_tc1_n119), .B(oc8051_sfr1_oc8051_tc1_n124), .Y(
        oc8051_sfr1_oc8051_tc1_n138) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u159 ( .A(oc8051_sfr1_oc8051_tc1_n174), .Y(oc8051_sfr1_oc8051_tc1_n110) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u158 ( .A(oc8051_sfr1_tmod[5]), .B(
        oc8051_sfr1_oc8051_tc1_n110), .Y(oc8051_sfr1_oc8051_tc1_n151) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u157 ( .A(
        oc8051_sfr1_oc8051_tc1_n192), .B(oc8051_sfr1_oc8051_tc1_n151), .S0(
        oc8051_sfr1_oc8051_tc1_n120), .Y(oc8051_sfr1_oc8051_tc1_n146) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u156 ( .A(
        oc8051_sfr1_oc8051_tc1_n233), .B(oc8051_sfr1_oc8051_tc1_n99), .Y(
        oc8051_sfr1_oc8051_tc1_n148) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u155 ( .A(oc8051_sfr1_tl1[3]), .B(
        oc8051_sfr1_tl1[2]), .C(oc8051_sfr1_tl1[1]), .D(oc8051_sfr1_tl1[0]), 
        .Y(oc8051_sfr1_oc8051_tc1_n149) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u154 ( .A(oc8051_sfr1_tl1[7]), .B(
        oc8051_sfr1_tl1[6]), .C(oc8051_sfr1_tl1[5]), .D(oc8051_sfr1_tl1[4]), 
        .Y(oc8051_sfr1_oc8051_tc1_n150) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u153 ( .A(
        oc8051_sfr1_oc8051_tc1_n149), .B(oc8051_sfr1_oc8051_tc1_n150), .Y(
        oc8051_sfr1_oc8051_tc1_n145) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u152 ( .A(oc8051_sfr1_tmod[5]), .B(
        oc8051_sfr1_oc8051_tc1_n119), .C(oc8051_sfr1_oc8051_tc1_n145), .Y(
        oc8051_sfr1_oc8051_tc1_n86) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u151 ( .A(oc8051_sfr1_oc8051_tc1_n86), 
        .Y(oc8051_sfr1_oc8051_tc1_n127) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u150 ( .A(
        oc8051_sfr1_oc8051_tc1_n148), .B(oc8051_sfr1_oc8051_tc1_n127), .S0(
        oc8051_sfr1_oc8051_tc1_n124), .Y(oc8051_sfr1_oc8051_tc1_n147) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u149 ( .A0(
        oc8051_sfr1_oc8051_tc1_n138), .A1(oc8051_sfr1_oc8051_tc1_n146), .B0(
        oc8051_sfr1_oc8051_tc1_n147), .Y(oc8051_sfr1_oc8051_tc1_n234) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u148 ( .A(oc8051_sfr1_oc8051_tc1_n92), .B(oc8051_sfr1_oc8051_tc1_n145), .Y(oc8051_sfr1_oc8051_tc1_n91) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u147 ( .A0(
        oc8051_sfr1_oc8051_tc1_n202), .A1(oc8051_sfr1_oc8051_tc1_n91), .B0(
        oc8051_sfr1_oc8051_tc1_n167), .B1(oc8051_sfr1_oc8051_tc1_n92), .Y(
        oc8051_sfr1_oc8051_tc1_n142) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u146 ( .A0(
        oc8051_sfr1_oc8051_tc1_n92), .A1(oc8051_sfr1_oc8051_tc1_n120), .B0(
        oc8051_sfr1_oc8051_tc1_n122), .C0(oc8051_sfr1_oc8051_tc1_n125), .Y(
        oc8051_sfr1_oc8051_tc1_n144) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u145 ( .A(
        oc8051_sfr1_oc8051_tc1_n119), .B(oc8051_sfr1_oc8051_tc1_n144), .Y(
        oc8051_sfr1_oc8051_tc1_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u144 ( .A(oc8051_sfr1_oc8051_tc1_n144), .Y(oc8051_sfr1_oc8051_tc1_n89) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u143 ( .A0(
        oc8051_sfr1_oc8051_tc1_n89), .A1(oc8051_sfr1_tl1[6]), .B0(
        oc8051_sfr1_oc8051_tc1_n90), .B1(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n143) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u142 ( .A0(
        oc8051_sfr1_oc8051_tc1_n142), .A1(oc8051_sfr1_oc8051_tc1_n85), .B0(
        oc8051_sfr1_oc8051_tc1_n86), .B1(oc8051_sfr1_oc8051_tc1_n113), .C0(
        oc8051_sfr1_oc8051_tc1_n143), .Y(oc8051_sfr1_oc8051_tc1_n235) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u141 ( .A0(
        oc8051_sfr1_oc8051_tc1_n201), .A1(oc8051_sfr1_oc8051_tc1_n91), .B0(
        oc8051_sfr1_oc8051_tc1_n166), .B1(oc8051_sfr1_oc8051_tc1_n92), .Y(
        oc8051_sfr1_oc8051_tc1_n139) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u140 ( .A0(
        oc8051_sfr1_oc8051_tc1_n89), .A1(oc8051_sfr1_tl1[5]), .B0(
        oc8051_sfr1_oc8051_tc1_n90), .B1(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n141) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u139 ( .A0(
        oc8051_sfr1_oc8051_tc1_n139), .A1(oc8051_sfr1_oc8051_tc1_n85), .B0(
        oc8051_sfr1_oc8051_tc1_n86), .B1(oc8051_sfr1_oc8051_tc1_n140), .C0(
        oc8051_sfr1_oc8051_tc1_n141), .Y(oc8051_sfr1_oc8051_tc1_n236) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u138 ( .A(oc8051_sfr1_tl1[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n136) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u137 ( .AN(
        oc8051_sfr1_oc8051_tc1_n91), .B(oc8051_sfr1_oc8051_tc1_n138), .Y(
        oc8051_sfr1_oc8051_tc1_n128) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u136 ( .A(oc8051_sfr1_oc8051_tc1_n92), .B(oc8051_sfr1_tmod[4]), .Y(oc8051_sfr1_oc8051_tc1_n121) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u135 ( .A(
        oc8051_sfr1_oc8051_tc1_n138), .B(oc8051_sfr1_oc8051_tc1_n121), .Y(
        oc8051_sfr1_oc8051_tc1_n129) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u134 ( .A0(oc8051_sfr1_th1[4]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n200), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n165), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n137) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u133 ( .A0(
        oc8051_sfr1_oc8051_tc1_n136), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n36), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n137), .Y(oc8051_sfr1_oc8051_tc1_n237) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u132 ( .A(oc8051_sfr1_tl1[3]), .Y(
        oc8051_sfr1_oc8051_tc1_n134) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u131 ( .A(wr_dat[3]), .Y(
        oc8051_sfr1_oc8051_tc1_n34) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u130 ( .A0(oc8051_sfr1_th1[3]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n199), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1640), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n135) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u129 ( .A0(
        oc8051_sfr1_oc8051_tc1_n134), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n34), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n135), .Y(oc8051_sfr1_oc8051_tc1_n238) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u128 ( .A(oc8051_sfr1_tl1[2]), .Y(
        oc8051_sfr1_oc8051_tc1_n132) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u127 ( .A(wr_dat[2]), .Y(
        oc8051_sfr1_oc8051_tc1_n32) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u126 ( .A0(oc8051_sfr1_th1[2]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n198), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1630), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n133) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u125 ( .A0(
        oc8051_sfr1_oc8051_tc1_n132), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n32), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n133), .Y(oc8051_sfr1_oc8051_tc1_n239) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u124 ( .A(oc8051_sfr1_tl1[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n130) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u123 ( .A0(oc8051_sfr1_th1[1]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n197), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1620), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n131) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u122 ( .A0(
        oc8051_sfr1_oc8051_tc1_n130), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n30), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n131), .Y(oc8051_sfr1_oc8051_tc1_n240) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u121 ( .A(oc8051_sfr1_tl1[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n123) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u120 ( .A0(oc8051_sfr1_th1[0]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n196), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1610), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n126) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u119 ( .A0(
        oc8051_sfr1_oc8051_tc1_n123), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n26), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n126), .Y(oc8051_sfr1_oc8051_tc1_n241) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u118 ( .A0(
        oc8051_sfr1_oc8051_tc1_n121), .A1(oc8051_sfr1_oc8051_tc1_n122), .B0(
        oc8051_sfr1_oc8051_tc1_n114), .Y(oc8051_sfr1_oc8051_tc1_n112) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u117 ( .A(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n9) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u116 ( .A(
        oc8051_sfr1_oc8051_tc1_n112), .B(oc8051_sfr1_oc8051_tc1_n120), .C(
        oc8051_sfr1_oc8051_tc1_n119), .Y(oc8051_sfr1_oc8051_tc1_n93) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u115 ( .A(oc8051_sfr1_oc8051_tc1_n93), 
        .Y(oc8051_sfr1_oc8051_tc1_n116) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u114 ( .A(
        oc8051_sfr1_oc8051_tc1_n119), .B(oc8051_sfr1_oc8051_tc1_n112), .C(
        oc8051_sfr1_tmod[4]), .Y(oc8051_sfr1_oc8051_tc1_n95) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u113 ( .A(oc8051_sfr1_oc8051_tc1_n95), 
        .Y(oc8051_sfr1_oc8051_tc1_n117) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u112 ( .A0(
        oc8051_sfr1_oc8051_tc1_n173), .A1(oc8051_sfr1_oc8051_tc1_n116), .B0(
        oc8051_sfr1_oc8051_tc1_n191), .B1(oc8051_sfr1_oc8051_tc1_n117), .Y(
        oc8051_sfr1_oc8051_tc1_n118) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u111 ( .A0(
        oc8051_sfr1_oc8051_tc1_n87), .A1(oc8051_sfr1_oc8051_tc1_n112), .B0(
        oc8051_sfr1_oc8051_tc1_n9), .B1(oc8051_sfr1_oc8051_tc1_n114), .C0(
        oc8051_sfr1_oc8051_tc1_n118), .Y(oc8051_sfr1_oc8051_tc1_n242) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u110 ( .A(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n40) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u109 ( .A0(
        oc8051_sfr1_oc8051_tc1_n172), .A1(oc8051_sfr1_oc8051_tc1_n116), .B0(
        oc8051_sfr1_oc8051_tc1_n190), .B1(oc8051_sfr1_oc8051_tc1_n117), .Y(
        oc8051_sfr1_oc8051_tc1_n115) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u108 ( .A0(
        oc8051_sfr1_oc8051_tc1_n112), .A1(oc8051_sfr1_oc8051_tc1_n113), .B0(
        oc8051_sfr1_oc8051_tc1_n40), .B1(oc8051_sfr1_oc8051_tc1_n114), .C0(
        oc8051_sfr1_oc8051_tc1_n115), .Y(oc8051_sfr1_oc8051_tc1_n243) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u107 ( .A(oc8051_sfr1_oc8051_tc1_n171), .Y(oc8051_sfr1_oc8051_tc1_n104) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u106 ( .A(oc8051_sfr1_oc8051_tc1_n112), .Y(oc8051_sfr1_oc8051_tc1_n98) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u105 ( .A0(oc8051_sfr1_th1[5]), 
        .A1(oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[5]), .Y(oc8051_sfr1_oc8051_tc1_n111) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u104 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n104), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n110), .C0(
        oc8051_sfr1_oc8051_tc1_n111), .Y(oc8051_sfr1_oc8051_tc1_n244) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u103 ( .A(oc8051_sfr1_oc8051_tc1_n170), .Y(oc8051_sfr1_oc8051_tc1_n101) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u102 ( .A(oc8051_sfr1_oc8051_tc1_n173), .Y(oc8051_sfr1_oc8051_tc1_n108) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u101 ( .A0(oc8051_sfr1_th1[4]), 
        .A1(oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[4]), .Y(oc8051_sfr1_oc8051_tc1_n109) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u100 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n101), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n108), .C0(
        oc8051_sfr1_oc8051_tc1_n109), .Y(oc8051_sfr1_oc8051_tc1_n245) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u99 ( .A(oc8051_sfr1_oc8051_tc1_n169), 
        .Y(oc8051_sfr1_oc8051_tc1_n96) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u98 ( .A(oc8051_sfr1_oc8051_tc1_n172), 
        .Y(oc8051_sfr1_oc8051_tc1_n106) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u97 ( .A0(oc8051_sfr1_th1[3]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[3]), .Y(oc8051_sfr1_oc8051_tc1_n107) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u96 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n96), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n106), .C0(
        oc8051_sfr1_oc8051_tc1_n107), .Y(oc8051_sfr1_oc8051_tc1_n246) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u95 ( .A(oc8051_sfr1_oc8051_tc1_n168), 
        .Y(oc8051_sfr1_oc8051_tc1_n103) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u94 ( .A0(oc8051_sfr1_th1[2]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[2]), .Y(oc8051_sfr1_oc8051_tc1_n105) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u93 ( .A0(
        oc8051_sfr1_oc8051_tc1_n103), .A1(oc8051_sfr1_oc8051_tc1_n93), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n104), .C0(
        oc8051_sfr1_oc8051_tc1_n105), .Y(oc8051_sfr1_oc8051_tc1_n247) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u92 ( .A(oc8051_sfr1_oc8051_tc1_n167), 
        .Y(oc8051_sfr1_oc8051_tc1_n100) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u91 ( .A0(oc8051_sfr1_th1[1]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[1]), .Y(oc8051_sfr1_oc8051_tc1_n102) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u90 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n100), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n101), .C0(
        oc8051_sfr1_oc8051_tc1_n102), .Y(oc8051_sfr1_oc8051_tc1_n248) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u89 ( .A(oc8051_sfr1_oc8051_tc1_n166), 
        .Y(oc8051_sfr1_oc8051_tc1_n94) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u88 ( .A0(oc8051_sfr1_th1[0]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[0]), .Y(oc8051_sfr1_oc8051_tc1_n97) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u87 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n94), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n96), .C0(
        oc8051_sfr1_oc8051_tc1_n97), .Y(oc8051_sfr1_oc8051_tc1_n249) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u86 ( .A0(
        oc8051_sfr1_oc8051_tc1_n203), .A1(oc8051_sfr1_oc8051_tc1_n91), .B0(
        oc8051_sfr1_oc8051_tc1_n168), .B1(oc8051_sfr1_oc8051_tc1_n92), .Y(
        oc8051_sfr1_oc8051_tc1_n84) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u85 ( .A0(
        oc8051_sfr1_oc8051_tc1_n89), .A1(oc8051_sfr1_tl1[7]), .B0(
        oc8051_sfr1_oc8051_tc1_n90), .B1(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n88) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u84 ( .A0(
        oc8051_sfr1_oc8051_tc1_n84), .A1(oc8051_sfr1_oc8051_tc1_n85), .B0(
        oc8051_sfr1_oc8051_tc1_n86), .B1(oc8051_sfr1_oc8051_tc1_n87), .C0(
        oc8051_sfr1_oc8051_tc1_n88), .Y(oc8051_sfr1_oc8051_tc1_n250) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u83 ( .A0(
        oc8051_sfr1_oc8051_tc1_n920), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n630), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n600), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n76) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u82 ( .A(oc8051_sfr1_oc8051_tc1_n82), .B(oc8051_sfr1_oc8051_tc1_n83), .Y(oc8051_sfr1_oc8051_tc1_n25) );
  OR3_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u81 ( .A(oc8051_sfr1_oc8051_tc1_n80), 
        .B(wr_addr[0]), .C(oc8051_sfr1_oc8051_tc1_n81), .Y(
        oc8051_sfr1_oc8051_tc1_n8) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u80 ( .A(oc8051_sfr1_oc8051_tc1_n25), .B(oc8051_sfr1_oc8051_tc1_n8), .Y(oc8051_sfr1_oc8051_tc1_n15) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u79 ( .A(oc8051_sfr1_oc8051_tc1_n79), 
        .B(oc8051_sfr1_tmod[0]), .Y(oc8051_sfr1_oc8051_tc1_n68) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u78 ( .A(oc8051_sfr1_oc8051_tc1_n15), 
        .Y(oc8051_sfr1_oc8051_tc1_n21) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u77 ( .A(oc8051_sfr1_tl0[3]), .B(
        oc8051_sfr1_tl0[2]), .C(oc8051_sfr1_tl0[1]), .D(oc8051_sfr1_tl0[0]), 
        .Y(oc8051_sfr1_oc8051_tc1_n77) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u76 ( .A(oc8051_sfr1_tl0[7]), .B(
        oc8051_sfr1_tl0[6]), .C(oc8051_sfr1_tl0[5]), .D(oc8051_sfr1_tl0[4]), 
        .Y(oc8051_sfr1_oc8051_tc1_n78) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u75 ( .A(oc8051_sfr1_oc8051_tc1_n77), 
        .B(oc8051_sfr1_oc8051_tc1_n78), .Y(oc8051_sfr1_oc8051_tc1_n71) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u74 ( .A(oc8051_sfr1_oc8051_tc1_n68), .B(oc8051_sfr1_oc8051_tc1_n21), .C(oc8051_sfr1_oc8051_tc1_n71), .Y(
        oc8051_sfr1_oc8051_tc1_n10) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u73 ( .A0(
        oc8051_sfr1_oc8051_tc1_n76), .A1(oc8051_sfr1_oc8051_tc1_n15), .B0(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n73) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u72 ( .A0(
        oc8051_sfr1_oc8051_tc1_n75), .A1(oc8051_sfr1_oc8051_tc1_n15), .B0(
        oc8051_sfr1_oc8051_tc1_n8), .Y(oc8051_sfr1_oc8051_tc1_n45) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u71 ( .AN(
        oc8051_sfr1_oc8051_tc1_n25), .B(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n74) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u70 ( .A(oc8051_sfr1_oc8051_tc1_n73), 
        .B(oc8051_sfr1_tf0), .S0(oc8051_sfr1_oc8051_tc1_n74), .Y(
        oc8051_sfr1_oc8051_tc1_n251) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u69 ( .A(oc8051_sfr1_oc8051_tc1_n27), 
        .Y(oc8051_sfr1_oc8051_tc1_n18) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u68 ( .A(oc8051_sfr1_oc8051_tc1_n15), 
        .B(oc8051_sfr1_oc8051_tc1_n18), .Y(oc8051_sfr1_oc8051_tc1_n4) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u67 ( .A(oc8051_sfr1_oc8051_tc1_n68), 
        .Y(oc8051_sfr1_oc8051_tc1_n19) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u66 ( .A(oc8051_sfr1_oc8051_tc1_n20), 
        .Y(oc8051_sfr1_oc8051_tc1_n72) );
  OA21A1OI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u65 ( .A0(
        oc8051_sfr1_oc8051_tc1_n19), .A1(oc8051_sfr1_oc8051_tc1_n71), .B0(
        oc8051_sfr1_oc8051_tc1_n72), .C0(oc8051_sfr1_oc8051_tc1_n15), .Y(
        oc8051_sfr1_oc8051_tc1_n6) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u64 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n40), .B0(oc8051_sfr1_oc8051_tc1_n217), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n70) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u63 ( .A0(
        oc8051_sfr1_oc8051_tc1_n530), .A1(oc8051_sfr1_oc8051_tc1_n4), .B0(
        oc8051_sfr1_oc8051_tc1_n900), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n70), .Y(oc8051_sfr1_oc8051_tc1_n65) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u62 ( .A0(
        oc8051_sfr1_oc8051_tc1_n68), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n69), .Y(oc8051_sfr1_oc8051_tc1_n67) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u61 ( .A0(
        oc8051_sfr1_oc8051_tc1_n66), .A1(oc8051_sfr1_oc8051_tc1_n67), .B0(
        oc8051_sfr1_oc8051_tc1_n15), .C0(oc8051_sfr1_oc8051_tc1_n8), .Y(
        oc8051_sfr1_oc8051_tc1_n3) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u60 ( .A(oc8051_sfr1_oc8051_tc1_n64), .B(oc8051_sfr1_oc8051_tc1_n65), .S0(oc8051_sfr1_oc8051_tc1_n3), .Y(
        oc8051_sfr1_oc8051_tc1_n252) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u59 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n38), .B0(oc8051_sfr1_oc8051_tc1_n218), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n63) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u58 ( .A0(
        oc8051_sfr1_oc8051_tc1_n520), .A1(oc8051_sfr1_oc8051_tc1_n4), .B0(
        oc8051_sfr1_oc8051_tc1_n890), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n63), .Y(oc8051_sfr1_oc8051_tc1_n62) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u57 ( .A(oc8051_sfr1_oc8051_tc1_n61), .B(oc8051_sfr1_oc8051_tc1_n62), .S0(oc8051_sfr1_oc8051_tc1_n3), .Y(
        oc8051_sfr1_oc8051_tc1_n253) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u56 ( .A(oc8051_sfr1_oc8051_tc1_n28), 
        .Y(oc8051_sfr1_oc8051_tc1_n17) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u55 ( .A0(
        oc8051_sfr1_oc8051_tc1_n17), .A1(oc8051_sfr1_oc8051_tc1_n18), .B0(
        oc8051_sfr1_oc8051_tc1_n15), .Y(oc8051_sfr1_oc8051_tc1_n46) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u54 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n36), .B0(oc8051_sfr1_oc8051_tc1_n219), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n60) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u53 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n510), .B0(
        oc8051_sfr1_oc8051_tc1_n880), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n60), .Y(oc8051_sfr1_oc8051_tc1_n59) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u52 ( .A(oc8051_sfr1_oc8051_tc1_n58), .B(oc8051_sfr1_oc8051_tc1_n59), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n254) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u51 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n34), .B0(oc8051_sfr1_oc8051_tc1_n220), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n57) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u50 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n500), .B0(
        oc8051_sfr1_oc8051_tc1_n870), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n57), .Y(oc8051_sfr1_oc8051_tc1_n56) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u49 ( .A(oc8051_sfr1_oc8051_tc1_n55), .B(oc8051_sfr1_oc8051_tc1_n56), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n255) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u48 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n32), .B0(oc8051_sfr1_oc8051_tc1_n221), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n54) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u47 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n490), .B0(
        oc8051_sfr1_oc8051_tc1_n860), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n54), .Y(oc8051_sfr1_oc8051_tc1_n53) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u46 ( .A(oc8051_sfr1_oc8051_tc1_n52), .B(oc8051_sfr1_oc8051_tc1_n53), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n256) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u45 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n30), .B0(oc8051_sfr1_oc8051_tc1_n222), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n51) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u44 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n480), .B0(
        oc8051_sfr1_oc8051_tc1_n850), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n51), .Y(oc8051_sfr1_oc8051_tc1_n50) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u43 ( .A(oc8051_sfr1_oc8051_tc1_n49), .B(oc8051_sfr1_oc8051_tc1_n50), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n257) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u42 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_0), .Y(oc8051_sfr1_oc8051_tc1_n47) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u41 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n26), .B0(oc8051_sfr1_oc8051_tc1_n223), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n48) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u40 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n47), .B0(
        oc8051_sfr1_oc8051_tc1_n840), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n48), .Y(oc8051_sfr1_oc8051_tc1_n44) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u39 ( .A(oc8051_sfr1_oc8051_tc1_n43), .B(oc8051_sfr1_oc8051_tc1_n44), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n258) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u38 ( .A0(
        oc8051_sfr1_oc8051_tc1_n42), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n15), .C0(oc8051_sfr1_oc8051_tc1_n25), .Y(
        oc8051_sfr1_oc8051_tc1_n22) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u37 ( .A0(
        oc8051_sfr1_oc8051_tc1_n20), .A1(oc8051_sfr1_oc8051_tc1_n540), .B0(
        oc8051_sfr1_oc8051_tc1_n620), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n590), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n41) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u36 ( .A(oc8051_sfr1_oc8051_tc1_n21), .B(oc8051_sfr1_oc8051_tc1_n22), .Y(oc8051_sfr1_oc8051_tc1_n24) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u35 ( .A0(
        oc8051_sfr1_oc8051_tc1_n216), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n41), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n9), .C1(oc8051_sfr1_oc8051_tc1_n25), .Y(
        oc8051_sfr1_oc8051_tc1_n259) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u34 ( .A0(
        oc8051_sfr1_oc8051_tc1_n530), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n610), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n580), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n39) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u33 ( .A0(
        oc8051_sfr1_oc8051_tc1_n217), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n39), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n40), .Y(
        oc8051_sfr1_oc8051_tc1_n260) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u32 ( .A0(
        oc8051_sfr1_oc8051_tc1_n520), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n600), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n570), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n37) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u31 ( .A0(
        oc8051_sfr1_oc8051_tc1_n218), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n37), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n38), .Y(
        oc8051_sfr1_oc8051_tc1_n261) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u30 ( .A0(
        oc8051_sfr1_oc8051_tc1_n510), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n590), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n560), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n35) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u29 ( .A0(
        oc8051_sfr1_oc8051_tc1_n219), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n35), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n36), .Y(
        oc8051_sfr1_oc8051_tc1_n262) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u28 ( .A0(
        oc8051_sfr1_oc8051_tc1_n500), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n580), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n28), .C1(oc8051_sfr1_oc8051_tc1_n550), .Y(
        oc8051_sfr1_oc8051_tc1_n33) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u27 ( .A0(
        oc8051_sfr1_oc8051_tc1_n220), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n33), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n34), .Y(
        oc8051_sfr1_oc8051_tc1_n263) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u26 ( .A0(
        oc8051_sfr1_oc8051_tc1_n490), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n570), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n28), .C1(oc8051_sfr1_oc8051_tc1_n540), .Y(
        oc8051_sfr1_oc8051_tc1_n31) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u25 ( .A0(
        oc8051_sfr1_oc8051_tc1_n221), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n31), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n32), .Y(
        oc8051_sfr1_oc8051_tc1_n264) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u24 ( .A0(
        oc8051_sfr1_oc8051_tc1_n480), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n560), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n530), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n29) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u23 ( .A0(
        oc8051_sfr1_oc8051_tc1_n222), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n29), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n30), .Y(
        oc8051_sfr1_oc8051_tc1_n265) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u22 ( .A0(
        oc8051_sfr1_oc8051_tc1_n470), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n550), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n520), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n23) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u21 ( .A0(
        oc8051_sfr1_oc8051_tc1_n223), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n23), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n26), .Y(
        oc8051_sfr1_oc8051_tc1_n266) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u20 ( .A(oc8051_sfr1_oc8051_tc1_n20), .B(oc8051_sfr1_oc8051_tc1_n21), .C(oc8051_sfr1_oc8051_tc1_n550), .Y(
        oc8051_sfr1_oc8051_tc1_n11) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u19 ( .A(oc8051_sfr1_oc8051_tc1_n17), .B(oc8051_sfr1_oc8051_tc1_n18), .C(oc8051_sfr1_oc8051_tc1_n19), .Y(
        oc8051_sfr1_oc8051_tc1_n13) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u18 ( .A(oc8051_sfr1_oc8051_tc1_n16), 
        .Y(oc8051_sfr1_oc8051_tc1_n14) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u17 ( .A(oc8051_sfr1_oc8051_tc1_n13), 
        .B(oc8051_sfr1_oc8051_tc1_n14), .C(oc8051_sfr1_oc8051_tc1_n15), .Y(
        oc8051_sfr1_oc8051_tc1_n12) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u16 ( .A(oc8051_sfr1_oc8051_tc1_n11), .B(oc8051_sfr1_oc8051_tc1_n232), .S0(oc8051_sfr1_oc8051_tc1_n12), .Y(
        oc8051_sfr1_oc8051_tc1_n267) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u15 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n9), .B0(oc8051_sfr1_oc8051_tc1_n216), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n7) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u14 ( .A0(
        oc8051_sfr1_oc8051_tc1_n540), .A1(oc8051_sfr1_oc8051_tc1_n4), .B0(
        oc8051_sfr1_oc8051_tc1_n910), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n7), .Y(oc8051_sfr1_oc8051_tc1_n2) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u13 ( .A(oc8051_sfr1_oc8051_tc1_n1), 
        .B(oc8051_sfr1_oc8051_tc1_n2), .S0(oc8051_sfr1_oc8051_tc1_n3), .Y(
        oc8051_sfr1_oc8051_tc1_n268) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u12 ( .A(oc8051_sfr1_oc8051_tc1_n216), 
        .Y(oc8051_sfr1_th0[7]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u11 ( .A(oc8051_sfr1_oc8051_tc1_n217), 
        .Y(oc8051_sfr1_th0[6]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u10 ( .A(oc8051_sfr1_oc8051_tc1_n218), 
        .Y(oc8051_sfr1_th0[5]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u9 ( .A(oc8051_sfr1_oc8051_tc1_n219), 
        .Y(oc8051_sfr1_th0[4]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u8 ( .A(oc8051_sfr1_oc8051_tc1_n220), 
        .Y(oc8051_sfr1_th0[3]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u7 ( .A(oc8051_sfr1_oc8051_tc1_n221), 
        .Y(oc8051_sfr1_th0[2]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u6 ( .A(oc8051_sfr1_oc8051_tc1_n222), 
        .Y(oc8051_sfr1_th0[1]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u5 ( .A(oc8051_sfr1_oc8051_tc1_n223), 
        .Y(oc8051_sfr1_th0[0]) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u4 ( .A(oc8051_sfr1_oc8051_tc1_n233), .B(oc8051_sfr1_oc8051_tc1_n232), .Y(oc8051_sfr1_tf1) );
  TIELO_X1M_A12TS oc8051_sfr1_oc8051_tc1_u3 ( .Y(oc8051_sfr1_oc8051_tc1_n5) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n259), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n216) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n260), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n217) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n261), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n218) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n264), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n221) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n265), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n222) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n266), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n223) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n262), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n219) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n263), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n220) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n241), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n228), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[4]) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_tf1_0_reg ( .D(
        oc8051_sfr1_oc8051_tc1_n267), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n232) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_tf1_1_reg ( .D(
        oc8051_sfr1_oc8051_tc1_n234), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n233) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n238), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n237), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n240), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n239), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n258), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n236), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n235), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n255), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n268), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n254), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n253), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n257), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n256), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n252), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n250), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n245), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n246), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n247), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n248), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n249), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n229), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n224), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n225), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n244), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n226), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n230), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n227), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n242), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n243), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n231), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tf0_reg ( .D(
        oc8051_sfr1_oc8051_tc1_n251), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tf0) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_t1_buff_reg ( .D(t1_i), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc1_t1_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_t0_buff_reg ( .D(t0_i), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc1_t0_buff) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1 ( .A(oc8051_sfr1_tl1[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n1610) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_13 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_13), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[13]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[14]), .S(oc8051_sfr1_oc8051_tc1_n174) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_14 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_14), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[14]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[15]), .S(oc8051_sfr1_oc8051_tc1_n190) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_15 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_15), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[15]), .CO(
        oc8051_sfr1_oc8051_tc1_n192), .S(oc8051_sfr1_oc8051_tc1_n191) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_5 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_5), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[6]), .S(oc8051_sfr1_oc8051_tc1_n166)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_6 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_6), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[7]), .S(oc8051_sfr1_oc8051_tc1_n167)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_7 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_7), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[8]), .S(oc8051_sfr1_oc8051_tc1_n168)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_8 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_8), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[8]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[9]), .S(oc8051_sfr1_oc8051_tc1_n169)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_9 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_9), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[9]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[10]), .S(oc8051_sfr1_oc8051_tc1_n170) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_10 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_10), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[10]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[11]), .S(oc8051_sfr1_oc8051_tc1_n171) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_11 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_11), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[11]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[12]), .S(oc8051_sfr1_oc8051_tc1_n172) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_12 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_12), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[12]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[13]), .S(oc8051_sfr1_oc8051_tc1_n173) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_1 ( .A(oc8051_sfr1_tl1[1]), 
        .B(oc8051_sfr1_tl1[0]), .CO(oc8051_sfr1_oc8051_tc1_r372_carry[2]), .S(
        oc8051_sfr1_oc8051_tc1_n1620) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_3 ( .A(oc8051_sfr1_tl1[3]), 
        .B(oc8051_sfr1_oc8051_tc1_r372_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[4]), .S(oc8051_sfr1_oc8051_tc1_n1640) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_2 ( .A(oc8051_sfr1_tl1[2]), 
        .B(oc8051_sfr1_oc8051_tc1_r372_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[3]), .S(oc8051_sfr1_oc8051_tc1_n1630) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_4 ( .A(oc8051_sfr1_tl1[4]), 
        .B(oc8051_sfr1_oc8051_tc1_r372_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[5]), .S(oc8051_sfr1_oc8051_tc1_n165)
         );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u2 ( .A(
        oc8051_sfr1_oc8051_tc1_add_220_carry[7]), .B(oc8051_sfr1_tl1[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n203) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1 ( .A(oc8051_sfr1_tl1[0]), 
        .Y(oc8051_sfr1_oc8051_tc1_n196) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_1 ( .A(oc8051_sfr1_tl1[1]), .B(oc8051_sfr1_tl1[0]), .CO(oc8051_sfr1_oc8051_tc1_add_220_carry[2]), .S(
        oc8051_sfr1_oc8051_tc1_n197) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_3 ( .A(oc8051_sfr1_tl1[3]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[4]), .S(
        oc8051_sfr1_oc8051_tc1_n199) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_2 ( .A(oc8051_sfr1_tl1[2]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[3]), .S(
        oc8051_sfr1_oc8051_tc1_n198) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_4 ( .A(oc8051_sfr1_tl1[4]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[5]), .S(
        oc8051_sfr1_oc8051_tc1_n200) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_5 ( .A(oc8051_sfr1_tl1[5]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[6]), .S(
        oc8051_sfr1_oc8051_tc1_n201) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_6 ( .A(oc8051_sfr1_tl1[6]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[7]), .S(
        oc8051_sfr1_oc8051_tc1_n202) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1 ( .A(oc8051_sfr1_tl0[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n840) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_1 ( .A(oc8051_sfr1_tl0[1]), 
        .B(oc8051_sfr1_tl0[0]), .CO(oc8051_sfr1_oc8051_tc1_r364_carry[2]), .S(
        oc8051_sfr1_oc8051_tc1_n850) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_2 ( .A(oc8051_sfr1_tl0[2]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[3]), .S(oc8051_sfr1_oc8051_tc1_n860)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_3 ( .A(oc8051_sfr1_tl0[3]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[4]), .S(oc8051_sfr1_oc8051_tc1_n870)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_4 ( .A(oc8051_sfr1_tl0[4]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[5]), .S(oc8051_sfr1_oc8051_tc1_n880)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_5 ( .A(oc8051_sfr1_tl0[5]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[6]), .S(oc8051_sfr1_oc8051_tc1_n890)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_6 ( .A(oc8051_sfr1_tl0[6]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[7]), .S(oc8051_sfr1_oc8051_tc1_n900)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_7 ( .A(oc8051_sfr1_tl0[7]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc1_n920), .S(oc8051_sfr1_oc8051_tc1_n910) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_0), .Y(oc8051_sfr1_oc8051_tc1_n470) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_1 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_1), .B(oc8051_sfr1_oc8051_tc1_u3_u1_z_0), .CO(oc8051_sfr1_oc8051_tc1_r360_carry[2]), .S(oc8051_sfr1_oc8051_tc1_n480)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_5 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_5), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[6]), .S(oc8051_sfr1_oc8051_tc1_n520)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_6 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_6), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[7]), .S(oc8051_sfr1_oc8051_tc1_n530)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_7 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_7), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[8]), .S(oc8051_sfr1_oc8051_tc1_n540)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_2 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_2), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[3]), .S(oc8051_sfr1_oc8051_tc1_n490)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_3 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_3), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[4]), .S(oc8051_sfr1_oc8051_tc1_n500)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_4 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_4), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[5]), .S(oc8051_sfr1_oc8051_tc1_n510)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_9 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_9), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[9]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[10]), .S(oc8051_sfr1_oc8051_tc1_n560) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_10 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_10), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[10]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[11]), .S(oc8051_sfr1_oc8051_tc1_n570) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_11 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_11), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[11]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[12]), .S(oc8051_sfr1_oc8051_tc1_n580) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_12 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_12), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[12]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[13]), .S(oc8051_sfr1_oc8051_tc1_n590) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_8 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_8), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[8]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[9]), .S(oc8051_sfr1_oc8051_tc1_n550)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_14 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_14), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[14]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[15]), .S(oc8051_sfr1_oc8051_tc1_n610) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_13 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_13), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[13]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[14]), .S(oc8051_sfr1_oc8051_tc1_n600) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_15 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_15), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[15]), .CO(
        oc8051_sfr1_oc8051_tc1_n630), .S(oc8051_sfr1_oc8051_tc1_n620) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u186 ( .AN(
        oc8051_sfr1_oc8051_tc21_t2ex_r), .B(t2ex_i), .Y(
        oc8051_sfr1_oc8051_tc21_n217) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u185 ( .AN(
        oc8051_sfr1_oc8051_tc21_t2_r), .B(t2_i), .Y(
        oc8051_sfr1_oc8051_tc21_n220) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u184 ( .A(oc8051_sfr1_t2con_3_), 
        .B(oc8051_sfr1_oc8051_tc21_neg_trans), .Y(oc8051_sfr1_oc8051_tc21_n115) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u183 ( .A(oc8051_sfr1_oc8051_tc21_n7), .Y(oc8051_sfr1_tclk) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u182 ( .A(oc8051_sfr1_oc8051_tc21_n8), .Y(oc8051_sfr1_rclk) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u181 ( .A(oc8051_sfr1_tclk), .B(
        oc8051_sfr1_rclk), .Y(oc8051_sfr1_oc8051_tc21_n116) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u180 ( .AN(
        oc8051_sfr1_oc8051_tc21_n116), .B(oc8051_sfr1_t2con_0_), .Y(
        oc8051_sfr1_oc8051_tc21_n11) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u179 ( .A(
        oc8051_sfr1_oc8051_tc21_n11), .Y(oc8051_sfr1_oc8051_tc21_n135) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u178 ( .AN(wr_addr[2]), .B(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_tc21_n34) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u177 ( .A(n_5_net_), .Y(
        oc8051_sfr1_oc8051_tc21_n139) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u176 ( .A(
        oc8051_sfr1_oc8051_tc21_n139), .B(wr_addr[5]), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n138) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u175 ( .A(wr_addr[6]), .B(
        wr_addr[3]), .C(wr_addr[7]), .D(oc8051_sfr1_oc8051_tc21_n138), .Y(
        oc8051_sfr1_oc8051_tc21_n127) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u174 ( .AN(
        oc8051_sfr1_oc8051_tc21_n127), .B(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_tc21_n114) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u173 ( .A(
        oc8051_sfr1_oc8051_tc21_n34), .B(oc8051_sfr1_oc8051_tc21_n114), .C(
        wr_addr[0]), .Y(oc8051_sfr1_oc8051_tc21_n83) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u172 ( .AN(
        oc8051_sfr1_oc8051_tc21_n114), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n113) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u171 ( .A(
        oc8051_sfr1_oc8051_tc21_n113), .B(oc8051_sfr1_oc8051_tc21_n34), .Y(
        oc8051_sfr1_oc8051_tc21_n77) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u170 ( .A(
        oc8051_sfr1_oc8051_tc21_n83), .B(oc8051_sfr1_oc8051_tc21_n77), .Y(
        oc8051_sfr1_oc8051_tc21_n2) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u169 ( .A(oc8051_sfr1_pres_ow), 
        .B(oc8051_sfr1_oc8051_tc21_tc2_event), .S0(oc8051_sfr1_t2con_1_), .Y(
        oc8051_sfr1_oc8051_tc21_n137) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u168 ( .AN(oc8051_sfr1_t2con_2_), 
        .B(oc8051_sfr1_oc8051_tc21_n137), .Y(oc8051_sfr1_oc8051_tc21_n136) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u167 ( .A0(
        oc8051_sfr1_oc8051_tc21_n115), .A1(oc8051_sfr1_oc8051_tc21_n135), .B0(
        oc8051_sfr1_oc8051_tc21_n2), .C0(oc8051_sfr1_oc8051_tc21_n136), .Y(
        oc8051_sfr1_oc8051_tc21_n79) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u166 ( .A(
        oc8051_sfr1_oc8051_tc21_n79), .B(oc8051_sfr1_oc8051_tc21_n116), .Y(
        oc8051_sfr1_oc8051_tc21_n129) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u165 ( .A(oc8051_sfr1_brate2), .B(
        oc8051_sfr1_oc8051_tc21_n850), .S0(oc8051_sfr1_oc8051_tc21_n129), .Y(
        oc8051_sfr1_oc8051_tc21_n128) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u164 ( .A(oc8051_sfr1_tl2[3]), .B(
        oc8051_sfr1_tl2[2]), .C(oc8051_sfr1_tl2[1]), .D(oc8051_sfr1_tl2[0]), 
        .Y(oc8051_sfr1_oc8051_tc21_n131) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u163 ( .A(oc8051_sfr1_tl2[7]), .B(
        oc8051_sfr1_tl2[6]), .C(oc8051_sfr1_tl2[5]), .D(oc8051_sfr1_tl2[4]), 
        .Y(oc8051_sfr1_oc8051_tc21_n132) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u162 ( .A(oc8051_sfr1_th2[3]), .B(
        oc8051_sfr1_th2[2]), .C(oc8051_sfr1_th2[1]), .D(oc8051_sfr1_th2[0]), 
        .Y(oc8051_sfr1_oc8051_tc21_n133) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u161 ( .A(oc8051_sfr1_th2[7]), .B(
        oc8051_sfr1_th2[6]), .C(oc8051_sfr1_th2[5]), .D(oc8051_sfr1_th2[4]), 
        .Y(oc8051_sfr1_oc8051_tc21_n134) );
  OR4_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u160 ( .A(
        oc8051_sfr1_oc8051_tc21_n131), .B(oc8051_sfr1_oc8051_tc21_n132), .C(
        oc8051_sfr1_oc8051_tc21_n133), .D(oc8051_sfr1_oc8051_tc21_n134), .Y(
        oc8051_sfr1_oc8051_tc21_n130) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u159 ( .A(
        oc8051_sfr1_oc8051_tc21_n130), .Y(oc8051_sfr1_oc8051_tc21_n100) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u158 ( .A(
        oc8051_sfr1_oc8051_tc21_n129), .B(oc8051_sfr1_oc8051_tc21_n100), .Y(
        oc8051_sfr1_oc8051_tc21_n101) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u157 ( .A(
        oc8051_sfr1_oc8051_tc21_n128), .B(oc8051_sfr1_oc8051_tc21_n101), .Y(
        oc8051_sfr1_oc8051_tc21_n150) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u156 ( .A(wr_addr[2]), .B(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_tc21_n19) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u155 ( .A(
        oc8051_sfr1_oc8051_tc21_n19), .B(oc8051_sfr1_oc8051_tc21_n113), .Y(
        oc8051_sfr1_oc8051_tc21_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u154 ( .A(
        oc8051_sfr1_oc8051_tc21_n17), .Y(oc8051_sfr1_oc8051_tc21_n122) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u153 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_tc21_n127), .Y(oc8051_sfr1_oc8051_tc21_n121) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u152 ( .A(
        oc8051_sfr1_oc8051_tc21_n121), .Y(oc8051_sfr1_oc8051_tc21_n120) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u151 ( .A(descy), .B(
        oc8051_sfr1_oc8051_tc21_n120), .Y(oc8051_sfr1_oc8051_tc21_n14) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u150 ( .A0(
        oc8051_sfr1_oc8051_tc21_n122), .A1(oc8051_sfr1_oc8051_tc21_n120), .B0(
        oc8051_sfr1_oc8051_tc21_n14), .Y(oc8051_sfr1_oc8051_tc21_n123) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u149 ( .A0(wr_dat[7]), .A1(
        oc8051_sfr1_oc8051_tc21_n122), .B0(oc8051_sfr1_oc8051_tc21_n123), .Y(
        oc8051_sfr1_oc8051_tc21_n124) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u148 ( .AN(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_tc21_n121), .Y(oc8051_sfr1_oc8051_tc21_n23) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u147 ( .A(wr_addr[1]), .B(
        wr_addr[2]), .C(oc8051_sfr1_oc8051_tc21_n23), .Y(
        oc8051_sfr1_oc8051_tc21_n126) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u146 ( .A0(
        oc8051_sfr1_oc8051_tc21_tf2_set), .A1(oc8051_sfr1_oc8051_tc21_n121), 
        .B0(oc8051_sfr1_oc8051_tc21_n122), .C0(oc8051_sfr1_oc8051_tc21_n126), 
        .Y(oc8051_sfr1_oc8051_tc21_n125) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u145 ( .A(
        oc8051_sfr1_oc8051_tc21_n124), .B(oc8051_sfr1_oc8051_tc21_n6), .S0(
        oc8051_sfr1_oc8051_tc21_n125), .Y(oc8051_sfr1_oc8051_tc21_n151) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u144 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_tc21_n122), .B0(oc8051_sfr1_oc8051_tc21_n123), .Y(
        oc8051_sfr1_oc8051_tc21_n117) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u143 ( .A(
        oc8051_sfr1_oc8051_tc21_n121), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n18) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u142 ( .A0(
        oc8051_sfr1_oc8051_tc21_n115), .A1(oc8051_sfr1_oc8051_tc21_tf2_set), 
        .A2(oc8051_sfr1_oc8051_tc21_n120), .B0(oc8051_sfr1_oc8051_tc21_n17), 
        .Y(oc8051_sfr1_oc8051_tc21_n119) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u141 ( .A0(
        oc8051_sfr1_oc8051_tc21_n18), .A1(wr_addr[2]), .A2(wr_addr[1]), .B0(
        oc8051_sfr1_oc8051_tc21_n119), .Y(oc8051_sfr1_oc8051_tc21_n118) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u140 ( .A(
        oc8051_sfr1_oc8051_tc21_n117), .B(oc8051_sfr1_oc8051_tc21_n5), .S0(
        oc8051_sfr1_oc8051_tc21_n118), .Y(oc8051_sfr1_oc8051_tc21_n152) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u139 ( .A(oc8051_sfr1_th2[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n97) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u138 ( .A(oc8051_sfr1_t2con_0_), 
        .B(oc8051_sfr1_oc8051_tc21_n116), .Y(oc8051_sfr1_oc8051_tc21_n99) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u137 ( .A(
        oc8051_sfr1_oc8051_tc21_n99), .Y(oc8051_sfr1_oc8051_tc21_n10) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u136 ( .A(
        oc8051_sfr1_oc8051_tc21_n115), .Y(oc8051_sfr1_oc8051_tc21_n102) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u135 ( .AN(wr_addr[1]), .B(
        wr_addr[2]), .Y(oc8051_sfr1_oc8051_tc21_n27) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u134 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_tc21_n114), .C(oc8051_sfr1_oc8051_tc21_n27), .Y(
        oc8051_sfr1_oc8051_tc21_n105) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u133 ( .A(
        oc8051_sfr1_oc8051_tc21_n27), .B(oc8051_sfr1_oc8051_tc21_n113), .Y(
        oc8051_sfr1_oc8051_tc21_n43) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u132 ( .A(
        oc8051_sfr1_oc8051_tc21_n10), .B(oc8051_sfr1_oc8051_tc21_n102), .C(
        oc8051_sfr1_oc8051_tc21_n105), .D(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n39) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u131 ( .A(oc8051_sfr1_rcap2h[7]), 
        .Y(oc8051_sfr1_oc8051_tc21_n112) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u130 ( .A(
        oc8051_sfr1_oc8051_tc21_n105), .B(oc8051_sfr1_oc8051_tc21_n39), .Y(
        oc8051_sfr1_oc8051_tc21_n104) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u129 ( .A(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n64) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u128 ( .A0(
        oc8051_sfr1_oc8051_tc21_n97), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n112), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n64), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n153) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u127 ( .A(oc8051_sfr1_th2[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n95) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u126 ( .A(oc8051_sfr1_rcap2h[6]), 
        .Y(oc8051_sfr1_oc8051_tc21_n111) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u125 ( .A(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n61) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u124 ( .A0(
        oc8051_sfr1_oc8051_tc21_n95), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n111), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n61), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n154) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u123 ( .A(oc8051_sfr1_th2[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n93) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u122 ( .A(oc8051_sfr1_rcap2h[5]), 
        .Y(oc8051_sfr1_oc8051_tc21_n110) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u121 ( .A(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n58) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u120 ( .A0(
        oc8051_sfr1_oc8051_tc21_n93), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n110), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n58), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n155) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u119 ( .A(oc8051_sfr1_th2[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n91) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u118 ( .A(oc8051_sfr1_rcap2h[4]), 
        .Y(oc8051_sfr1_oc8051_tc21_n109) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u117 ( .A(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n55) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u116 ( .A0(
        oc8051_sfr1_oc8051_tc21_n91), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n109), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n55), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n156) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u115 ( .A(oc8051_sfr1_th2[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n89) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u114 ( .A(oc8051_sfr1_rcap2h[3]), 
        .Y(oc8051_sfr1_oc8051_tc21_n108) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u113 ( .A(wr_dat[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n52) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u112 ( .A0(
        oc8051_sfr1_oc8051_tc21_n89), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n108), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n52), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n157) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u111 ( .A(oc8051_sfr1_th2[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n87) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u110 ( .A(oc8051_sfr1_rcap2h[2]), 
        .Y(oc8051_sfr1_oc8051_tc21_n107) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u109 ( .A(wr_dat[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n49) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u108 ( .A0(
        oc8051_sfr1_oc8051_tc21_n87), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n107), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n49), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n158) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u107 ( .A(oc8051_sfr1_th2[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u106 ( .A(oc8051_sfr1_rcap2h[1]), 
        .Y(oc8051_sfr1_oc8051_tc21_n106) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u105 ( .A(wr_dat[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n46) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u104 ( .A0(
        oc8051_sfr1_oc8051_tc21_n85), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n106), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n46), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u103 ( .A(oc8051_sfr1_th2[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n81) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u102 ( .A(oc8051_sfr1_rcap2h[0]), 
        .Y(oc8051_sfr1_oc8051_tc21_n103) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u101 ( .A(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n42) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u100 ( .A0(
        oc8051_sfr1_oc8051_tc21_n81), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n103), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n42), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n160) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u99 ( .A(
        oc8051_sfr1_oc8051_tc21_n11), .B(oc8051_sfr1_oc8051_tc21_n102), .C(
        oc8051_sfr1_oc8051_tc21_n2), .Y(oc8051_sfr1_oc8051_tc21_n80) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u98 ( .A(
        oc8051_sfr1_oc8051_tc21_n79), .B(oc8051_sfr1_oc8051_tc21_n83), .C(
        oc8051_sfr1_oc8051_tc21_n80), .Y(oc8051_sfr1_oc8051_tc21_n82) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u97 ( .A(oc8051_sfr1_oc8051_tc21_n79), .Y(oc8051_sfr1_oc8051_tc21_n12) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u96 ( .A(
        oc8051_sfr1_oc8051_tc21_n100), .B(oc8051_sfr1_oc8051_tc21_n11), .C(
        oc8051_sfr1_oc8051_tc21_n12), .Y(oc8051_sfr1_oc8051_tc21_n9) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u95 ( .A(
        oc8051_sfr1_oc8051_tc21_n101), .B(oc8051_sfr1_oc8051_tc21_n9), .C(
        oc8051_sfr1_oc8051_tc21_n80), .Y(oc8051_sfr1_oc8051_tc21_n78) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u94 ( .A0(
        oc8051_sfr1_oc8051_tc21_n99), .A1(oc8051_sfr1_oc8051_tc21_n100), .B0(
        oc8051_sfr1_oc8051_tc21_n79), .Y(oc8051_sfr1_oc8051_tc21_n68) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u93 ( .A0(oc8051_sfr1_rcap2h[7]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n840), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n98) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u92 ( .A0(
        oc8051_sfr1_oc8051_tc21_n97), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n64), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n98), .Y(oc8051_sfr1_oc8051_tc21_n161) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u91 ( .A0(oc8051_sfr1_rcap2h[6]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n830), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n96) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u90 ( .A0(
        oc8051_sfr1_oc8051_tc21_n95), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n61), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n96), .Y(oc8051_sfr1_oc8051_tc21_n162) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u89 ( .A0(oc8051_sfr1_rcap2h[5]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n820), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n94) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u88 ( .A0(
        oc8051_sfr1_oc8051_tc21_n93), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n58), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n94), .Y(oc8051_sfr1_oc8051_tc21_n163) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u87 ( .A0(oc8051_sfr1_rcap2h[4]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n810), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n92) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u86 ( .A0(
        oc8051_sfr1_oc8051_tc21_n91), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n55), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n92), .Y(oc8051_sfr1_oc8051_tc21_n164) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u85 ( .A0(oc8051_sfr1_rcap2h[3]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n800), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n90) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u84 ( .A0(
        oc8051_sfr1_oc8051_tc21_n89), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n52), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n90), .Y(oc8051_sfr1_oc8051_tc21_n165) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u83 ( .A0(oc8051_sfr1_rcap2h[2]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n790), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n88) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u82 ( .A0(
        oc8051_sfr1_oc8051_tc21_n87), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n49), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n88), .Y(oc8051_sfr1_oc8051_tc21_n166) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u81 ( .A0(oc8051_sfr1_rcap2h[1]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n780), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n86) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u80 ( .A0(
        oc8051_sfr1_oc8051_tc21_n85), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n46), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n86), .Y(oc8051_sfr1_oc8051_tc21_n167) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u79 ( .A0(oc8051_sfr1_rcap2h[0]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n770), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n84) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u78 ( .A0(
        oc8051_sfr1_oc8051_tc21_n81), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n42), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n84), .Y(oc8051_sfr1_oc8051_tc21_n168) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u77 ( .A(oc8051_sfr1_tl2[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n62) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u76 ( .A(
        oc8051_sfr1_oc8051_tc21_n79), .B(oc8051_sfr1_oc8051_tc21_n77), .C(
        oc8051_sfr1_oc8051_tc21_n80), .Y(oc8051_sfr1_oc8051_tc21_n65) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u75 ( .A(oc8051_sfr1_oc8051_tc21_n78), .Y(oc8051_sfr1_oc8051_tc21_n66) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u74 ( .A(oc8051_sfr1_rcap2l[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n63) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u73 ( .A(oc8051_sfr1_oc8051_tc21_n77), .Y(oc8051_sfr1_oc8051_tc21_n69) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u72 ( .A0(
        oc8051_sfr1_oc8051_tc21_n760), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n76) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u71 ( .A0(
        oc8051_sfr1_oc8051_tc21_n62), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n63), .C0(
        oc8051_sfr1_oc8051_tc21_n76), .Y(oc8051_sfr1_oc8051_tc21_n169) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u70 ( .A(oc8051_sfr1_tl2[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n59) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u69 ( .A(oc8051_sfr1_rcap2l[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n60) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u68 ( .A0(
        oc8051_sfr1_oc8051_tc21_n750), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n75) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u67 ( .A0(
        oc8051_sfr1_oc8051_tc21_n59), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n60), .C0(
        oc8051_sfr1_oc8051_tc21_n75), .Y(oc8051_sfr1_oc8051_tc21_n170) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u66 ( .A(oc8051_sfr1_tl2[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n56) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u65 ( .A(oc8051_sfr1_rcap2l[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n57) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u64 ( .A0(
        oc8051_sfr1_oc8051_tc21_n740), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n74) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u63 ( .A0(
        oc8051_sfr1_oc8051_tc21_n56), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n57), .C0(
        oc8051_sfr1_oc8051_tc21_n74), .Y(oc8051_sfr1_oc8051_tc21_n171) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u62 ( .A(oc8051_sfr1_tl2[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n53) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u61 ( .A(oc8051_sfr1_rcap2l[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n54) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u60 ( .A0(
        oc8051_sfr1_oc8051_tc21_n730), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n73) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u59 ( .A0(
        oc8051_sfr1_oc8051_tc21_n53), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n54), .C0(
        oc8051_sfr1_oc8051_tc21_n73), .Y(oc8051_sfr1_oc8051_tc21_n172) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u58 ( .A(oc8051_sfr1_tl2[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n50) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u57 ( .A(oc8051_sfr1_rcap2l[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n51) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u56 ( .A0(
        oc8051_sfr1_oc8051_tc21_n720), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n72) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u55 ( .A0(
        oc8051_sfr1_oc8051_tc21_n50), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n51), .C0(
        oc8051_sfr1_oc8051_tc21_n72), .Y(oc8051_sfr1_oc8051_tc21_n173) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u54 ( .A(oc8051_sfr1_tl2[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n47) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u53 ( .A(oc8051_sfr1_rcap2l[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n48) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u52 ( .A0(
        oc8051_sfr1_oc8051_tc21_n710), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n71) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u51 ( .A0(
        oc8051_sfr1_oc8051_tc21_n47), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n48), .C0(
        oc8051_sfr1_oc8051_tc21_n71), .Y(oc8051_sfr1_oc8051_tc21_n174) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u50 ( .A(oc8051_sfr1_tl2[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n44) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u49 ( .A(oc8051_sfr1_rcap2l[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n45) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u48 ( .A0(
        oc8051_sfr1_oc8051_tc21_n700), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n70) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u47 ( .A0(
        oc8051_sfr1_oc8051_tc21_n44), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n45), .C0(
        oc8051_sfr1_oc8051_tc21_n70), .Y(oc8051_sfr1_oc8051_tc21_n175) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u46 ( .A(oc8051_sfr1_tl2[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n38) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u45 ( .A(oc8051_sfr1_rcap2l[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n41) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u44 ( .A0(
        oc8051_sfr1_oc8051_tc21_n690), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n67) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u43 ( .A0(
        oc8051_sfr1_oc8051_tc21_n38), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n41), .C0(
        oc8051_sfr1_oc8051_tc21_n67), .Y(oc8051_sfr1_oc8051_tc21_n176) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u42 ( .A(
        oc8051_sfr1_oc8051_tc21_n43), .B(oc8051_sfr1_oc8051_tc21_n39), .Y(
        oc8051_sfr1_oc8051_tc21_n40) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u41 ( .A0(
        oc8051_sfr1_oc8051_tc21_n62), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n63), .C0(
        oc8051_sfr1_oc8051_tc21_n43), .C1(oc8051_sfr1_oc8051_tc21_n64), .Y(
        oc8051_sfr1_oc8051_tc21_n177) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u40 ( .A0(
        oc8051_sfr1_oc8051_tc21_n59), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n60), .C0(
        oc8051_sfr1_oc8051_tc21_n43), .C1(oc8051_sfr1_oc8051_tc21_n61), .Y(
        oc8051_sfr1_oc8051_tc21_n178) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u39 ( .A0(
        oc8051_sfr1_oc8051_tc21_n56), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n57), .C0(
        oc8051_sfr1_oc8051_tc21_n58), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n179) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u38 ( .A0(
        oc8051_sfr1_oc8051_tc21_n53), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n54), .C0(
        oc8051_sfr1_oc8051_tc21_n55), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n180) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u37 ( .A0(
        oc8051_sfr1_oc8051_tc21_n50), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n51), .C0(
        oc8051_sfr1_oc8051_tc21_n52), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n181) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u36 ( .A0(
        oc8051_sfr1_oc8051_tc21_n47), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n48), .C0(
        oc8051_sfr1_oc8051_tc21_n49), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n182) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u35 ( .A0(
        oc8051_sfr1_oc8051_tc21_n44), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n45), .C0(
        oc8051_sfr1_oc8051_tc21_n46), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n183) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u34 ( .A0(
        oc8051_sfr1_oc8051_tc21_n38), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n41), .C0(
        oc8051_sfr1_oc8051_tc21_n42), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n184) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u33 ( .A(
        oc8051_sfr1_oc8051_tc21_n23), .B(oc8051_sfr1_oc8051_tc21_n34), .Y(
        oc8051_sfr1_oc8051_tc21_n35) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u32 ( .A(
        oc8051_sfr1_oc8051_tc21_n35), .B(oc8051_sfr1_rclk), .Y(
        oc8051_sfr1_oc8051_tc21_n37) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u31 ( .A(wr_dat[5]), .B(
        oc8051_sfr1_oc8051_tc21_n37), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n36) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u30 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n35), .B0(
        oc8051_sfr1_oc8051_tc21_n36), .Y(oc8051_sfr1_oc8051_tc21_n185) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u29 ( .A(
        oc8051_sfr1_oc8051_tc21_n18), .B(oc8051_sfr1_oc8051_tc21_n34), .Y(
        oc8051_sfr1_oc8051_tc21_n31) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u28 ( .A(
        oc8051_sfr1_oc8051_tc21_n31), .B(oc8051_sfr1_tclk), .Y(
        oc8051_sfr1_oc8051_tc21_n33) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u27 ( .A(wr_dat[4]), .B(
        oc8051_sfr1_oc8051_tc21_n33), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n32) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u26 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n31), .B0(
        oc8051_sfr1_oc8051_tc21_n32), .Y(oc8051_sfr1_oc8051_tc21_n186) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u25 ( .A(
        oc8051_sfr1_oc8051_tc21_n27), .B(oc8051_sfr1_oc8051_tc21_n23), .Y(
        oc8051_sfr1_oc8051_tc21_n28) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u24 ( .A(
        oc8051_sfr1_oc8051_tc21_n28), .B(oc8051_sfr1_t2con_3_), .Y(
        oc8051_sfr1_oc8051_tc21_n30) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u23 ( .A(wr_dat[3]), .B(
        oc8051_sfr1_oc8051_tc21_n30), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n29) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u22 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n28), .B0(
        oc8051_sfr1_oc8051_tc21_n29), .Y(oc8051_sfr1_oc8051_tc21_n187) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u21 ( .A(
        oc8051_sfr1_oc8051_tc21_n27), .B(oc8051_sfr1_oc8051_tc21_n18), .Y(
        oc8051_sfr1_oc8051_tc21_n24) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u20 ( .A(
        oc8051_sfr1_oc8051_tc21_n24), .B(oc8051_sfr1_t2con_2_), .Y(
        oc8051_sfr1_oc8051_tc21_n26) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u19 ( .A(wr_dat[2]), .B(
        oc8051_sfr1_oc8051_tc21_n26), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n25) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u18 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n24), .B0(
        oc8051_sfr1_oc8051_tc21_n25), .Y(oc8051_sfr1_oc8051_tc21_n188) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u17 ( .A(
        oc8051_sfr1_oc8051_tc21_n23), .B(oc8051_sfr1_oc8051_tc21_n19), .Y(
        oc8051_sfr1_oc8051_tc21_n20) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u16 ( .A(
        oc8051_sfr1_oc8051_tc21_n20), .B(oc8051_sfr1_t2con_1_), .Y(
        oc8051_sfr1_oc8051_tc21_n22) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u15 ( .A(wr_dat[1]), .B(
        oc8051_sfr1_oc8051_tc21_n22), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n21) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u14 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n20), .B0(
        oc8051_sfr1_oc8051_tc21_n21), .Y(oc8051_sfr1_oc8051_tc21_n189) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u13 ( .A(
        oc8051_sfr1_oc8051_tc21_n18), .B(oc8051_sfr1_oc8051_tc21_n19), .Y(
        oc8051_sfr1_oc8051_tc21_n13) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u12 ( .A(
        oc8051_sfr1_oc8051_tc21_n13), .B(oc8051_sfr1_t2con_0_), .Y(
        oc8051_sfr1_oc8051_tc21_n16) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u11 ( .A(wr_dat[0]), .B(
        oc8051_sfr1_oc8051_tc21_n16), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n15) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u10 ( .A0(
        oc8051_sfr1_oc8051_tc21_n13), .A1(oc8051_sfr1_oc8051_tc21_n14), .B0(
        oc8051_sfr1_oc8051_tc21_n15), .Y(oc8051_sfr1_oc8051_tc21_n190) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u9 ( .A(
        oc8051_sfr1_oc8051_tc21_tf2_set), .Y(oc8051_sfr1_oc8051_tc21_n3) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u8 ( .A0(
        oc8051_sfr1_oc8051_tc21_n10), .A1(oc8051_sfr1_oc8051_tc21_n11), .B0(
        oc8051_sfr1_oc8051_tc21_n12), .C0(oc8051_sfr1_oc8051_tc21_n850), .Y(
        oc8051_sfr1_oc8051_tc21_n4) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u7 ( .A0(
        oc8051_sfr1_oc8051_tc21_n2), .A1(oc8051_sfr1_oc8051_tc21_n3), .B0(
        oc8051_sfr1_oc8051_tc21_n4), .C0(oc8051_sfr1_oc8051_tc21_n9), .Y(
        oc8051_sfr1_oc8051_tc21_n191) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u6 ( .A(oc8051_sfr1_oc8051_tc21_n5), 
        .Y(oc8051_sfr1_t2con_6_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u5 ( .A(oc8051_sfr1_oc8051_tc21_n6), 
        .Y(oc8051_sfr1_t2con_7_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u4 ( .A(oc8051_sfr1_oc8051_tc21_n5), .B(oc8051_sfr1_oc8051_tc21_n6), .Y(oc8051_sfr1_tc2_int) );
  TIELO_X1M_A12TS oc8051_sfr1_oc8051_tc21_u3 ( .Y(oc8051_sfr1_oc8051_tc21_n1)
         );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n152), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n5) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n151), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n6) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n186), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n7) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n185), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n8) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n176), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n169), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n173), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n161), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n165), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n172), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n164), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n168), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n171), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n175), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n170), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n174), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n163), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n167), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n162), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n166), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n190), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n189), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n187), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n188), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tf2_set_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n191), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_tc21_tf2_set) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n153), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n154), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n155), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n156), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n157), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n158), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n159), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n160), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_brate2_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n150), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_brate2) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n183), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n177), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n178), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n179), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n180), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n181), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n182), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n184), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tc2_event_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n220), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_tc21_tc2_event) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_neg_trans_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n217), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_tc21_neg_trans) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2_r_reg ( .D(t2_i), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc21_t2_r) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2ex_r_reg ( .D(t2ex_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc21_t2ex_r) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1 ( .A(oc8051_sfr1_tl2[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n690) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_1 ( .A(oc8051_sfr1_tl2[1]), 
        .B(oc8051_sfr1_tl2[0]), .CO(oc8051_sfr1_oc8051_tc21_r320_carry[2]), 
        .S(oc8051_sfr1_oc8051_tc21_n700) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_2 ( .A(oc8051_sfr1_tl2[2]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[3]), .S(
        oc8051_sfr1_oc8051_tc21_n710) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_3 ( .A(oc8051_sfr1_tl2[3]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[4]), .S(
        oc8051_sfr1_oc8051_tc21_n720) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_4 ( .A(oc8051_sfr1_tl2[4]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[5]), .S(
        oc8051_sfr1_oc8051_tc21_n730) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_5 ( .A(oc8051_sfr1_tl2[5]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[6]), .S(
        oc8051_sfr1_oc8051_tc21_n740) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_6 ( .A(oc8051_sfr1_tl2[6]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[7]), .S(
        oc8051_sfr1_oc8051_tc21_n750) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_7 ( .A(oc8051_sfr1_tl2[7]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[8]), .S(
        oc8051_sfr1_oc8051_tc21_n760) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_8 ( .A(oc8051_sfr1_th2[0]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[8]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[9]), .S(
        oc8051_sfr1_oc8051_tc21_n770) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_9 ( .A(oc8051_sfr1_th2[1]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[9]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[10]), .S(
        oc8051_sfr1_oc8051_tc21_n780) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_10 ( .A(oc8051_sfr1_th2[2]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[10]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[11]), .S(
        oc8051_sfr1_oc8051_tc21_n790) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_11 ( .A(oc8051_sfr1_th2[3]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[11]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[12]), .S(
        oc8051_sfr1_oc8051_tc21_n800) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_12 ( .A(oc8051_sfr1_th2[4]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[12]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[13]), .S(
        oc8051_sfr1_oc8051_tc21_n810) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_13 ( .A(oc8051_sfr1_th2[5]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[13]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[14]), .S(
        oc8051_sfr1_oc8051_tc21_n820) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_14 ( .A(oc8051_sfr1_th2[6]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[14]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[15]), .S(
        oc8051_sfr1_oc8051_tc21_n830) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_15 ( .A(oc8051_sfr1_th2[7]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[15]), .CO(
        oc8051_sfr1_oc8051_tc21_n850), .S(oc8051_sfr1_oc8051_tc21_n840) );
endmodule

