
module cpu8080 ( addr, data_in, data_out, readmem, writemem, readio, writeio, intr, inta, 
        waitr, reset, clock );
  output [15:0] addr;

  input [7:0] data_in;
  output [7:0] data_out;

  input intr, waitr, reset, clock;
  output readmem, writemem, readio, writeio, inta;
  wire   n46, n233, n234, n235, n236, n237, aluoprb_0_, alucin, alucout,
         aluzout, alusout, alupar, aluaxc, ei, eienb, carry, regfil_2__7_,
         regfil_2__6_, regfil_2__5_, regfil_2__4_, regfil_2__3_, regfil_2__2_,
         regfil_2__1_, regfil_2__0_, regfil_6__7_, regfil_6__6_, regfil_6__5_,
         regfil_6__4_, regfil_6__3_, regfil_6__2_, regfil_6__1_, regfil_6__0_,
         regfil_7__0_, auxcar, n240, n241, n242, n243, n244, n245, n246, n247,
         sign, zero, parity, intcyc, n963, n964, n965, n966, n967, n968, n969,
         n970, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n26580, n26590, n26600, n26610,
         n26620, n26630, n26640, n26650, n26660, n26670, n26680, n26690,
         n26700, n26710, n26720, n30100, n30110, n30120, n30130, n30140,
         n30150, n30160, n30170, n30180, n30190, n30200, n30210, n30220,
         n30230, n30240, n31370, n31390, n31400, n31410, n31420, n31430,
         n31440, n31450, n31460, n31470, n31480, n31490, n31500, n31510,
         n31520, n35710, n35720, n35730, n35740, n35750, u3_u79_z_0,
         u3_u79_z_1, u3_u79_z_2, u3_u79_z_3, u3_u79_z_4, u3_u79_z_5,
         u3_u79_z_6, u3_u79_z_7, u3_u79_z_8, u3_u79_z_9, u3_u79_z_10,
         u3_u79_z_11, u3_u79_z_12, u3_u79_z_13, u3_u79_z_14, u3_u79_z_15,
         u3_u80_z_0, u3_u80_z_1, u3_u80_z_2, u3_u80_z_3, u3_u80_z_4,
         u3_u80_z_5, u3_u80_z_6, u3_u80_z_7, u3_u80_z_8, u3_u80_z_9,
         u3_u80_z_10, u3_u80_z_11, u3_u80_z_12, u3_u80_z_13, u3_u80_z_14,
         u3_u80_z_15, u3_u84_z_0, u3_u84_z_1, u3_u84_z_2, u3_u84_z_3,
         u3_u84_z_4, u3_u84_z_5, u3_u84_z_6, u3_u84_z_7, u3_u84_z_8,
         u3_u84_z_9, u3_u84_z_10, u3_u84_z_11, u3_u84_z_12, u3_u84_z_13,
         u3_u84_z_14, u3_u84_z_15, u3_u85_z_1, u3_u85_z_2, u3_u85_z_3,
         u3_u85_z_4, u3_u85_z_5, u3_u85_z_6, u3_u85_z_7, u3_u85_z_8,
         u3_u87_z_0, u3_u88_z_0, u3_u88_z_1, u3_u88_z_2, u3_u88_z_3,
         u3_u88_z_4, u3_u88_z_5, u3_u88_z_6, u3_u88_z_7, u3_u88_z_8,
         u3_u88_z_9, u3_u88_z_10, u3_u88_z_11, u3_u88_z_12, u3_u88_z_13,
         u3_u88_z_14, u3_u88_z_15, u3_u92_z_0, u3_u92_z_1, u3_u92_z_2,
         u3_u92_z_3, u3_u92_z_4, u3_u92_z_5, u3_u92_z_6, u3_u92_z_7,
         u3_u93_z_6, u3_u94_z_0, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n26581, n26591, n26601, n26611,
         n26621, n26631, n26641, n26651, n26661, n26671, n26681, n26691,
         n26701, n26711, n26721, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, r1226_sum_1_, r1226_sum_2_, r1226_sum_3_,
         r1226_sum_4_, r1226_sum_5_, r1226_sum_6_, r1226_sum_7_, r1226_sum_8_,
         r1226_sum_9_, r1226_sum_10_, r1226_sum_11_, r1226_sum_12_,
         r1226_sum_13_, r1226_sum_14_, r1226_sum_15_, r1298_carry_1_,
         r1298_carry_2_, r1298_carry_3_, r1298_carry_4_, r1298_carry_5_,
         r1298_carry_6_, r1298_carry_7_, r1298_carry_8_, r1298_carry_9_,
         r1298_carry_10_, r1298_carry_11_, r1298_carry_12_, r1298_carry_13_,
         r1298_carry_14_, r1298_carry_15_, r1606_b_as_0_, r1606_b_as_2_,
         r1606_b_as_6_, r1606_carry_1_, r1606_carry_2_, r1606_carry_3_,
         r1606_carry_4_, r1606_carry_5_, r1606_carry_6_, r1606_carry_7_,
         r1606_carry_8_, r1606_sum_0_, r1606_sum_1_, r1606_sum_2_,
         r1606_sum_3_, r1606_sum_4_, r1606_sum_5_, r1606_sum_6_, r1606_sum_7_,
         r1606_sum_8_, r201_carry_1_, r201_carry_2_, r201_carry_3_,
         r201_carry_4_, r201_carry_5_, r201_carry_6_, r201_carry_7_,
         r201_carry_8_, r201_carry_9_, r201_carry_10_, r201_carry_11_,
         r201_carry_12_, r201_carry_13_, r201_carry_14_, r201_carry_15_,
         r201_sum_0_, r201_sum_1_, r201_sum_2_, r201_sum_3_, r201_sum_4_,
         r201_sum_5_, r201_sum_6_, r201_sum_7_, r201_sum_8_, r201_sum_9_,
         r201_sum_10_, r201_sum_11_, r201_sum_12_, r201_sum_13_, r201_sum_14_,
         r201_sum_15_, r201_a_0_, r201_a_9_, r201_a_10_, r201_a_11_,
         r201_a_12_, r201_a_13_, r201_a_14_, r201_a_15_, r194_carry_1_,
         r194_carry_2_, r194_carry_3_, r194_carry_4_, r194_carry_5_,
         r194_carry_6_, r194_carry_7_, r194_carry_8_, r194_carry_9_,
         r194_carry_10_, r194_carry_11_, r194_carry_12_, r194_carry_13_,
         r194_carry_14_, r194_carry_15_, r194_sum_0_, r194_sum_1_, r194_sum_2_,
         r194_sum_3_, r194_sum_4_, r194_sum_5_, r194_sum_6_, r194_sum_7_,
         r194_sum_8_, r194_sum_9_, r194_sum_10_, r194_sum_11_, r194_sum_12_,
         r194_sum_13_, r194_sum_14_, r194_sum_15_, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n30101, n30111, n30121, n30131, n30141,
         n30151, n30161, n30171, n30181, n30191, n30201, n30211, n30221,
         n30231, n30241, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n31371, n3138, n31391, n31401,
         n31411, n31421, n31431, n31441, n31451, n31461, n31471, n31481,
         n31491, n31501, n31511, n31521, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n35711, n35721, n35731, n35741, n35751, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4313, n4314, n4315, n4316, n4318,
         alu_n42, alu_n41, alu_n40, alu_n39, alu_n38, alu_n37, alu_n35,
         alu_n34, alu_n33, alu_n32, alu_n31, alu_n30, alu_n29, alu_n28,
         alu_n27, alu_n26, alu_n25, alu_n24, alu_n23, alu_n22, alu_n21,
         alu_n20, alu_n19, alu_n18, alu_n17, alu_n16, alu_n15, alu_n14,
         alu_n13, alu_n12, alu_n11, alu_n10, alu_n9, alu_n8, alu_n7, alu_n6,
         alu_n5, alu_n4, alu_n3, alu_n2, alu_n1, alu_n36, alu_u2_u4_z_0,
         alu_u2_u3_z_0, alu_n100, alu_n99, alu_n98, alu_n97, alu_n96, alu_n95,
         alu_n94, alu_n93, alu_n92, alu_n91, alu_resi_0_, alu_resi_1_,
         alu_resi_2_, alu_resi_4_, alu_resi_6_, alu_n330, alu_n320, alu_n310,
         alu_n300, alu_n290, alu_n280, alu_n270, alu_n260, alu_n250, alu_n240,
         alu_n230, alu_n220, alu_n210, alu_n200, alu_n190, alu_n180, alu_n170,
         alu_n160, alu_n150, alu_n140, alu_n130, alu_n120, alu_n110, alu_n101,
         alu_r24_b_as_0_, alu_r24_b_as_1_, alu_r24_b_as_2_, alu_r24_b_as_3_,
         alu_r24_b_as_4_, alu_r24_b_as_5_, alu_r24_b_as_6_, alu_r24_b_as_7_,
         alu_r373_n13, alu_r373_n12, alu_r373_n11, alu_r373_n10, alu_r373_n9,
         alu_r373_n8, alu_r373_n7, alu_r373_n6, alu_r373_n5, alu_r373_n4,
         alu_r373_n3, alu_r373_n2, alu_r373_n1, alu_r373_carry_4_, r1610_n1,
         r1610_carry_2_, r1610_carry_3_, r1610_carry_4_, r1610_carry_5_,
         r1610_carry_6_, r1610_carry_7_, r1610_carry_8_, r1610_carry_9_,
         r1610_carry_10_, r1610_carry_11_, r1610_carry_12_, r1610_carry_13_,
         r1610_carry_14_, r1610_carry_15_;
  wire   [7:0] alures;
  wire   [7:0] aluopra;
  wire   [2:0] alusel;
  wire   [15:0] pc;
  wire   [5:0] state;
  wire   [7:6] opcode;
  wire   [15:1] sp;
  wire   [5:0] statesel;
  wire   [15:0] raddrhold;
  wire   [7:0] rdatahold;
  wire   [7:0] rdatahold2;
  wire   [1:0] popdes;
  wire   [2:0] regd;
  wire   [7:0] datao;
  wire   [1:0] r201_b_as;
  wire   [1:0] r194_b_as;
  wire   [8:0] alu_r24_carry;

  ADDF_X1M_A12TR r1298_u1_1 ( .A(sp[1]), .B(n4307), .CI(r1298_carry_1_), .CO(
        r1298_carry_2_), .S(n26580) );
  ADDF_X1M_A12TR r1298_u1_2 ( .A(sp[2]), .B(r1298_carry_1_), .CI(
        r1298_carry_2_), .CO(r1298_carry_3_), .S(n26590) );
  ADDF_X1M_A12TR r1298_u1_3 ( .A(sp[3]), .B(r1298_carry_1_), .CI(
        r1298_carry_3_), .CO(r1298_carry_4_), .S(n26600) );
  ADDF_X1M_A12TR r1298_u1_4 ( .A(sp[4]), .B(r1298_carry_1_), .CI(
        r1298_carry_4_), .CO(r1298_carry_5_), .S(n26610) );
  ADDF_X1M_A12TR r1298_u1_5 ( .A(sp[5]), .B(r1298_carry_1_), .CI(
        r1298_carry_5_), .CO(r1298_carry_6_), .S(n26620) );
  ADDF_X1M_A12TR r1298_u1_6 ( .A(sp[6]), .B(r1298_carry_1_), .CI(
        r1298_carry_6_), .CO(r1298_carry_7_), .S(n26630) );
  ADDF_X1M_A12TR r1298_u1_7 ( .A(sp[7]), .B(r1298_carry_1_), .CI(
        r1298_carry_7_), .CO(r1298_carry_8_), .S(n26640) );
  ADDF_X1M_A12TR r1298_u1_8 ( .A(sp[8]), .B(r1298_carry_1_), .CI(
        r1298_carry_8_), .CO(r1298_carry_9_), .S(n26650) );
  ADDF_X1M_A12TR r1298_u1_9 ( .A(sp[9]), .B(r1298_carry_1_), .CI(
        r1298_carry_9_), .CO(r1298_carry_10_), .S(n26660) );
  ADDF_X1M_A12TR r1298_u1_10 ( .A(sp[10]), .B(r1298_carry_1_), .CI(
        r1298_carry_10_), .CO(r1298_carry_11_), .S(n26670) );
  ADDF_X1M_A12TR r1298_u1_11 ( .A(sp[11]), .B(r1298_carry_1_), .CI(
        r1298_carry_11_), .CO(r1298_carry_12_), .S(n26680) );
  ADDF_X1M_A12TR r1298_u1_12 ( .A(sp[12]), .B(r1298_carry_1_), .CI(
        r1298_carry_12_), .CO(r1298_carry_13_), .S(n26690) );
  ADDF_X1M_A12TR r1298_u1_13 ( .A(sp[13]), .B(r1298_carry_1_), .CI(
        r1298_carry_13_), .CO(r1298_carry_14_), .S(n26700) );
  ADDF_X1M_A12TR r1298_u1_14 ( .A(sp[14]), .B(r1298_carry_1_), .CI(
        r1298_carry_14_), .CO(r1298_carry_15_), .S(n26710) );
  ADDF_X1M_A12TR r1298_u1_15 ( .A(sp[15]), .B(r1298_carry_1_), .CI(
        r1298_carry_15_), .CO(), .S(n26720) );
  ADDF_X1M_A12TR r1606_u1_0 ( .A(u3_u92_z_0), .B(r1606_b_as_0_), .CI(
        u3_u94_z_0), .CO(r1606_carry_1_), .S(r1606_sum_0_) );
  ADDF_X1M_A12TR r1606_u1_1 ( .A(u3_u92_z_1), .B(r1606_b_as_2_), .CI(
        r1606_carry_1_), .CO(r1606_carry_2_), .S(r1606_sum_1_) );
  ADDF_X1M_A12TR r1606_u1_2 ( .A(u3_u92_z_2), .B(r1606_b_as_2_), .CI(
        r1606_carry_2_), .CO(r1606_carry_3_), .S(r1606_sum_2_) );
  ADDF_X1M_A12TR r1606_u1_3 ( .A(u3_u92_z_3), .B(u3_u94_z_0), .CI(
        r1606_carry_3_), .CO(r1606_carry_4_), .S(r1606_sum_3_) );
  ADDF_X1M_A12TR r1606_u1_4 ( .A(u3_u92_z_4), .B(u3_u94_z_0), .CI(
        r1606_carry_4_), .CO(r1606_carry_5_), .S(r1606_sum_4_) );
  ADDF_X1M_A12TR r1606_u1_5 ( .A(u3_u92_z_5), .B(r1606_b_as_6_), .CI(
        r1606_carry_5_), .CO(r1606_carry_6_), .S(r1606_sum_5_) );
  ADDF_X1M_A12TR r1606_u1_6 ( .A(u3_u92_z_6), .B(r1606_b_as_6_), .CI(
        r1606_carry_6_), .CO(r1606_carry_7_), .S(r1606_sum_6_) );
  ADDF_X1M_A12TR r1606_u1_7 ( .A(u3_u92_z_7), .B(u3_u94_z_0), .CI(
        r1606_carry_7_), .CO(r1606_carry_8_), .S(r1606_sum_7_) );
  ADDF_X1M_A12TR r201_u1_0 ( .A(r201_a_0_), .B(r201_b_as[0]), .CI(u3_u87_z_0), 
        .CO(r201_carry_1_), .S(r201_sum_0_) );
  ADDF_X1M_A12TR r201_u1_1 ( .A(u3_u85_z_1), .B(r201_b_as[1]), .CI(
        r201_carry_1_), .CO(r201_carry_2_), .S(r201_sum_1_) );
  ADDF_X1M_A12TR r201_u1_2 ( .A(u3_u85_z_2), .B(u3_u87_z_0), .CI(r201_carry_2_), .CO(r201_carry_3_), .S(r201_sum_2_) );
  ADDF_X1M_A12TR r201_u1_3 ( .A(u3_u85_z_3), .B(u3_u87_z_0), .CI(r201_carry_3_), .CO(r201_carry_4_), .S(r201_sum_3_) );
  ADDF_X1M_A12TR r201_u1_4 ( .A(u3_u85_z_4), .B(u3_u87_z_0), .CI(r201_carry_4_), .CO(r201_carry_5_), .S(r201_sum_4_) );
  ADDF_X1M_A12TR r201_u1_5 ( .A(u3_u85_z_5), .B(u3_u87_z_0), .CI(r201_carry_5_), .CO(r201_carry_6_), .S(r201_sum_5_) );
  ADDF_X1M_A12TR r201_u1_6 ( .A(u3_u85_z_6), .B(u3_u87_z_0), .CI(r201_carry_6_), .CO(r201_carry_7_), .S(r201_sum_6_) );
  ADDF_X1M_A12TR r201_u1_7 ( .A(u3_u85_z_7), .B(u3_u87_z_0), .CI(r201_carry_7_), .CO(r201_carry_8_), .S(r201_sum_7_) );
  ADDF_X1M_A12TR r201_u1_8 ( .A(u3_u85_z_8), .B(u3_u87_z_0), .CI(r201_carry_8_), .CO(r201_carry_9_), .S(r201_sum_8_) );
  ADDF_X1M_A12TR r201_u1_9 ( .A(r201_a_9_), .B(u3_u87_z_0), .CI(r201_carry_9_), 
        .CO(r201_carry_10_), .S(r201_sum_9_) );
  ADDF_X1M_A12TR r201_u1_10 ( .A(r201_a_10_), .B(u3_u87_z_0), .CI(
        r201_carry_10_), .CO(r201_carry_11_), .S(r201_sum_10_) );
  ADDF_X1M_A12TR r201_u1_11 ( .A(r201_a_11_), .B(u3_u87_z_0), .CI(
        r201_carry_11_), .CO(r201_carry_12_), .S(r201_sum_11_) );
  ADDF_X1M_A12TR r201_u1_12 ( .A(r201_a_12_), .B(u3_u87_z_0), .CI(
        r201_carry_12_), .CO(r201_carry_13_), .S(r201_sum_12_) );
  ADDF_X1M_A12TR r201_u1_13 ( .A(r201_a_13_), .B(u3_u87_z_0), .CI(
        r201_carry_13_), .CO(r201_carry_14_), .S(r201_sum_13_) );
  ADDF_X1M_A12TR r201_u1_14 ( .A(r201_a_14_), .B(u3_u87_z_0), .CI(
        r201_carry_14_), .CO(r201_carry_15_), .S(r201_sum_14_) );
  ADDF_X1M_A12TR r201_u1_15 ( .A(r201_a_15_), .B(u3_u87_z_0), .CI(
        r201_carry_15_), .CO(), .S(r201_sum_15_) );
  ADDF_X1M_A12TR r194_u1_1 ( .A(u3_u88_z_1), .B(r194_b_as[1]), .CI(
        r194_carry_1_), .CO(r194_carry_2_), .S(r194_sum_1_) );
  DFFQ_X1M_A12TR writeio_reg ( .D(n2723), .CK(clock), .Q(writeio) );
  DFFQ_X1M_A12TR addr_reg_15_ ( .D(n2516), .CK(clock), .Q(addr[15]) );
  DFFQ_X1M_A12TR addr_reg_14_ ( .D(n2515), .CK(clock), .Q(addr[14]) );
  DFFQ_X1M_A12TR addr_reg_13_ ( .D(n2514), .CK(clock), .Q(addr[13]) );
  DFFQ_X1M_A12TR addr_reg_12_ ( .D(n2513), .CK(clock), .Q(addr[12]) );
  DFFQ_X1M_A12TR addr_reg_11_ ( .D(n2512), .CK(clock), .Q(addr[11]) );
  DFFQ_X1M_A12TR addr_reg_10_ ( .D(n2511), .CK(clock), .Q(addr[10]) );
  DFFQ_X1M_A12TR addr_reg_9_ ( .D(n2510), .CK(clock), .Q(addr[9]) );
  DFFQ_X1M_A12TR addr_reg_8_ ( .D(n2509), .CK(clock), .Q(addr[8]) );
  DFFQ_X1M_A12TR addr_reg_7_ ( .D(n2508), .CK(clock), .Q(addr[7]) );
  DFFQ_X1M_A12TR addr_reg_6_ ( .D(n2507), .CK(clock), .Q(addr[6]) );
  DFFQ_X1M_A12TR addr_reg_5_ ( .D(n2506), .CK(clock), .Q(addr[5]) );
  DFFQ_X1M_A12TR addr_reg_4_ ( .D(n2505), .CK(clock), .Q(addr[4]) );
  DFFQ_X1M_A12TR addr_reg_3_ ( .D(n2504), .CK(clock), .Q(addr[3]) );
  DFFQ_X1M_A12TR addr_reg_2_ ( .D(n2503), .CK(clock), .Q(addr[2]) );
  DFFQ_X1M_A12TR addr_reg_1_ ( .D(n2502), .CK(clock), .Q(addr[1]) );
  DFFQ_X1M_A12TR addr_reg_0_ ( .D(n2501), .CK(clock), .Q(addr[0]) );
  DFFQ_X1M_A12TR readio_reg ( .D(n2500), .CK(clock), .Q(readio) );
  DFFQ_X1M_A12TR writemem_reg ( .D(n2724), .CK(clock), .Q(writemem) );
  DFFQ_X1M_A12TR alucin_reg ( .D(n2692), .CK(clock), .Q(alucin) );
  DFFQ_X1M_A12TR raddrhold_reg_8_ ( .D(n26581), .CK(clock), .Q(raddrhold[8])
         );
  DFFQ_X1M_A12TR raddrhold_reg_9_ ( .D(n2657), .CK(clock), .Q(raddrhold[9]) );
  DFFQ_X1M_A12TR raddrhold_reg_10_ ( .D(n2656), .CK(clock), .Q(raddrhold[10])
         );
  DFFQ_X1M_A12TR raddrhold_reg_11_ ( .D(n2655), .CK(clock), .Q(raddrhold[11])
         );
  DFFQ_X1M_A12TR raddrhold_reg_13_ ( .D(n2653), .CK(clock), .Q(raddrhold[13])
         );
  DFFQ_X1M_A12TR raddrhold_reg_14_ ( .D(n2652), .CK(clock), .Q(raddrhold[14])
         );
  DFFQ_X1M_A12TR raddrhold_reg_12_ ( .D(n2654), .CK(clock), .Q(raddrhold[12])
         );
  DFFQ_X1M_A12TR raddrhold_reg_15_ ( .D(n2736), .CK(clock), .Q(raddrhold[15])
         );
  DFFQ_X1M_A12TR auxcar_reg ( .D(n2639), .CK(clock), .Q(auxcar) );
  DFFQ_X1M_A12TR eienb_reg ( .D(n2683), .CK(clock), .Q(eienb) );
  DFFQ_X1M_A12TR ei_reg ( .D(n2682), .CK(clock), .Q(ei) );
  DFFQ_X1M_A12TR sign_reg ( .D(n2641), .CK(clock), .Q(sign) );
  DFFQ_X1M_A12TR raddrhold_reg_1_ ( .D(n26651), .CK(clock), .Q(raddrhold[1])
         );
  DFFQ_X1M_A12TR raddrhold_reg_2_ ( .D(n26641), .CK(clock), .Q(raddrhold[2])
         );
  DFFQ_X1M_A12TR raddrhold_reg_3_ ( .D(n26631), .CK(clock), .Q(raddrhold[3])
         );
  DFFQ_X1M_A12TR raddrhold_reg_4_ ( .D(n26621), .CK(clock), .Q(raddrhold[4])
         );
  DFFQ_X1M_A12TR raddrhold_reg_5_ ( .D(n26611), .CK(clock), .Q(raddrhold[5])
         );
  DFFQ_X1M_A12TR raddrhold_reg_6_ ( .D(n26601), .CK(clock), .Q(raddrhold[6])
         );
  DFFQ_X1M_A12TR raddrhold_reg_7_ ( .D(n26591), .CK(clock), .Q(raddrhold[7])
         );
  DFFQ_X1M_A12TR intcyc_reg ( .D(n2681), .CK(clock), .Q(intcyc) );
  DFFQ_X1M_A12TR raddrhold_reg_0_ ( .D(n26661), .CK(clock), .Q(raddrhold[0])
         );
  DFFQ_X1M_A12TR popdes_reg_1_ ( .D(n2684), .CK(clock), .Q(popdes[1]) );
  DFFQ_X1M_A12TR popdes_reg_0_ ( .D(n2685), .CK(clock), .Q(popdes[0]) );
  DFFQ_X1M_A12TR opcode_reg_6_ ( .D(n2694), .CK(clock), .Q(opcode[6]) );
  DFFQ_X1M_A12TR opcode_reg_7_ ( .D(n2693), .CK(clock), .Q(opcode[7]) );
  DFFQ_X1M_A12TR regfil_reg_6__6_ ( .D(n2617), .CK(clock), .Q(regfil_6__6_) );
  DFFQ_X1M_A12TR regfil_reg_6__4_ ( .D(n2619), .CK(clock), .Q(regfil_6__4_) );
  DFFQ_X1M_A12TR regfil_reg_6__0_ ( .D(n2623), .CK(clock), .Q(regfil_6__0_) );
  DFFQ_X1M_A12TR regfil_reg_6__7_ ( .D(n2616), .CK(clock), .Q(regfil_6__7_) );
  DFFQ_X1M_A12TR regfil_reg_6__5_ ( .D(n2618), .CK(clock), .Q(regfil_6__5_) );
  DFFQ_X1M_A12TR regfil_reg_6__3_ ( .D(n2620), .CK(clock), .Q(regfil_6__3_) );
  DFFQ_X1M_A12TR regfil_reg_6__2_ ( .D(n2621), .CK(clock), .Q(regfil_6__2_) );
  DFFQ_X1M_A12TR regfil_reg_6__1_ ( .D(n2622), .CK(clock), .Q(regfil_6__1_) );
  DFFQ_X1M_A12TR sp_reg_0_ ( .D(n2554), .CK(clock), .Q(n31370) );
  DFFQ_X1M_A12TR carry_reg ( .D(n2733), .CK(clock), .Q(carry) );
  DFFQ_X1M_A12TR zero_reg ( .D(n2642), .CK(clock), .Q(zero) );
  DFFQ_X1M_A12TR parity_reg ( .D(n2643), .CK(clock), .Q(parity) );
  DFFQ_X1M_A12TR regd_reg_1_ ( .D(n2687), .CK(clock), .Q(regd[1]) );
  DFFQ_X1M_A12TR regd_reg_0_ ( .D(n2688), .CK(clock), .Q(regd[0]) );
  DFFQ_X1M_A12TR rdatahold2_reg_0_ ( .D(n2719), .CK(clock), .Q(rdatahold2[0])
         );
  DFFQ_X1M_A12TR aluoprb_reg_0_ ( .D(n2651), .CK(clock), .Q(aluoprb_0_) );
  DFFQ_X1M_A12TR pc_reg_15_ ( .D(n2735), .CK(clock), .Q(pc[15]) );
  DFFQ_X1M_A12TR datao_reg_0_ ( .D(n2721), .CK(clock), .Q(datao[0]) );
  DFFQ_X1M_A12TR datao_reg_4_ ( .D(n2709), .CK(clock), .Q(datao[4]) );
  DFFQ_X1M_A12TR datao_reg_7_ ( .D(n2739), .CK(clock), .Q(datao[7]) );
  DFFQ_X1M_A12TR datao_reg_6_ ( .D(n2703), .CK(clock), .Q(datao[6]) );
  DFFQ_X1M_A12TR datao_reg_1_ ( .D(n2718), .CK(clock), .Q(datao[1]) );
  DFFQ_X1M_A12TR datao_reg_2_ ( .D(n2715), .CK(clock), .Q(datao[2]) );
  DFFQ_X1M_A12TR datao_reg_3_ ( .D(n2712), .CK(clock), .Q(datao[3]) );
  DFFQ_X1M_A12TR datao_reg_5_ ( .D(n2706), .CK(clock), .Q(datao[5]) );
  DFFQ_X1M_A12TR regd_reg_2_ ( .D(n2686), .CK(clock), .Q(regd[2]) );
  DFFQ_X1M_A12TR rdatahold2_reg_5_ ( .D(n2704), .CK(clock), .Q(rdatahold2[5])
         );
  DFFQ_X1M_A12TR rdatahold2_reg_3_ ( .D(n2710), .CK(clock), .Q(rdatahold2[3])
         );
  DFFQ_X1M_A12TR rdatahold2_reg_1_ ( .D(n2716), .CK(clock), .Q(rdatahold2[1])
         );
  DFFQ_X1M_A12TR regfil_reg_1__0_ ( .D(n2584), .CK(clock), .Q(n1167) );
  DFFQ_X1M_A12TR regfil_reg_7__4_ ( .D(n2634), .CK(clock), .Q(n1105) );
  DFFQ_X1M_A12TR regfil_reg_1__1_ ( .D(n2583), .CK(clock), .Q(n1168) );
  DFFQ_X1M_A12TR regfil_reg_1__5_ ( .D(n2579), .CK(clock), .Q(n1172) );
  DFFQ_X1M_A12TR regfil_reg_1__3_ ( .D(n2581), .CK(clock), .Q(n1170) );
  DFFQ_X1M_A12TR regfil_reg_1__6_ ( .D(n2578), .CK(clock), .Q(n1173) );
  DFFQ_X1M_A12TR regfil_reg_1__4_ ( .D(n2580), .CK(clock), .Q(n1171) );
  DFFQ_X1M_A12TR regfil_reg_1__2_ ( .D(n2582), .CK(clock), .Q(n1169) );
  DFFQ_X1M_A12TR rdatahold2_reg_7_ ( .D(n2725), .CK(clock), .Q(rdatahold2[7])
         );
  DFFQ_X1M_A12TR regfil_reg_1__7_ ( .D(n2640), .CK(clock), .Q(n1174) );
  DFFQ_X1M_A12TR rdatahold2_reg_4_ ( .D(n2707), .CK(clock), .Q(rdatahold2[4])
         );
  DFFQ_X1M_A12TR regfil_reg_0__0_ ( .D(n2577), .CK(clock), .Q(n1175) );
  DFFQ_X1M_A12TR regfil_reg_7__7_ ( .D(n2738), .CK(clock), .Q(n1108) );
  DFFQ_X1M_A12TR regfil_reg_7__3_ ( .D(n2635), .CK(clock), .Q(n1104) );
  DFFQ_X1M_A12TR regfil_reg_0__7_ ( .D(n2737), .CK(clock), .Q(n1182) );
  DFFQ_X1M_A12TR regfil_reg_0__4_ ( .D(n2573), .CK(clock), .Q(n1179) );
  DFFQ_X1M_A12TR regfil_reg_0__5_ ( .D(n2572), .CK(clock), .Q(n1180) );
  DFFQ_X1M_A12TR regfil_reg_0__3_ ( .D(n2574), .CK(clock), .Q(n1178) );
  DFFQ_X1M_A12TR regfil_reg_0__2_ ( .D(n2575), .CK(clock), .Q(n1177) );
  DFFQ_X1M_A12TR regfil_reg_0__1_ ( .D(n2576), .CK(clock), .Q(n1176) );
  DFFQ_X1M_A12TR regfil_reg_0__6_ ( .D(n2571), .CK(clock), .Q(n1181) );
  DFFQ_X1M_A12TR regfil_reg_7__6_ ( .D(n2632), .CK(clock), .Q(n1107) );
  DFFQ_X1M_A12TR regfil_reg_7__2_ ( .D(n2636), .CK(clock), .Q(n1103) );
  DFFQ_X1M_A12TR rdatahold2_reg_6_ ( .D(n2701), .CK(clock), .Q(rdatahold2[6])
         );
  DFFQ_X1M_A12TR rdatahold2_reg_2_ ( .D(n2713), .CK(clock), .Q(rdatahold2[2])
         );
  DFFQ_X1M_A12TR regfil_reg_7__5_ ( .D(n2633), .CK(clock), .Q(n1106) );
  DFFQ_X1M_A12TR regfil_reg_7__1_ ( .D(n2637), .CK(clock), .Q(n1102) );
  DFFQ_X1M_A12TR regfil_reg_7__0_ ( .D(n2638), .CK(clock), .Q(regfil_7__0_) );
  DFFQ_X1M_A12TR aluopra_reg_7_ ( .D(n2624), .CK(clock), .Q(aluopra[7]) );
  DFFQ_X1M_A12TR aluopra_reg_5_ ( .D(n2626), .CK(clock), .Q(aluopra[5]) );
  DFFQ_X1M_A12TR aluopra_reg_6_ ( .D(n2625), .CK(clock), .Q(aluopra[6]) );
  DFFQ_X1M_A12TR aluopra_reg_4_ ( .D(n2627), .CK(clock), .Q(aluopra[4]) );
  DFFQ_X1M_A12TR regfil_reg_2__0_ ( .D(n2591), .CK(clock), .Q(regfil_2__0_) );
  DFFQ_X1M_A12TR regfil_reg_2__4_ ( .D(n2587), .CK(clock), .Q(regfil_2__4_) );
  DFFQ_X1M_A12TR regfil_reg_2__7_ ( .D(n2734), .CK(clock), .Q(regfil_2__7_) );
  DFFQ_X1M_A12TR regfil_reg_2__5_ ( .D(n2586), .CK(clock), .Q(regfil_2__5_) );
  DFFQ_X1M_A12TR regfil_reg_2__3_ ( .D(n2588), .CK(clock), .Q(regfil_2__3_) );
  DFFQ_X1M_A12TR regfil_reg_2__2_ ( .D(n2589), .CK(clock), .Q(regfil_2__2_) );
  DFFQ_X1M_A12TR regfil_reg_2__1_ ( .D(n2590), .CK(clock), .Q(regfil_2__1_) );
  DFFQ_X1M_A12TR regfil_reg_2__6_ ( .D(n2585), .CK(clock), .Q(regfil_2__6_) );
  DFFQ_X1M_A12TR regfil_reg_3__5_ ( .D(n2594), .CK(clock), .Q(n1662) );
  DFFQ_X1M_A12TR regfil_reg_3__3_ ( .D(n2596), .CK(clock), .Q(n1660) );
  DFFQ_X1M_A12TR regfil_reg_3__0_ ( .D(n2599), .CK(clock), .Q(n1657) );
  DFFQ_X1M_A12TR regfil_reg_3__6_ ( .D(n2593), .CK(clock), .Q(n1663) );
  DFFQ_X1M_A12TR regfil_reg_3__4_ ( .D(n2595), .CK(clock), .Q(n1661) );
  DFFQ_X1M_A12TR regfil_reg_3__2_ ( .D(n2597), .CK(clock), .Q(n1659) );
  DFFQ_X1M_A12TR regfil_reg_3__7_ ( .D(n2592), .CK(clock), .Q(n1664) );
  DFFQ_X1M_A12TR regfil_reg_3__1_ ( .D(n2598), .CK(clock), .Q(n1658) );
  DFFQ_X1M_A12TR rdatahold_reg_5_ ( .D(n2705), .CK(clock), .Q(rdatahold[5]) );
  DFFQ_X1M_A12TR rdatahold_reg_3_ ( .D(n2711), .CK(clock), .Q(rdatahold[3]) );
  DFFQ_X1M_A12TR state_reg_3_ ( .D(n2728), .CK(clock), .Q(state[3]) );
  DFFQ_X1M_A12TR pc_reg_12_ ( .D(n2558), .CK(clock), .Q(pc[12]) );
  DFFQ_X1M_A12TR pc_reg_13_ ( .D(n2557), .CK(clock), .Q(pc[13]) );
  DFFQ_X1M_A12TR pc_reg_11_ ( .D(n2559), .CK(clock), .Q(pc[11]) );
  DFFQ_X1M_A12TR pc_reg_10_ ( .D(n2560), .CK(clock), .Q(pc[10]) );
  DFFQ_X1M_A12TR pc_reg_9_ ( .D(n2561), .CK(clock), .Q(pc[9]) );
  DFFQ_X1M_A12TR pc_reg_14_ ( .D(n2556), .CK(clock), .Q(pc[14]) );
  DFFQ_X1M_A12TR pc_reg_8_ ( .D(n2562), .CK(clock), .Q(pc[8]) );
  DFFQ_X1M_A12TR regfil_reg_4__4_ ( .D(n2603), .CK(clock), .Q(n1162) );
  DFFQ_X1M_A12TR regfil_reg_4__0_ ( .D(n2607), .CK(clock), .Q(n1158) );
  DFFQ_X1M_A12TR regfil_reg_4__7_ ( .D(n2600), .CK(clock), .Q(n1165) );
  DFFQ_X1M_A12TR regfil_reg_4__5_ ( .D(n2602), .CK(clock), .Q(n1163) );
  DFFQ_X1M_A12TR regfil_reg_4__3_ ( .D(n2604), .CK(clock), .Q(n1161) );
  DFFQ_X1M_A12TR regfil_reg_4__2_ ( .D(n2605), .CK(clock), .Q(n1160) );
  DFFQ_X1M_A12TR regfil_reg_4__1_ ( .D(n2606), .CK(clock), .Q(n1159) );
  DFFQ_X1M_A12TR regfil_reg_4__6_ ( .D(n2601), .CK(clock), .Q(n1164) );
  DFFQ_X1M_A12TR rdatahold_reg_0_ ( .D(n2720), .CK(clock), .Q(rdatahold[0]) );
  DFFQ_X1M_A12TR rdatahold_reg_4_ ( .D(n2708), .CK(clock), .Q(rdatahold[4]) );
  DFFQ_X1M_A12TR rdatahold_reg_6_ ( .D(n2702), .CK(clock), .Q(rdatahold[6]) );
  DFFQ_X1M_A12TR rdatahold_reg_2_ ( .D(n2714), .CK(clock), .Q(rdatahold[2]) );
  DFFQ_X1M_A12TR rdatahold_reg_1_ ( .D(n2717), .CK(clock), .Q(rdatahold[1]) );
  DFFQ_X1M_A12TR rdatahold_reg_7_ ( .D(n2726), .CK(clock), .Q(rdatahold[7]) );
  DFFQ_X1M_A12TR aluopra_reg_2_ ( .D(n2629), .CK(clock), .Q(aluopra[2]) );
  DFFQ_X1M_A12TR pc_reg_6_ ( .D(n2564), .CK(clock), .Q(pc[6]) );
  DFFQ_X1M_A12TR pc_reg_7_ ( .D(n2563), .CK(clock), .Q(pc[7]) );
  DFFQ_X1M_A12TR pc_reg_2_ ( .D(n2568), .CK(clock), .Q(pc[2]) );
  DFFQ_X1M_A12TR pc_reg_3_ ( .D(n2567), .CK(clock), .Q(pc[3]) );
  DFFQ_X1M_A12TR pc_reg_5_ ( .D(n2565), .CK(clock), .Q(pc[5]) );
  DFFQ_X1M_A12TR regfil_reg_5__1_ ( .D(n2614), .CK(clock), .Q(n1151) );
  DFFQ_X1M_A12TR state_reg_5_ ( .D(n2732), .CK(clock), .Q(state[5]) );
  DFFQ_X1M_A12TR pc_reg_1_ ( .D(n2569), .CK(clock), .Q(pc[1]) );
  DFFQ_X1M_A12TR regfil_reg_5__5_ ( .D(n2610), .CK(clock), .Q(n1155) );
  DFFQ_X1M_A12TR regfil_reg_5__3_ ( .D(n2612), .CK(clock), .Q(n1153) );
  DFFQ_X1M_A12TR regfil_reg_5__0_ ( .D(n2615), .CK(clock), .Q(n1150) );
  DFFQ_X1M_A12TR aluopra_reg_0_ ( .D(n2631), .CK(clock), .Q(aluopra[0]) );
  DFFQ_X1M_A12TR pc_reg_4_ ( .D(n2566), .CK(clock), .Q(pc[4]) );
  DFFQ_X1M_A12TR regfil_reg_5__6_ ( .D(n2609), .CK(clock), .Q(n1156) );
  DFFQ_X1M_A12TR regfil_reg_5__2_ ( .D(n2613), .CK(clock), .Q(n1152) );
  DFFQ_X1M_A12TR regfil_reg_5__7_ ( .D(n2608), .CK(clock), .Q(n1157) );
  DFFQ_X1M_A12TR regfil_reg_5__4_ ( .D(n2611), .CK(clock), .Q(n1154) );
  DFFQN_X1M_A12TR wdatahold2_reg_0_ ( .D(n2741), .CK(clock), .QN(n2498) );
  DFFQN_X1M_A12TR wdatahold2_reg_7_ ( .D(n2517), .CK(clock), .QN(n2491) );
  DFFQN_X1M_A12TR wdatahold2_reg_1_ ( .D(n2523), .CK(clock), .QN(n2497) );
  DFFQN_X1M_A12TR wdatahold2_reg_5_ ( .D(n2519), .CK(clock), .QN(n2493) );
  DFFQN_X1M_A12TR wdatahold2_reg_3_ ( .D(n2521), .CK(clock), .QN(n2495) );
  DFFQN_X1M_A12TR wdatahold2_reg_2_ ( .D(n2522), .CK(clock), .QN(n2496) );
  DFFQN_X1M_A12TR wdatahold2_reg_6_ ( .D(n2518), .CK(clock), .QN(n2492) );
  DFFQN_X1M_A12TR wdatahold2_reg_4_ ( .D(n2520), .CK(clock), .QN(n2494) );
  DFFQ_X1M_A12TR pc_reg_0_ ( .D(n2570), .CK(clock), .Q(pc[0]) );
  DFFQ_X1M_A12TR aluopra_reg_3_ ( .D(n2628), .CK(clock), .Q(aluopra[3]) );
  DFFQ_X1M_A12TR aluopra_reg_1_ ( .D(n2630), .CK(clock), .Q(aluopra[1]) );
  DFFQ_X1M_A12TR sp_reg_15_ ( .D(n2555), .CK(clock), .Q(sp[15]) );
  DFFQ_X1M_A12TR state_reg_2_ ( .D(n2729), .CK(clock), .Q(state[2]) );
  DFFQN_X1M_A12TR aluoprb_reg_6_ ( .D(n2645), .CK(clock), .QN(n2464) );
  DFFQN_X1M_A12TR aluoprb_reg_4_ ( .D(n2647), .CK(clock), .QN(n2463) );
  DFFQN_X1M_A12TR aluoprb_reg_7_ ( .D(n2644), .CK(clock), .QN(n2462) );
  DFFQN_X1M_A12TR aluoprb_reg_5_ ( .D(n2646), .CK(clock), .QN(n2460) );
  DFFQN_X1M_A12TR aluoprb_reg_3_ ( .D(n2648), .CK(clock), .QN(n2459) );
  DFFQN_X1M_A12TR aluoprb_reg_2_ ( .D(n2649), .CK(clock), .QN(n2458) );
  DFFQN_X1M_A12TR aluoprb_reg_1_ ( .D(n2650), .CK(clock), .QN(n2457) );
  DFFQN_X1M_A12TR waddrhold_reg_15_ ( .D(n2524), .CK(clock), .QN(n2467) );
  DFFQN_X1M_A12TR waddrhold_reg_1_ ( .D(n2538), .CK(clock), .QN(n2481) );
  DFFQN_X1M_A12TR waddrhold_reg_2_ ( .D(n2537), .CK(clock), .QN(n2480) );
  DFFQN_X1M_A12TR waddrhold_reg_3_ ( .D(n2536), .CK(clock), .QN(n2479) );
  DFFQN_X1M_A12TR waddrhold_reg_4_ ( .D(n2535), .CK(clock), .QN(n2478) );
  DFFQN_X1M_A12TR waddrhold_reg_5_ ( .D(n2534), .CK(clock), .QN(n2477) );
  DFFQN_X1M_A12TR waddrhold_reg_6_ ( .D(n2533), .CK(clock), .QN(n2476) );
  DFFQN_X1M_A12TR waddrhold_reg_7_ ( .D(n2532), .CK(clock), .QN(n2475) );
  DFFQN_X1M_A12TR waddrhold_reg_8_ ( .D(n2531), .CK(clock), .QN(n2474) );
  DFFQN_X1M_A12TR waddrhold_reg_9_ ( .D(n2530), .CK(clock), .QN(n2473) );
  DFFQN_X1M_A12TR waddrhold_reg_10_ ( .D(n2529), .CK(clock), .QN(n2472) );
  DFFQN_X1M_A12TR waddrhold_reg_11_ ( .D(n2528), .CK(clock), .QN(n2471) );
  DFFQN_X1M_A12TR waddrhold_reg_12_ ( .D(n2527), .CK(clock), .QN(n2470) );
  DFFQN_X1M_A12TR waddrhold_reg_13_ ( .D(n2526), .CK(clock), .QN(n2469) );
  DFFQN_X1M_A12TR waddrhold_reg_14_ ( .D(n2525), .CK(clock), .QN(n2468) );
  DFFQN_X1M_A12TR wdatahold_reg_0_ ( .D(n2673), .CK(clock), .QN(n2490) );
  DFFQN_X1M_A12TR wdatahold_reg_4_ ( .D(n26691), .CK(clock), .QN(n2486) );
  DFFQN_X1M_A12TR wdatahold_reg_7_ ( .D(n2740), .CK(clock), .QN(n2483) );
  DFFQN_X1M_A12TR wdatahold_reg_1_ ( .D(n26721), .CK(clock), .QN(n2489) );
  DFFQN_X1M_A12TR wdatahold_reg_2_ ( .D(n26711), .CK(clock), .QN(n2488) );
  DFFQN_X1M_A12TR wdatahold_reg_3_ ( .D(n26701), .CK(clock), .QN(n2487) );
  DFFQN_X1M_A12TR wdatahold_reg_5_ ( .D(n26681), .CK(clock), .QN(n2485) );
  DFFQN_X1M_A12TR wdatahold_reg_6_ ( .D(n26671), .CK(clock), .QN(n2484) );
  DFFQ_X1M_A12TR statesel_reg_5_ ( .D(n2679), .CK(clock), .Q(statesel[5]) );
  DFFQN_X1M_A12TR dataeno_reg ( .D(n2722), .CK(clock), .QN(n2465) );
  DFFQN_X1M_A12TR readmem_reg ( .D(n2680), .CK(clock), .QN(n2461) );
  DFFQN_X1M_A12TR inta_reg ( .D(n2499), .CK(clock), .QN(n2456) );
  DFFQ_X1M_A12TR statesel_reg_2_ ( .D(n2676), .CK(clock), .Q(statesel[2]) );
  DFFQ_X1M_A12TR sp_reg_1_ ( .D(n2553), .CK(clock), .Q(sp[1]) );
  DFFQN_X1M_A12TR waddrhold_reg_0_ ( .D(n2539), .CK(clock), .QN(n2482) );
  DFFQ_X1M_A12TR sp_reg_14_ ( .D(n2540), .CK(clock), .Q(sp[14]) );
  DFFQ_X1M_A12TR sp_reg_13_ ( .D(n2541), .CK(clock), .Q(sp[13]) );
  DFFQ_X1M_A12TR sp_reg_2_ ( .D(n2552), .CK(clock), .Q(sp[2]) );
  DFFQ_X1M_A12TR sp_reg_3_ ( .D(n2551), .CK(clock), .Q(sp[3]) );
  DFFQ_X1M_A12TR sp_reg_4_ ( .D(n2550), .CK(clock), .Q(sp[4]) );
  DFFQ_X1M_A12TR sp_reg_5_ ( .D(n2549), .CK(clock), .Q(sp[5]) );
  DFFQ_X1M_A12TR sp_reg_6_ ( .D(n2548), .CK(clock), .Q(sp[6]) );
  DFFQ_X1M_A12TR sp_reg_7_ ( .D(n2547), .CK(clock), .Q(sp[7]) );
  DFFQ_X1M_A12TR sp_reg_8_ ( .D(n2546), .CK(clock), .Q(sp[8]) );
  DFFQ_X1M_A12TR sp_reg_9_ ( .D(n2545), .CK(clock), .Q(sp[9]) );
  DFFQ_X1M_A12TR sp_reg_10_ ( .D(n2544), .CK(clock), .Q(sp[10]) );
  DFFQ_X1M_A12TR sp_reg_11_ ( .D(n2543), .CK(clock), .Q(sp[11]) );
  DFFQ_X1M_A12TR sp_reg_12_ ( .D(n2542), .CK(clock), .Q(sp[12]) );
  DFFQ_X1M_A12TR statesel_reg_3_ ( .D(n2675), .CK(clock), .Q(statesel[3]) );
  DFFQ_X1M_A12TR state_reg_4_ ( .D(n2727), .CK(clock), .Q(state[4]) );
  DFFQ_X1M_A12TR statesel_reg_4_ ( .D(n2674), .CK(clock), .Q(statesel[4]) );
  DFFQ_X1M_A12TR statesel_reg_1_ ( .D(n2677), .CK(clock), .Q(statesel[1]) );
  DFFQ_X1M_A12TR statesel_reg_0_ ( .D(n2678), .CK(clock), .Q(statesel[0]) );
  BUFZ_X1M_A12TR data_tri_0_ ( .A(datao[0]), .OE(n4310), .Y(data_out[0]) );
  BUFZ_X1M_A12TR data_tri_1_ ( .A(datao[1]), .OE(n4310), .Y(data_out[1]) );
  BUFZ_X1M_A12TR data_tri_2_ ( .A(datao[2]), .OE(n4310), .Y(data_out[2]) );
  BUFZ_X1M_A12TR data_tri_3_ ( .A(datao[3]), .OE(n4310), .Y(data_out[3]) );
  BUFZ_X1M_A12TR data_tri_4_ ( .A(datao[4]), .OE(n4310), .Y(data_out[4]) );
  BUFZ_X1M_A12TR data_tri_5_ ( .A(datao[5]), .OE(n4310), .Y(data_out[5]) );
  BUFZ_X1M_A12TR data_tri_6_ ( .A(datao[6]), .OE(n4310), .Y(data_out[6]) );
  BUFZ_X1M_A12TR data_tri_7_ ( .A(datao[7]), .OE(n4310), .Y(data_out[7]) );
  DFFQ_X1M_A12TR alusel_reg_0_ ( .D(n2691), .CK(clock), .Q(alusel[0]) );
  DFFQ_X1M_A12TR alusel_reg_1_ ( .D(n2690), .CK(clock), .Q(alusel[1]) );
  DFFQ_X1M_A12TR state_reg_0_ ( .D(n2731), .CK(clock), .Q(state[0]) );
  DFFQ_X1M_A12TR state_reg_1_ ( .D(n2730), .CK(clock), .Q(u3_u93_z_6) );
  DFFQ_X1M_A12TR alusel_reg_2_ ( .D(n2689), .CK(clock), .Q(alusel[2]) );
  DFFQ_X1M_A12TR opcode_reg_2_ ( .D(n2698), .CK(clock), .Q(n235) );
  DFFQ_X1M_A12TR opcode_reg_5_ ( .D(n2695), .CK(clock), .Q(n237) );
  DFFQ_X1M_A12TR opcode_reg_0_ ( .D(n2700), .CK(clock), .Q(n233) );
  DFFQ_X1M_A12TR opcode_reg_4_ ( .D(n2696), .CK(clock), .Q(n46) );
  DFFQ_X1M_A12TR opcode_reg_1_ ( .D(n2699), .CK(clock), .Q(n234) );
  DFFQ_X1M_A12TR opcode_reg_3_ ( .D(n2697), .CK(clock), .Q(n236) );
  XOR3_X0P5M_A12TR r194_u1_15 ( .A(u3_u88_z_15), .B(n2742), .C(r194_carry_15_), 
        .Y(r194_sum_15_) );
  ADDF_X1M_A12TR r194_u1_0 ( .A(u3_u88_z_0), .B(r194_b_as[0]), .CI(n2742), 
        .CO(r194_carry_1_), .S(r194_sum_0_) );
  ADDF_X1M_A12TR r194_u1_8 ( .A(u3_u88_z_8), .B(n2742), .CI(r194_carry_8_), 
        .CO(r194_carry_9_), .S(r194_sum_8_) );
  ADDF_X1M_A12TR r194_u1_12 ( .A(u3_u88_z_12), .B(n2742), .CI(r194_carry_12_), 
        .CO(r194_carry_13_), .S(r194_sum_12_) );
  ADDF_X1M_A12TR r194_u1_13 ( .A(u3_u88_z_13), .B(n2742), .CI(r194_carry_13_), 
        .CO(r194_carry_14_), .S(r194_sum_13_) );
  ADDF_X1M_A12TR r194_u1_11 ( .A(u3_u88_z_11), .B(n2742), .CI(r194_carry_11_), 
        .CO(r194_carry_12_), .S(r194_sum_11_) );
  ADDF_X1M_A12TR r194_u1_10 ( .A(u3_u88_z_10), .B(n2742), .CI(r194_carry_10_), 
        .CO(r194_carry_11_), .S(r194_sum_10_) );
  ADDF_X1M_A12TR r194_u1_9 ( .A(u3_u88_z_9), .B(n2742), .CI(r194_carry_9_), 
        .CO(r194_carry_10_), .S(r194_sum_9_) );
  ADDF_X1M_A12TR r194_u1_14 ( .A(u3_u88_z_14), .B(n2742), .CI(r194_carry_14_), 
        .CO(r194_carry_15_), .S(r194_sum_14_) );
  ADDF_X1M_A12TR r194_u1_6 ( .A(u3_u88_z_6), .B(n2742), .CI(r194_carry_6_), 
        .CO(r194_carry_7_), .S(r194_sum_6_) );
  ADDF_X1M_A12TR r194_u1_7 ( .A(u3_u88_z_7), .B(n2742), .CI(r194_carry_7_), 
        .CO(r194_carry_8_), .S(r194_sum_7_) );
  ADDF_X1M_A12TR r194_u1_2 ( .A(u3_u88_z_2), .B(n2742), .CI(r194_carry_2_), 
        .CO(r194_carry_3_), .S(r194_sum_2_) );
  ADDF_X1M_A12TR r194_u1_3 ( .A(u3_u88_z_3), .B(n2742), .CI(r194_carry_3_), 
        .CO(r194_carry_4_), .S(r194_sum_3_) );
  ADDF_X1M_A12TR r194_u1_5 ( .A(u3_u88_z_5), .B(n2742), .CI(r194_carry_5_), 
        .CO(r194_carry_6_), .S(r194_sum_5_) );
  ADDF_X1M_A12TR r194_u1_4 ( .A(u3_u88_z_4), .B(n2742), .CI(r194_carry_4_), 
        .CO(r194_carry_5_), .S(r194_sum_4_) );
  AO21B_X1M_A12TR u1900 ( .A0(n30111), .A1(n3321), .B0N(n2823), .Y(n2742) );
  INV_X1M_A12TR u1901 ( .A(u3_u93_z_6), .Y(n2823) );
  NAND3_X2M_A12TR u1902 ( .A(n3568), .B(n3356), .C(n3191), .Y(r1298_carry_1_)
         );
  AOI211_X2M_A12TR u1903 ( .A0(n3042), .A1(n4293), .B0(n3642), .C0(n3857), .Y(
        u3_u87_z_0) );
  XOR2_X1M_A12TR u1904 ( .A(u3_u94_z_0), .B(r1606_carry_8_), .Y(r1606_sum_8_)
         );
  XOR2_X1M_A12TR u1905 ( .A(u3_u84_z_1), .B(u3_u84_z_0), .Y(r1226_sum_1_) );
  XOR2_X1M_A12TR u1906 ( .A(u3_u84_z_3), .B(n2744), .Y(r1226_sum_3_) );
  XOR2_X1M_A12TR u1907 ( .A(u3_u84_z_5), .B(n2746), .Y(r1226_sum_5_) );
  XOR2_X1M_A12TR u1908 ( .A(u3_u84_z_7), .B(n2748), .Y(r1226_sum_7_) );
  XOR2_X1M_A12TR u1909 ( .A(u3_u84_z_8), .B(n2749), .Y(r1226_sum_8_) );
  XOR2_X1M_A12TR u1910 ( .A(u3_u84_z_4), .B(n2745), .Y(r1226_sum_4_) );
  XOR2_X1M_A12TR u1911 ( .A(u3_u84_z_14), .B(n2755), .Y(r1226_sum_14_) );
  XOR2_X1M_A12TR u1912 ( .A(u3_u84_z_9), .B(n2750), .Y(r1226_sum_9_) );
  XOR2_X1M_A12TR u1913 ( .A(u3_u84_z_10), .B(n2751), .Y(r1226_sum_10_) );
  XOR2_X1M_A12TR u1914 ( .A(u3_u84_z_2), .B(n2743), .Y(r1226_sum_2_) );
  XOR2_X1M_A12TR u1915 ( .A(u3_u84_z_11), .B(n2752), .Y(r1226_sum_11_) );
  XOR2_X1M_A12TR u1916 ( .A(u3_u84_z_13), .B(n2754), .Y(r1226_sum_13_) );
  XOR2_X1M_A12TR u1917 ( .A(u3_u84_z_6), .B(n2747), .Y(r1226_sum_6_) );
  XOR2_X1M_A12TR u1918 ( .A(u3_u84_z_12), .B(n2753), .Y(r1226_sum_12_) );
  AND2_X1M_A12TR u1919 ( .A(u3_u84_z_1), .B(u3_u84_z_0), .Y(n2743) );
  AND2_X1M_A12TR u1920 ( .A(u3_u84_z_2), .B(n2743), .Y(n2744) );
  AND2_X1M_A12TR u1921 ( .A(u3_u84_z_3), .B(n2744), .Y(n2745) );
  AND2_X1M_A12TR u1922 ( .A(u3_u84_z_4), .B(n2745), .Y(n2746) );
  AND2_X1M_A12TR u1923 ( .A(u3_u84_z_5), .B(n2746), .Y(n2747) );
  AND2_X1M_A12TR u1924 ( .A(u3_u84_z_6), .B(n2747), .Y(n2748) );
  AND2_X1M_A12TR u1925 ( .A(u3_u84_z_7), .B(n2748), .Y(n2749) );
  AND2_X1M_A12TR u1926 ( .A(u3_u84_z_8), .B(n2749), .Y(n2750) );
  AND2_X1M_A12TR u1927 ( .A(u3_u84_z_9), .B(n2750), .Y(n2751) );
  AND2_X1M_A12TR u1928 ( .A(u3_u84_z_10), .B(n2751), .Y(n2752) );
  AND2_X1M_A12TR u1929 ( .A(u3_u84_z_11), .B(n2752), .Y(n2753) );
  AND2_X1M_A12TR u1930 ( .A(u3_u84_z_12), .B(n2753), .Y(n2754) );
  AND2_X1M_A12TR u1931 ( .A(u3_u84_z_13), .B(n2754), .Y(n2755) );
  XNOR2_X1M_A12TR u1932 ( .A(u3_u84_z_15), .B(n2802), .Y(r1226_sum_15_) );
  NAND2_X1M_A12TR u1933 ( .A(u3_u84_z_14), .B(n2755), .Y(n2802) );
  XOR2_X1M_A12TR u1934 ( .A(statesel[3]), .B(n2774), .Y(n35730) );
  XOR2_X1M_A12TR u1935 ( .A(statesel[1]), .B(statesel[0]), .Y(n35710) );
  XOR2_X1M_A12TR u1936 ( .A(statesel[5]), .B(n2800), .Y(n35750) );
  XOR2_X1M_A12TR u1937 ( .A(statesel[2]), .B(n2772), .Y(n35720) );
  XOR2_X1M_A12TR u1938 ( .A(statesel[4]), .B(n2773), .Y(n35740) );
  XOR2_X1M_A12TR u1939 ( .A(sp[15]), .B(n2801), .Y(n31520) );
  NOR2_X1M_A12TR u1940 ( .A(n2799), .B(sp[14]), .Y(n2801) );
  MXT2_X1M_A12TR u1941 ( .A(n2756), .B(n2757), .S0(n235), .Y(n244) );
  MXT4_X1M_A12TR u1942 ( .A(n1178), .B(regfil_2__3_), .C(n1170), .D(n1660), 
        .S0(n234), .S1(n233), .Y(n2756) );
  MXT4_X1M_A12TR u1943 ( .A(n1161), .B(regfil_6__3_), .C(n1153), .D(n1104), 
        .S0(n234), .S1(n233), .Y(n2757) );
  MXT2_X1M_A12TR u1944 ( .A(n2758), .B(n2759), .S0(n235), .Y(n242) );
  MXT4_X1M_A12TR u1945 ( .A(n1180), .B(regfil_2__5_), .C(n1172), .D(n1662), 
        .S0(n234), .S1(n233), .Y(n2758) );
  MXT4_X1M_A12TR u1946 ( .A(n1163), .B(regfil_6__5_), .C(n1155), .D(n1106), 
        .S0(n234), .S1(n233), .Y(n2759) );
  MXT2_X1M_A12TR u1947 ( .A(n2760), .B(n2761), .S0(n235), .Y(n241) );
  MXT4_X1M_A12TR u1948 ( .A(n1181), .B(regfil_2__6_), .C(n1173), .D(n1663), 
        .S0(n234), .S1(n233), .Y(n2760) );
  MXT4_X1M_A12TR u1949 ( .A(n1164), .B(regfil_6__6_), .C(n1156), .D(n1107), 
        .S0(n234), .S1(n233), .Y(n2761) );
  MXT2_X1M_A12TR u1950 ( .A(n2762), .B(n2763), .S0(n235), .Y(n246) );
  MXT4_X1M_A12TR u1951 ( .A(n1176), .B(regfil_2__1_), .C(n1168), .D(n1658), 
        .S0(n234), .S1(n233), .Y(n2762) );
  MXT4_X1M_A12TR u1952 ( .A(n1159), .B(regfil_6__1_), .C(n1151), .D(n1102), 
        .S0(n234), .S1(n233), .Y(n2763) );
  MXT2_X1M_A12TR u1953 ( .A(n2764), .B(n2765), .S0(n235), .Y(n245) );
  MXT4_X1M_A12TR u1954 ( .A(n1177), .B(regfil_2__2_), .C(n1169), .D(n1659), 
        .S0(n234), .S1(n233), .Y(n2764) );
  MXT4_X1M_A12TR u1955 ( .A(n1160), .B(regfil_6__2_), .C(n1152), .D(n1103), 
        .S0(n234), .S1(n233), .Y(n2765) );
  MXT2_X1M_A12TR u1956 ( .A(n2766), .B(n2767), .S0(n235), .Y(n247) );
  MXT4_X1M_A12TR u1957 ( .A(n1175), .B(regfil_2__0_), .C(n1167), .D(n1657), 
        .S0(n234), .S1(n233), .Y(n2766) );
  MXT4_X1M_A12TR u1958 ( .A(n1158), .B(regfil_6__0_), .C(n1150), .D(
        regfil_7__0_), .S0(n234), .S1(n233), .Y(n2767) );
  MXT2_X1M_A12TR u1959 ( .A(n2768), .B(n2769), .S0(n235), .Y(n243) );
  MXT4_X1M_A12TR u1960 ( .A(n1179), .B(regfil_2__4_), .C(n1171), .D(n1661), 
        .S0(n234), .S1(n233), .Y(n2768) );
  MXT4_X1M_A12TR u1961 ( .A(n1162), .B(regfil_6__4_), .C(n1154), .D(n1105), 
        .S0(n234), .S1(n233), .Y(n2769) );
  MXT2_X1M_A12TR u1962 ( .A(n2770), .B(n2771), .S0(n235), .Y(n240) );
  MXT4_X1M_A12TR u1963 ( .A(n1182), .B(regfil_2__7_), .C(n1174), .D(n1664), 
        .S0(n234), .S1(n233), .Y(n2770) );
  MXT4_X1M_A12TR u1964 ( .A(n1165), .B(regfil_6__7_), .C(n1157), .D(n1108), 
        .S0(n234), .S1(n233), .Y(n2771) );
  XNOR2_X1M_A12TR u1965 ( .A(sp[12]), .B(n2797), .Y(n31490) );
  XNOR2_X1M_A12TR u1966 ( .A(sp[11]), .B(n2796), .Y(n31480) );
  XNOR2_X1M_A12TR u1967 ( .A(sp[10]), .B(n2795), .Y(n31470) );
  XNOR2_X1M_A12TR u1968 ( .A(sp[9]), .B(n2794), .Y(n31460) );
  XNOR2_X1M_A12TR u1969 ( .A(sp[8]), .B(n2793), .Y(n31450) );
  XNOR2_X1M_A12TR u1970 ( .A(sp[7]), .B(n2792), .Y(n31440) );
  XNOR2_X1M_A12TR u1971 ( .A(sp[6]), .B(n2791), .Y(n31430) );
  XNOR2_X1M_A12TR u1972 ( .A(sp[5]), .B(n2790), .Y(n31420) );
  XNOR2_X1M_A12TR u1973 ( .A(sp[4]), .B(n2789), .Y(n31410) );
  XNOR2_X1M_A12TR u1974 ( .A(sp[3]), .B(n2788), .Y(n31400) );
  XNOR2_X1M_A12TR u1975 ( .A(sp[2]), .B(sp[1]), .Y(n31390) );
  XNOR2_X1M_A12TR u1976 ( .A(sp[13]), .B(n2798), .Y(n31500) );
  XNOR2_X1M_A12TR u1977 ( .A(sp[14]), .B(n2799), .Y(n31510) );
  MXIT2_X0P7M_A12TR u1978 ( .A(n2812), .B(n2813), .S0(n237), .Y(n966) );
  MXIT2_X0P7M_A12TR u1979 ( .A(n2804), .B(n2805), .S0(n237), .Y(n970) );
  MXIT2_X0P7M_A12TR u1980 ( .A(n2816), .B(n2817), .S0(n237), .Y(n964) );
  MXIT2_X0P7M_A12TR u1981 ( .A(n2806), .B(n2807), .S0(n237), .Y(n969) );
  MXIT2_X0P7M_A12TR u1982 ( .A(n2808), .B(n2809), .S0(n237), .Y(n968) );
  MXIT2_X0P7M_A12TR u1983 ( .A(n2810), .B(n2811), .S0(n237), .Y(n967) );
  MXIT2_X0P7M_A12TR u1984 ( .A(n2814), .B(n2815), .S0(n237), .Y(n965) );
  MXIT2_X0P7M_A12TR u1985 ( .A(n2818), .B(n2819), .S0(n237), .Y(n963) );
  XNOR2_X1M_A12TR u1986 ( .A(pc[1]), .B(pc[0]), .Y(n30100) );
  XNOR2_X1M_A12TR u1987 ( .A(pc[15]), .B(n2803), .Y(n30240) );
  NAND2_X1M_A12TR u1988 ( .A(pc[14]), .B(n2787), .Y(n2803) );
  XOR2_X1M_A12TR u1989 ( .A(pc[5]), .B(n2776), .Y(n30140) );
  XOR2_X1M_A12TR u1990 ( .A(pc[3]), .B(n2779), .Y(n30120) );
  XOR2_X1M_A12TR u1991 ( .A(pc[4]), .B(n2777), .Y(n30130) );
  XOR2_X1M_A12TR u1992 ( .A(pc[8]), .B(n2781), .Y(n30170) );
  XOR2_X1M_A12TR u1993 ( .A(pc[14]), .B(n2787), .Y(n30230) );
  XOR2_X1M_A12TR u1994 ( .A(pc[9]), .B(n2782), .Y(n30180) );
  XOR2_X1M_A12TR u1995 ( .A(pc[10]), .B(n2783), .Y(n30190) );
  XOR2_X1M_A12TR u1996 ( .A(pc[11]), .B(n2784), .Y(n30200) );
  XOR2_X1M_A12TR u1997 ( .A(pc[13]), .B(n2786), .Y(n30220) );
  XOR2_X1M_A12TR u1998 ( .A(pc[12]), .B(n2785), .Y(n30210) );
  XOR2_X1M_A12TR u1999 ( .A(pc[7]), .B(n2780), .Y(n30160) );
  XOR2_X1M_A12TR u2000 ( .A(pc[2]), .B(n2775), .Y(n30110) );
  XOR2_X1M_A12TR u2001 ( .A(pc[6]), .B(n2778), .Y(n30150) );
  MXIT4_X1M_A12TR u2002 ( .A(n1162), .B(regfil_6__4_), .C(n1154), .D(n1105), 
        .S0(n46), .S1(n236), .Y(n2813) );
  MXIT4_X1M_A12TR u2003 ( .A(n1158), .B(regfil_6__0_), .C(n1150), .D(
        regfil_7__0_), .S0(n46), .S1(n236), .Y(n2805) );
  MXIT4_X1M_A12TR u2004 ( .A(n1164), .B(regfil_6__6_), .C(n1156), .D(n1107), 
        .S0(n46), .S1(n236), .Y(n2817) );
  MXIT4_X1M_A12TR u2005 ( .A(n1159), .B(regfil_6__1_), .C(n1151), .D(n1102), 
        .S0(n46), .S1(n236), .Y(n2807) );
  MXIT4_X1M_A12TR u2006 ( .A(n1160), .B(regfil_6__2_), .C(n1152), .D(n1103), 
        .S0(n46), .S1(n236), .Y(n2809) );
  MXIT4_X1M_A12TR u2007 ( .A(n1161), .B(regfil_6__3_), .C(n1153), .D(n1104), 
        .S0(n46), .S1(n236), .Y(n2811) );
  MXIT4_X1M_A12TR u2008 ( .A(n1163), .B(regfil_6__5_), .C(n1155), .D(n1106), 
        .S0(n46), .S1(n236), .Y(n2815) );
  MXIT4_X1M_A12TR u2009 ( .A(n1165), .B(regfil_6__7_), .C(n1157), .D(n1108), 
        .S0(n46), .S1(n236), .Y(n2819) );
  MXIT4_X1M_A12TR u2010 ( .A(n1179), .B(regfil_2__4_), .C(n1171), .D(n1661), 
        .S0(n46), .S1(n236), .Y(n2812) );
  MXIT4_X1M_A12TR u2011 ( .A(n1175), .B(regfil_2__0_), .C(n1167), .D(n1657), 
        .S0(n46), .S1(n236), .Y(n2804) );
  MXIT4_X1M_A12TR u2012 ( .A(n1181), .B(regfil_2__6_), .C(n1173), .D(n1663), 
        .S0(n46), .S1(n236), .Y(n2816) );
  MXIT4_X1M_A12TR u2013 ( .A(n1176), .B(regfil_2__1_), .C(n1168), .D(n1658), 
        .S0(n46), .S1(n236), .Y(n2806) );
  MXIT4_X1M_A12TR u2014 ( .A(n1177), .B(regfil_2__2_), .C(n1169), .D(n1659), 
        .S0(n46), .S1(n236), .Y(n2808) );
  MXIT4_X1M_A12TR u2015 ( .A(n1178), .B(regfil_2__3_), .C(n1170), .D(n1660), 
        .S0(n46), .S1(n236), .Y(n2810) );
  MXIT4_X1M_A12TR u2016 ( .A(n1180), .B(regfil_2__5_), .C(n1172), .D(n1662), 
        .S0(n46), .S1(n236), .Y(n2814) );
  MXIT4_X1M_A12TR u2017 ( .A(n1182), .B(regfil_2__7_), .C(n1174), .D(n1664), 
        .S0(n46), .S1(n236), .Y(n2818) );
  AND2_X1M_A12TR u2018 ( .A(statesel[1]), .B(statesel[0]), .Y(n2772) );
  AND2_X1M_A12TR u2019 ( .A(statesel[3]), .B(n2774), .Y(n2773) );
  AND2_X1M_A12TR u2020 ( .A(statesel[2]), .B(n2772), .Y(n2774) );
  OR2_X1M_A12TR u2021 ( .A(pc[0]), .B(pc[1]), .Y(n2775) );
  AND2_X1M_A12TR u2022 ( .A(pc[4]), .B(n2777), .Y(n2776) );
  AND2_X1M_A12TR u2023 ( .A(pc[3]), .B(n2779), .Y(n2777) );
  AND2_X1M_A12TR u2024 ( .A(pc[5]), .B(n2776), .Y(n2778) );
  AND2_X1M_A12TR u2025 ( .A(pc[2]), .B(n2775), .Y(n2779) );
  AND2_X1M_A12TR u2026 ( .A(pc[6]), .B(n2778), .Y(n2780) );
  AND2_X1M_A12TR u2027 ( .A(pc[7]), .B(n2780), .Y(n2781) );
  AND2_X1M_A12TR u2028 ( .A(pc[8]), .B(n2781), .Y(n2782) );
  AND2_X1M_A12TR u2029 ( .A(pc[9]), .B(n2782), .Y(n2783) );
  AND2_X1M_A12TR u2030 ( .A(pc[10]), .B(n2783), .Y(n2784) );
  AND2_X1M_A12TR u2031 ( .A(pc[11]), .B(n2784), .Y(n2785) );
  AND2_X1M_A12TR u2032 ( .A(pc[12]), .B(n2785), .Y(n2786) );
  AND2_X1M_A12TR u2033 ( .A(pc[13]), .B(n2786), .Y(n2787) );
  OR2_X1M_A12TR u2034 ( .A(sp[1]), .B(sp[2]), .Y(n2788) );
  OR2_X1M_A12TR u2035 ( .A(n2788), .B(sp[3]), .Y(n2789) );
  OR2_X1M_A12TR u2036 ( .A(n2789), .B(sp[4]), .Y(n2790) );
  OR2_X1M_A12TR u2037 ( .A(n2790), .B(sp[5]), .Y(n2791) );
  OR2_X1M_A12TR u2038 ( .A(n2791), .B(sp[6]), .Y(n2792) );
  OR2_X1M_A12TR u2039 ( .A(n2792), .B(sp[7]), .Y(n2793) );
  OR2_X1M_A12TR u2040 ( .A(n2793), .B(sp[8]), .Y(n2794) );
  OR2_X1M_A12TR u2041 ( .A(n2794), .B(sp[9]), .Y(n2795) );
  OR2_X1M_A12TR u2042 ( .A(n2795), .B(sp[10]), .Y(n2796) );
  OR2_X1M_A12TR u2043 ( .A(n2796), .B(sp[11]), .Y(n2797) );
  OR2_X1M_A12TR u2044 ( .A(n2797), .B(sp[12]), .Y(n2798) );
  OR2_X1M_A12TR u2045 ( .A(n2798), .B(sp[13]), .Y(n2799) );
  AND2_X1M_A12TR u2046 ( .A(statesel[4]), .B(n2773), .Y(n2800) );
  TIELO_X1M_A12TR u2047 ( .Y(n4318) );
  NAND2_X0P5A_A12TR u2048 ( .A(n2820), .B(n2821), .Y(r201_b_as[1]) );
  AOI31_X0P5M_A12TR u2049 ( .A0(n2822), .A1(n2823), .A2(n2824), .B0(u3_u87_z_0), .Y(r201_b_as[0]) );
  NAND4_X0P5A_A12TR u2050 ( .A(n2825), .B(n2826), .C(n2827), .D(n2828), .Y(
        n2822) );
  OAI22_X0P5M_A12TR u2051 ( .A0(n2829), .A1(n2830), .B0(n2831), .B1(n2832), 
        .Y(n2827) );
  OAI222_X0P5M_A12TR u2052 ( .A0(n2824), .A1(n2833), .B0(n2820), .B1(n2834), 
        .C0(n2823), .C1(n2835), .Y(r201_a_9_) );
  OAI222_X0P5M_A12TR u2053 ( .A0(n2824), .A1(n2836), .B0(n2820), .B1(n2837), 
        .C0(n2823), .C1(n2838), .Y(r201_a_15_) );
  OAI222_X0P5M_A12TR u2054 ( .A0(n2824), .A1(n2839), .B0(n2820), .B1(n2840), 
        .C0(n2823), .C1(n2841), .Y(r201_a_14_) );
  OAI222_X0P5M_A12TR u2055 ( .A0(n2824), .A1(n2842), .B0(n2820), .B1(n2843), 
        .C0(n2823), .C1(n2844), .Y(r201_a_13_) );
  OAI222_X0P5M_A12TR u2056 ( .A0(n2824), .A1(n2845), .B0(n2820), .B1(n2846), 
        .C0(n2823), .C1(n2847), .Y(r201_a_12_) );
  OAI222_X0P5M_A12TR u2057 ( .A0(n2824), .A1(n2848), .B0(n2820), .B1(n2849), 
        .C0(n2823), .C1(n2850), .Y(r201_a_11_) );
  OAI222_X0P5M_A12TR u2058 ( .A0(n2824), .A1(n2851), .B0(n2820), .B1(n2852), 
        .C0(n2823), .C1(n2853), .Y(r201_a_10_) );
  OAI222_X0P5M_A12TR u2059 ( .A0(n2824), .A1(n2854), .B0(n2820), .B1(n2855), 
        .C0(n2823), .C1(n2856), .Y(r201_a_0_) );
  INV_X0P5B_A12TR u2060 ( .A(raddrhold[0]), .Y(n2856) );
  XOR2_X0P5M_A12TR u2061 ( .A(n2742), .B(n2857), .Y(r194_b_as[1]) );
  NAND2B_X0P5M_A12TR u2062 ( .AN(n2858), .B(n2859), .Y(n2857) );
  XOR2_X0P5M_A12TR u2063 ( .A(n2742), .B(n2860), .Y(r194_b_as[0]) );
  OAI211_X0P5M_A12TR u2064 ( .A0(n2861), .A1(state[5]), .B0(n2862), .C0(n2863), 
        .Y(n2860) );
  NAND2B_X0P5M_A12TR u2065 ( .AN(u3_u94_z_0), .B(n2823), .Y(r1606_b_as_6_) );
  INV_X0P5B_A12TR u2066 ( .A(n2864), .Y(r1606_b_as_2_) );
  AOI31_X0P5M_A12TR u2067 ( .A0(n2865), .A1(n2823), .A2(n2866), .B0(u3_u94_z_0), .Y(n2864) );
  AOI31_X0P5M_A12TR u2068 ( .A0(n2867), .A1(n2868), .A2(n2869), .B0(u3_u93_z_6), .Y(r1606_b_as_0_) );
  INV_X0P5B_A12TR u2069 ( .A(n2464), .Y(n4308) );
  INV_X0P5B_A12TR u2070 ( .A(n2463), .Y(n4309) );
  INV_X0P5B_A12TR u2071 ( .A(n2465), .Y(n4310) );
  INV_X0P5B_A12TR u2072 ( .A(n2462), .Y(n4311) );
  INV_X0P5B_A12TR u2073 ( .A(n2461), .Y(readmem) );
  INV_X0P5B_A12TR u2074 ( .A(n2460), .Y(n4313) );
  INV_X0P5B_A12TR u2075 ( .A(n2459), .Y(n4314) );
  INV_X0P5B_A12TR u2076 ( .A(n2458), .Y(n4315) );
  INV_X0P5B_A12TR u2077 ( .A(n2457), .Y(n4316) );
  INV_X0P5B_A12TR u2078 ( .A(n2456), .Y(inta) );
  OAI21_X0P5M_A12TR u2079 ( .A0(n2870), .A1(n2871), .B0(n2872), .Y(n2741) );
  MXIT2_X0P5M_A12TR u2080 ( .A(n2873), .B(n2874), .S0(n2875), .Y(n2872) );
  OAI211_X0P5M_A12TR u2081 ( .A0(n2876), .A1(n2877), .B0(n2878), .C0(n2879), 
        .Y(n2873) );
  AOI222_X0P5M_A12TR u2082 ( .A0(r1226_sum_8_), .A1(n2825), .B0(n1175), .B1(
        n2880), .C0(pc[8]), .C1(n2881), .Y(n2879) );
  AOI22_X0P5M_A12TR u2083 ( .A0(regfil_2__0_), .A1(n2882), .B0(n30170), .B1(
        n2883), .Y(n2878) );
  OAI21_X0P5M_A12TR u2084 ( .A0(n2830), .A1(n2884), .B0(n2885), .Y(n2740) );
  MXIT2_X0P5M_A12TR u2085 ( .A(n2886), .B(n2887), .S0(n2888), .Y(n2885) );
  OAI211_X0P5M_A12TR u2086 ( .A0(n2889), .A1(n2890), .B0(n2891), .C0(n2892), 
        .Y(n2887) );
  AOI222_X0P5M_A12TR u2087 ( .A0(state[4]), .A1(rdatahold[7]), .B0(n240), .B1(
        n2893), .C0(alures[7]), .C1(state[0]), .Y(n2892) );
  AOI21_X0P5M_A12TR u2088 ( .A0(n2894), .A1(n2895), .B0(n2896), .Y(n2891) );
  AOI31_X0P5M_A12TR u2089 ( .A0(n2897), .A1(n2898), .A2(n2899), .B0(n2900), 
        .Y(n2896) );
  AOI222_X0P5M_A12TR u2090 ( .A0(r1226_sum_7_), .A1(n2825), .B0(pc[7]), .B1(
        n2881), .C0(n1157), .C1(n2901), .Y(n2899) );
  AOI22_X0P5M_A12TR u2091 ( .A0(n1664), .A1(n2882), .B0(n30160), .B1(n2883), 
        .Y(n2898) );
  AOI22_X0P5M_A12TR u2092 ( .A0(sign), .A1(n2902), .B0(n1174), .B1(n2880), .Y(
        n2897) );
  INV_X0P5B_A12TR u2093 ( .A(n2483), .Y(n2886) );
  OAI221_X0P5M_A12TR u2094 ( .A0(n2483), .A1(n2903), .B0(n2830), .B1(n2904), 
        .C0(n2905), .Y(n2739) );
  NAND2_X0P5A_A12TR u2095 ( .A(datao[7]), .B(n2906), .Y(n2905) );
  OAI21_X0P5M_A12TR u2096 ( .A0(n2907), .A1(n2908), .B0(n2909), .Y(n2738) );
  MXIT2_X0P5M_A12TR u2097 ( .A(n2910), .B(n1108), .S0(n2911), .Y(n2909) );
  OAI221_X0P5M_A12TR u2098 ( .A0(n2912), .A1(n2913), .B0(n2914), .B1(n2915), 
        .C0(n2916), .Y(n2910) );
  AOI222_X0P5M_A12TR u2099 ( .A0(r1606_sum_7_), .A1(n2917), .B0(data_in[7]), .B1(
        n2918), .C0(n2919), .C1(n240), .Y(n2916) );
  AOI211_X0P5M_A12TR u2100 ( .A0(regfil_7__0_), .A1(n2920), .B0(n2921), .C0(
        n2922), .Y(n2907) );
  AO22_X0P5M_A12TR u2101 ( .A0(n2830), .A1(n2923), .B0(n2924), .B1(r201_sum_7_), .Y(n2921) );
  MXIT2_X0P5M_A12TR u2102 ( .A(n2925), .B(n2926), .S0(n2927), .Y(n2737) );
  AOI221_X0P5M_A12TR u2103 ( .A0(r201_sum_15_), .A1(n2928), .B0(rdatahold[7]), 
        .B1(n2929), .C0(n2930), .Y(n2926) );
  NAND4_X0P5A_A12TR u2104 ( .A(n2931), .B(n2932), .C(n2933), .D(n2934), .Y(
        n2736) );
  AOI22_X0P5M_A12TR u2105 ( .A0(n2935), .A1(n1182), .B0(r1226_sum_15_), .B1(
        n2936), .Y(n2934) );
  AOI22_X0P5M_A12TR u2106 ( .A0(n2937), .A1(regfil_2__7_), .B0(n2938), .B1(
        n1165), .Y(n2933) );
  AOI22_X0P5M_A12TR u2107 ( .A0(n2939), .A1(rdatahold[7]), .B0(sp[15]), .B1(
        n2940), .Y(n2932) );
  AOI22_X0P5M_A12TR u2108 ( .A0(n2941), .A1(r201_sum_15_), .B0(raddrhold[15]), 
        .B1(n2942), .Y(n2931) );
  OAI211_X0P5M_A12TR u2109 ( .A0(n2837), .A1(n2943), .B0(n2944), .C0(n2945), 
        .Y(n2735) );
  AOI221_X0P5M_A12TR u2110 ( .A0(n2946), .A1(r201_sum_15_), .B0(n2947), .B1(
        r1226_sum_15_), .C0(n2948), .Y(n2945) );
  AO22_X0P5M_A12TR u2111 ( .A0(n2949), .A1(n30240), .B0(n1165), .B1(n2950), 
        .Y(n2948) );
  AOI22_X0P5M_A12TR u2112 ( .A0(n2951), .A1(rdatahold[7]), .B0(r194_sum_15_), 
        .B1(n2952), .Y(n2944) );
  OAI221_X0P5M_A12TR u2113 ( .A0(n2953), .A1(n2954), .B0(n2955), .B1(n2956), 
        .C0(n2957), .Y(n2734) );
  MXIT2_X0P5M_A12TR u2114 ( .A(regfil_2__7_), .B(n2958), .S0(n2959), .Y(n2957)
         );
  OAI221_X0P5M_A12TR u2115 ( .A0(n2960), .A1(n2961), .B0(n2962), .B1(n2912), 
        .C0(n2963), .Y(n2958) );
  INV_X0P5B_A12TR u2116 ( .A(n2964), .Y(n2963) );
  INV_X0P5B_A12TR u2117 ( .A(r194_sum_15_), .Y(n2955) );
  INV_X0P5B_A12TR u2118 ( .A(r201_sum_15_), .Y(n2953) );
  MXIT2_X0P5M_A12TR u2119 ( .A(n2965), .B(n2832), .S0(n2966), .Y(n2733) );
  OA21A1OI2_X0P5M_A12TR u2120 ( .A0(n2924), .A1(n2967), .B0(n2968), .C0(n2969), 
        .Y(n2966) );
  NOR2_X0P5A_A12TR u2121 ( .A(reset), .B(n2970), .Y(n2969) );
  AOI221_X0P5M_A12TR u2122 ( .A0(alucout), .A1(n2971), .B0(r1606_sum_8_), .B1(
        n2972), .C0(n2973), .Y(n2965) );
  MXIT2_X0P5M_A12TR u2123 ( .A(n2974), .B(n2975), .S0(state[0]), .Y(n2973) );
  NAND2_X0P5A_A12TR u2124 ( .A(n2976), .B(n2823), .Y(n2974) );
  OAI211_X0P5M_A12TR u2125 ( .A0(n2977), .A1(n2978), .B0(n2979), .C0(n2980), 
        .Y(n2976) );
  AOI22_X0P5M_A12TR u2126 ( .A0(n1334), .A1(n2981), .B0(n2982), .B1(
        regfil_7__0_), .Y(n2980) );
  AOI31_X0P5M_A12TR u2127 ( .A0(n2825), .A1(n2832), .A2(n2983), .B0(n2984), 
        .Y(n2979) );
  NOR2_X0P5A_A12TR u2128 ( .A(n2985), .B(n2986), .Y(n2732) );
  AOI22_X0P5M_A12TR u2129 ( .A0(n2987), .A1(n2988), .B0(n2989), .B1(n2865), 
        .Y(n2985) );
  OAI31_X0P5M_A12TR u2130 ( .A0(n2990), .A1(n2991), .A2(n2992), .B0(n2993), 
        .Y(n2987) );
  MXIT2_X0P5M_A12TR u2131 ( .A(n2994), .B(n2995), .S0(statesel[1]), .Y(n2993)
         );
  NOR3_X0P5A_A12TR u2132 ( .A(n2996), .B(statesel[5]), .C(n2997), .Y(n2995) );
  OAI211_X0P5M_A12TR u2133 ( .A0(n2992), .A1(n2998), .B0(n2999), .C0(n3000), 
        .Y(n2994) );
  NAND3_X0P5A_A12TR u2134 ( .A(statesel[5]), .B(n3001), .C(n3002), .Y(n2999)
         );
  INV_X0P5B_A12TR u2135 ( .A(n3003), .Y(n2991) );
  MXIT2_X0P5M_A12TR u2136 ( .A(n3004), .B(n3005), .S0(n3006), .Y(n2731) );
  AND4_X0P5M_A12TR u2137 ( .A(n3007), .B(n3008), .C(n3009), .D(n30101), .Y(
        n3005) );
  AOI31_X0P5M_A12TR u2138 ( .A0(n2972), .A1(n30111), .A2(n30121), .B0(reset), 
        .Y(n30101) );
  OAI21_X0P5M_A12TR u2139 ( .A0(state[0]), .A1(n30131), .B0(n30141), .Y(n30121) );
  OA21A1OI2_X0P5M_A12TR u2140 ( .A0(n30151), .A1(n30161), .B0(n30171), .C0(
        n30181), .Y(n3009) );
  NOR3_X0P5A_A12TR u2141 ( .A(n30191), .B(u3_u93_z_6), .C(n30201), .Y(n30181)
         );
  INV_X0P5B_A12TR u2142 ( .A(n30211), .Y(n30151) );
  AOI22_X0P5M_A12TR u2143 ( .A0(n30221), .A1(n30231), .B0(n30241), .B1(n3025), 
        .Y(n3008) );
  NAND4_X0P5A_A12TR u2144 ( .A(n3026), .B(n3027), .C(n3028), .D(n3029), .Y(
        n3025) );
  OA21A1OI2_X0P5M_A12TR u2145 ( .A0(n3030), .A1(n3031), .B0(n3032), .C0(n3033), 
        .Y(n3029) );
  AOI21_X0P5M_A12TR u2146 ( .A0(n3034), .A1(n3035), .B0(n3036), .Y(n3033) );
  AOI211_X0P5M_A12TR u2147 ( .A0(n3037), .A1(n3038), .B0(n3039), .C0(n3040), 
        .Y(n3035) );
  AOI22_X0P5M_A12TR u2148 ( .A0(n3041), .A1(n3042), .B0(n236), .B1(n233), .Y(
        n3034) );
  OR3_X0P5M_A12TR u2149 ( .A(n3043), .B(n3044), .C(n3045), .Y(n3028) );
  OAI221_X0P5M_A12TR u2150 ( .A0(n3046), .A1(n3047), .B0(statesel[5]), .B1(
        n3048), .C0(n3049), .Y(n30231) );
  AOI32_X0P5M_A12TR u2151 ( .A0(n3050), .A1(n3051), .A2(statesel[3]), .B0(
        n3052), .B1(n3053), .Y(n3049) );
  INV_X0P5B_A12TR u2152 ( .A(n2996), .Y(n3053) );
  AO1B2_X0P5M_A12TR u2153 ( .B0(n3054), .B1(n3055), .A0N(n3056), .Y(n3050) );
  AOI211_X0P5M_A12TR u2154 ( .A0(n3054), .A1(n3057), .B0(n3058), .C0(n3059), 
        .Y(n3048) );
  OA21A1OI2_X0P5M_A12TR u2155 ( .A0(n3057), .A1(n3060), .B0(n3061), .C0(
        statesel[2]), .Y(n3059) );
  MXIT2_X0P5M_A12TR u2156 ( .A(n3062), .B(n3063), .S0(statesel[1]), .Y(n3058)
         );
  NAND2_X0P5A_A12TR u2157 ( .A(n3064), .B(n3047), .Y(n3063) );
  NAND2_X0P5A_A12TR u2158 ( .A(n3065), .B(statesel[4]), .Y(n3062) );
  AOI211_X0P5M_A12TR u2159 ( .A0(n3064), .A1(statesel[5]), .B0(n3066), .C0(
        n3067), .Y(n3046) );
  OA21A1OI2_X0P5M_A12TR u2160 ( .A0(statesel[3]), .A1(n2992), .B0(n3068), .C0(
        n3051), .Y(n3067) );
  INV_X0P5B_A12TR u2161 ( .A(n2998), .Y(n3064) );
  OAI221_X0P5M_A12TR u2162 ( .A0(n3069), .A1(n3070), .B0(n30201), .B1(n2972), 
        .C0(n3071), .Y(n30221) );
  INV_X0P5B_A12TR u2163 ( .A(n3072), .Y(n30201) );
  AOI22_X0P5M_A12TR u2164 ( .A0(n3073), .A1(n3074), .B0(n3075), .B1(n3076), 
        .Y(n3007) );
  OAI22_X0P5M_A12TR u2165 ( .A0(n2823), .A1(n3006), .B0(n3077), .B1(n2986), 
        .Y(n2730) );
  AOI221_X0P5M_A12TR u2166 ( .A0(n3078), .A1(n30141), .B0(n30241), .B1(n3079), 
        .C0(n3080), .Y(n3077) );
  OAI211_X0P5M_A12TR u2167 ( .A0(n3081), .A1(n3082), .B0(n3083), .C0(n3084), 
        .Y(n3080) );
  OAI211_X0P5M_A12TR u2168 ( .A0(n3085), .A1(n3076), .B0(state[0]), .C0(n2918), 
        .Y(n3083) );
  OA21A1OI2_X0P5M_A12TR u2169 ( .A0(n3081), .A1(n3086), .B0(n3087), .C0(
        state[5]), .Y(n3085) );
  AOI31_X0P5M_A12TR u2170 ( .A0(n3087), .A1(n30111), .A2(n3088), .B0(n3089), 
        .Y(n3082) );
  OA211_X0P5M_A12TR u2171 ( .A0(n2992), .A1(n3061), .B0(n3090), .C0(n3091), 
        .Y(n3081) );
  AOI211_X0P5M_A12TR u2172 ( .A0(n3092), .A1(n3051), .B0(n3093), .C0(n3094), 
        .Y(n3091) );
  MXIT2_X0P5M_A12TR u2173 ( .A(n3095), .B(n3096), .S0(n3055), .Y(n3094) );
  NOR2_X0P5A_A12TR u2174 ( .A(n3097), .B(statesel[0]), .Y(n3055) );
  OR2_X0P5M_A12TR u2175 ( .A(n3098), .B(n3051), .Y(n3096) );
  NAND2_X0P5A_A12TR u2176 ( .A(n3054), .B(statesel[3]), .Y(n3095) );
  MXIT2_X0P5M_A12TR u2177 ( .A(n3099), .B(n3100), .S0(statesel[2]), .Y(n3093)
         );
  AOI222_X0P5M_A12TR u2178 ( .A0(statesel[4]), .A1(statesel[1]), .B0(n3101), 
        .B1(n3057), .C0(n3102), .C1(n3047), .Y(n3099) );
  INV_X0P5B_A12TR u2179 ( .A(n3103), .Y(n3092) );
  OA21A1OI2_X0P5M_A12TR u2180 ( .A0(n3101), .A1(n3097), .B0(n3104), .C0(n3105), 
        .Y(n3090) );
  NOR2_X0P5A_A12TR u2181 ( .A(n2996), .B(n3068), .Y(n3105) );
  NAND2_X0P5A_A12TR u2182 ( .A(statesel[2]), .B(n3065), .Y(n2996) );
  OAI211_X0P5M_A12TR u2183 ( .A0(n3106), .A1(n3036), .B0(n3107), .C0(n3108), 
        .Y(n3079) );
  AND3_X0P5M_A12TR u2184 ( .A(n3109), .B(n3110), .C(n3111), .Y(n3108) );
  OA21A1OI2_X0P5M_A12TR u2185 ( .A0(n3045), .A1(n3043), .B0(n3112), .C0(n3113), 
        .Y(n3107) );
  INV_X0P5B_A12TR u2186 ( .A(n3114), .Y(n3106) );
  OAI22_X0P5M_A12TR u2187 ( .A0(n2972), .A1(n3006), .B0(n3115), .B1(n2986), 
        .Y(n2729) );
  AOI211_X0P5M_A12TR u2188 ( .A0(n3116), .A1(n30111), .B0(n3117), .C0(n3118), 
        .Y(n3115) );
  AOI31_X0P5M_A12TR u2189 ( .A0(n3119), .A1(n3027), .A2(n3120), .B0(n3121), 
        .Y(n3118) );
  AOI21_X0P5M_A12TR u2190 ( .A0(n3122), .A1(n3123), .B0(n3124), .Y(n3120) );
  OAI211_X0P5M_A12TR u2191 ( .A0(n3125), .A1(n3037), .B0(n3126), .C0(n3127), 
        .Y(n3119) );
  OAI21_X0P5M_A12TR u2192 ( .A0(n2984), .A1(n3128), .B0(n3129), .Y(n3126) );
  OAI211_X0P5M_A12TR u2193 ( .A0(n3130), .A1(n3131), .B0(n3132), .C0(n3133), 
        .Y(n3117) );
  NAND3_X0P5A_A12TR u2194 ( .A(n3074), .B(n3134), .C(n3135), .Y(n3132) );
  AOI22_X0P5M_A12TR u2195 ( .A0(n3136), .A1(n3072), .B0(n2918), .B1(n3076), 
        .Y(n3131) );
  INV_X0P5B_A12TR u2196 ( .A(n31371), .Y(n3130) );
  OAI21_X0P5M_A12TR u2197 ( .A0(state[2]), .A1(n3138), .B0(n31391), .Y(n3116)
         );
  OAI211_X0P5M_A12TR u2198 ( .A0(u3_u93_z_6), .A1(n31371), .B0(n3087), .C0(
        n3088), .Y(n31391) );
  AOI32_X0P5M_A12TR u2199 ( .A0(n31401), .A1(n31371), .A2(n3135), .B0(n3073), 
        .B1(n30141), .Y(n3138) );
  NAND3B_X0P5M_A12TR u2200 ( .AN(n31411), .B(n31421), .C(n31431), .Y(n31371)
         );
  AOI21_X0P5M_A12TR u2201 ( .A0(n31441), .A1(n3051), .B0(n31451), .Y(n31431)
         );
  AOI211_X0P5M_A12TR u2202 ( .A0(n31461), .A1(n2990), .B0(n3057), .C0(n3097), 
        .Y(n31451) );
  MXIT2_X0P5M_A12TR u2203 ( .A(n3054), .B(n31471), .S0(statesel[0]), .Y(n31461) );
  NOR2_X0P5A_A12TR u2204 ( .A(statesel[4]), .B(n3051), .Y(n31471) );
  OAI22_X0P5M_A12TR u2205 ( .A0(n2997), .A1(n2998), .B0(n31481), .B1(n3047), 
        .Y(n31441) );
  AOI22_X0P5M_A12TR u2206 ( .A0(n3098), .A1(n3052), .B0(n3102), .B1(n31491), 
        .Y(n31481) );
  NOR2_X0P5A_A12TR u2207 ( .A(n31491), .B(statesel[3]), .Y(n3098) );
  MXIT2_X0P5M_A12TR u2208 ( .A(n31501), .B(n31511), .S0(statesel[0]), .Y(
        n31421) );
  NOR2_X0P5A_A12TR u2209 ( .A(n2998), .B(n3068), .Y(n31511) );
  OAI21_X0P5M_A12TR u2210 ( .A0(n3051), .A1(n2992), .B0(n31521), .Y(n31501) );
  OAI22_X0P5M_A12TR u2211 ( .A0(n3153), .A1(n3006), .B0(n3154), .B1(n2986), 
        .Y(n2728) );
  AOI211_X0P5M_A12TR u2212 ( .A0(n3075), .A1(n3155), .B0(n3156), .C0(n3157), 
        .Y(n3154) );
  MXIT2_X0P5M_A12TR u2213 ( .A(n3158), .B(n3159), .S0(state[0]), .Y(n3157) );
  AOI22_X0P5M_A12TR u2214 ( .A0(n3155), .A1(n2972), .B0(n31401), .B1(n2971), 
        .Y(n3159) );
  NAND2_X0P5A_A12TR u2215 ( .A(n2894), .B(n2971), .Y(n3158) );
  AO21A1AI2_X0P5M_A12TR u2216 ( .A0(n3160), .A1(n3161), .B0(n3162), .C0(n3163), 
        .Y(n3156) );
  OAI21_X0P5M_A12TR u2217 ( .A0(n3164), .A1(n3124), .B0(n30241), .Y(n3163) );
  INV_X0P5B_A12TR u2218 ( .A(n3121), .Y(n30241) );
  INV_X0P5B_A12TR u2219 ( .A(n2988), .Y(n3162) );
  NAND2_X0P5A_A12TR u2220 ( .A(n3165), .B(n3071), .Y(n2988) );
  OA22_X0P5M_A12TR u2221 ( .A0(n3166), .A1(n3086), .B0(n3167), .B1(n3168), .Y(
        n3071) );
  MXIT2_X0P5M_A12TR u2222 ( .A(n3169), .B(n3170), .S0(statesel[0]), .Y(n3161)
         );
  AO21A1AI2_X0P5M_A12TR u2223 ( .A0(n3057), .A1(n31491), .B0(n3068), .C0(n3171), .Y(n3170) );
  NAND4_X0P5A_A12TR u2224 ( .A(statesel[5]), .B(n3001), .C(n3051), .D(n3057), 
        .Y(n3171) );
  NOR2B_X0P5M_A12TR u2225 ( .AN(n3104), .B(statesel[4]), .Y(n3169) );
  AOI21_X0P5M_A12TR u2226 ( .A0(statesel[1]), .A1(n3172), .B0(n31411), .Y(
        n3160) );
  AO1B2_X0P5M_A12TR u2227 ( .B0(n3173), .B1(statesel[1]), .A0N(n3174), .Y(
        n31411) );
  OAI31_X0P5M_A12TR u2228 ( .A0(n3175), .A1(n3176), .A2(n3104), .B0(n3097), 
        .Y(n3174) );
  NOR2_X0P5A_A12TR u2229 ( .A(n2998), .B(statesel[1]), .Y(n3104) );
  NAND2_X0P5A_A12TR u2230 ( .A(statesel[2]), .B(statesel[3]), .Y(n2998) );
  INV_X0P5B_A12TR u2231 ( .A(n3000), .Y(n3176) );
  OAI21_X0P5M_A12TR u2232 ( .A0(n2990), .A1(n3060), .B0(n3177), .Y(n3175) );
  NAND4_X0P5A_A12TR u2233 ( .A(statesel[3]), .B(statesel[4]), .C(n3047), .D(
        n3051), .Y(n3177) );
  NAND2_X0P5A_A12TR u2234 ( .A(statesel[1]), .B(n31491), .Y(n2990) );
  OAI21_X0P5M_A12TR u2235 ( .A0(n3056), .A1(statesel[3]), .B0(n3103), .Y(n3173) );
  AOI31_X0P5M_A12TR u2236 ( .A0(statesel[4]), .A1(n3097), .A2(n31491), .B0(
        n3066), .Y(n3056) );
  OAI221_X0P5M_A12TR u2237 ( .A0(n2992), .A1(n3061), .B0(statesel[0]), .B1(
        n31521), .C0(n3178), .Y(n3172) );
  AOI32_X0P5M_A12TR u2238 ( .A0(statesel[3]), .A1(statesel[5]), .A2(n3054), 
        .B0(n3002), .B1(n2997), .Y(n3178) );
  OAI22_X0P5M_A12TR u2239 ( .A0(n3179), .A1(n3006), .B0(n3180), .B1(n2986), 
        .Y(n2727) );
  NAND2_X0P5A_A12TR u2240 ( .A(n3181), .B(n3006), .Y(n2986) );
  AOI211_X0P5M_A12TR u2241 ( .A0(n3075), .A1(state[4]), .B0(n3182), .C0(n3183), 
        .Y(n3180) );
  AOI31_X0P5M_A12TR u2242 ( .A0(n3184), .A1(n3185), .A2(n3186), .B0(n3121), 
        .Y(n3183) );
  NAND3_X0P5A_A12TR u2243 ( .A(n2859), .B(n3004), .C(n30131), .Y(n3121) );
  AOI21_X0P5M_A12TR u2244 ( .A0(n3127), .A1(n3187), .B0(n3188), .Y(n3186) );
  OAI22_X0P5M_A12TR u2245 ( .A0(n3189), .A1(n3190), .B0(n3038), .B1(n3191), 
        .Y(n3187) );
  INV_X0P5B_A12TR u2246 ( .A(n3113), .Y(n3185) );
  AOI211_X0P5M_A12TR u2247 ( .A0(n3192), .A1(n3032), .B0(n233), .C0(n3193), 
        .Y(n3113) );
  OA211_X0P5M_A12TR u2248 ( .A0(sign), .A1(n3038), .B0(n3194), .C0(n3195), .Y(
        n3032) );
  AOI221_X0P5M_A12TR u2249 ( .A0(parity), .A1(n3196), .B0(zero), .B1(n2920), 
        .C0(n2922), .Y(n3195) );
  NOR2_X0P5A_A12TR u2250 ( .A(n3197), .B(n2832), .Y(n2922) );
  MXIT2_X0P5M_A12TR u2251 ( .A(n3198), .B(n3199), .S0(n236), .Y(n3194) );
  NOR2_X0P5A_A12TR u2252 ( .A(n3200), .B(n3201), .Y(n3199) );
  OAI222_X0P5M_A12TR u2253 ( .A0(parity), .A1(n3042), .B0(carry), .B1(n2831), 
        .C0(zero), .C1(n2829), .Y(n3198) );
  OAI211_X0P5M_A12TR u2254 ( .A0(n2920), .A1(n3128), .B0(n3043), .C0(n3112), 
        .Y(n3184) );
  AO21A1AI2_X0P5M_A12TR u2255 ( .A0(n46), .A1(n234), .B0(n236), .C0(n3202), 
        .Y(n3043) );
  MXIT2_X0P5M_A12TR u2256 ( .A(n3203), .B(n3204), .S0(n234), .Y(n3202) );
  NAND3_X0P5A_A12TR u2257 ( .A(n3205), .B(n3206), .C(n3207), .Y(n3182) );
  AO21A1AI2_X0P5M_A12TR u2258 ( .A0(n3155), .A1(state[0]), .B0(n3208), .C0(
        n2918), .Y(n3207) );
  OAI31_X0P5M_A12TR u2259 ( .A0(n3086), .A1(state[5]), .A2(n3209), .B0(n3210), 
        .Y(n3208) );
  INV_X0P5B_A12TR u2260 ( .A(n3211), .Y(n3209) );
  AO21A1AI2_X0P5M_A12TR u2261 ( .A0(n3212), .A1(n3087), .B0(n3089), .C0(n3211), 
        .Y(n3206) );
  OAI21_X0P5M_A12TR u2262 ( .A0(n3061), .A1(n3068), .B0(n3213), .Y(n3211) );
  MXIT2_X0P5M_A12TR u2263 ( .A(n3214), .B(n3215), .S0(statesel[1]), .Y(n3213)
         );
  OAI221_X0P5M_A12TR u2264 ( .A0(statesel[5]), .A1(n3216), .B0(n3100), .B1(
        n31491), .C0(n3000), .Y(n3215) );
  NAND2_X0P5A_A12TR u2265 ( .A(n3054), .B(n3065), .Y(n3000) );
  AOI22_X0P5M_A12TR u2266 ( .A0(n3097), .A1(n3101), .B0(n3003), .B1(n3052), 
        .Y(n3100) );
  NOR2_X0P5A_A12TR u2267 ( .A(n3097), .B(statesel[4]), .Y(n3052) );
  NOR2_X0P5A_A12TR u2268 ( .A(n3002), .B(n3065), .Y(n3003) );
  INV_X0P5B_A12TR u2269 ( .A(n3061), .Y(n3065) );
  AOI22_X0P5M_A12TR u2270 ( .A0(n3002), .A1(n3001), .B0(n3047), .B1(n31491), 
        .Y(n3216) );
  NOR2_X0P5A_A12TR u2271 ( .A(n3057), .B(n3047), .Y(n3002) );
  OAI211_X0P5M_A12TR u2272 ( .A0(statesel[0]), .A1(n3217), .B0(n3103), .C0(
        n3218), .Y(n3214) );
  AO21A1AI2_X0P5M_A12TR u2273 ( .A0(n3101), .A1(n3097), .B0(n3066), .C0(n3057), 
        .Y(n3218) );
  INV_X0P5B_A12TR u2274 ( .A(n31521), .Y(n3066) );
  NAND2_X0P5A_A12TR u2275 ( .A(statesel[2]), .B(n3102), .Y(n31521) );
  INV_X0P5B_A12TR u2276 ( .A(n2992), .Y(n3102) );
  INV_X0P5B_A12TR u2277 ( .A(n3060), .Y(n3101) );
  NAND2_X0P5A_A12TR u2278 ( .A(statesel[0]), .B(statesel[4]), .Y(n3060) );
  NAND3_X0P5A_A12TR u2279 ( .A(statesel[0]), .B(statesel[5]), .C(n3054), .Y(
        n3103) );
  INV_X0P5B_A12TR u2280 ( .A(n3001), .Y(n3054) );
  NAND2_X0P5A_A12TR u2281 ( .A(n2997), .B(n31491), .Y(n3001) );
  INV_X0P5B_A12TR u2282 ( .A(n3219), .Y(n3217) );
  AO21A1AI2_X0P5M_A12TR u2283 ( .A0(n2992), .A1(n3057), .B0(statesel[2]), .C0(
        n3068), .Y(n3219) );
  NAND2_X0P5A_A12TR u2284 ( .A(statesel[5]), .B(statesel[4]), .Y(n2992) );
  NAND2_X0P5A_A12TR u2285 ( .A(n2997), .B(n3097), .Y(n3068) );
  NAND2_X0P5A_A12TR u2286 ( .A(n3057), .B(n3047), .Y(n3061) );
  INV_X0P5B_A12TR u2287 ( .A(statesel[0]), .Y(n3047) );
  INV_X0P5B_A12TR u2288 ( .A(n3165), .Y(n3089) );
  AO21A1AI2_X0P5M_A12TR u2289 ( .A0(state[0]), .A1(n3087), .B0(n3220), .C0(
        n2971), .Y(n3205) );
  NAND4_X0P5A_A12TR u2290 ( .A(n3221), .B(n3222), .C(n3223), .D(n3224), .Y(
        n3006) );
  NOR3_X0P5A_A12TR u2291 ( .A(n3225), .B(state[5]), .C(n3226), .Y(n3224) );
  AO21A1AI2_X0P5M_A12TR u2292 ( .A0(n3227), .A1(n3228), .B0(n3229), .C0(n3230), 
        .Y(n3225) );
  OA21A1OI2_X0P5M_A12TR u2293 ( .A0(n3231), .A1(n3087), .B0(state[0]), .C0(
        n3232), .Y(n3223) );
  NOR2_X0P5A_A12TR u2294 ( .A(state[4]), .B(n3070), .Y(n3232) );
  OAI31_X0P5M_A12TR u2295 ( .A0(n3155), .A1(state[0]), .A2(n3220), .B0(n3233), 
        .Y(n3222) );
  INV_X0P5B_A12TR u2296 ( .A(n3210), .Y(n3220) );
  MXIT2_X0P5M_A12TR u2297 ( .A(n2912), .B(n3234), .S0(n3235), .Y(n2726) );
  MXIT2_X0P5M_A12TR u2298 ( .A(n3236), .B(n2912), .S0(n3235), .Y(n2725) );
  NOR2_X0P5A_A12TR u2299 ( .A(reset), .B(n3237), .Y(n2724) );
  MXIT2_X0P5M_A12TR u2300 ( .A(u3_u93_z_6), .B(writemem), .S0(n3238), .Y(n3237) );
  AOI32_X0P5M_A12TR u2301 ( .A0(n3073), .A1(state[2]), .A2(n3239), .B0(n3240), 
        .B1(n3241), .Y(n3238) );
  INV_X0P5B_A12TR u2302 ( .A(n3242), .Y(n3240) );
  MXT2_X0P5M_A12TR u2303 ( .A(n3243), .B(writeio), .S0(n3244), .Y(n2723) );
  AOI21_X0P5M_A12TR u2304 ( .A0(n3245), .A1(n3246), .B0(reset), .Y(n3244) );
  AOI21_X0P5M_A12TR u2305 ( .A0(waitr), .A1(state[0]), .B0(n30171), .Y(n3245)
         );
  NOR2_X0P5A_A12TR u2306 ( .A(state[0]), .B(reset), .Y(n3243) );
  MXIT2_X0P5M_A12TR u2307 ( .A(n2465), .B(n3247), .S0(n3248), .Y(n2722) );
  OAI221_X0P5M_A12TR u2308 ( .A0(n3168), .A1(n30171), .B0(n3166), .B1(n3179), 
        .C0(n3249), .Y(n3248) );
  AOI31_X0P5M_A12TR u2309 ( .A0(n3239), .A1(u3_u93_z_6), .A2(n3088), .B0(reset), .Y(n3249) );
  AO21A1AI2_X0P5M_A12TR u2310 ( .A0(n3135), .A1(n3155), .B0(n2894), .C0(n3181), 
        .Y(n3247) );
  OAI221_X0P5M_A12TR u2311 ( .A0(n2490), .A1(n2903), .B0(n2877), .B1(n2904), 
        .C0(n3250), .Y(n2721) );
  NAND2_X0P5A_A12TR u2312 ( .A(datao[0]), .B(n2906), .Y(n3250) );
  MXIT2_X0P5M_A12TR u2313 ( .A(n3251), .B(n3252), .S0(n3235), .Y(n2720) );
  MXIT2_X0P5M_A12TR u2314 ( .A(n2975), .B(n3251), .S0(n3235), .Y(n2719) );
  OAI221_X0P5M_A12TR u2315 ( .A0(n2489), .A1(n2903), .B0(n2904), .B1(n3253), 
        .C0(n3254), .Y(n2718) );
  NAND2_X0P5A_A12TR u2316 ( .A(datao[1]), .B(n2906), .Y(n3254) );
  MXIT2_X0P5M_A12TR u2317 ( .A(n3255), .B(n3256), .S0(n3235), .Y(n2717) );
  MXIT2_X0P5M_A12TR u2318 ( .A(n3257), .B(n3255), .S0(n3235), .Y(n2716) );
  OAI221_X0P5M_A12TR u2319 ( .A0(n2488), .A1(n2903), .B0(n2904), .B1(n3258), 
        .C0(n3259), .Y(n2715) );
  NAND2_X0P5A_A12TR u2320 ( .A(datao[2]), .B(n2906), .Y(n3259) );
  MXIT2_X0P5M_A12TR u2321 ( .A(n3260), .B(n3261), .S0(n3235), .Y(n2714) );
  MXIT2_X0P5M_A12TR u2322 ( .A(n3262), .B(n3260), .S0(n3235), .Y(n2713) );
  OAI221_X0P5M_A12TR u2323 ( .A0(n2487), .A1(n2903), .B0(n3263), .B1(n2904), 
        .C0(n3264), .Y(n2712) );
  NAND2_X0P5A_A12TR u2324 ( .A(datao[3]), .B(n2906), .Y(n3264) );
  MXIT2_X0P5M_A12TR u2325 ( .A(n3265), .B(n3266), .S0(n3235), .Y(n2711) );
  MXIT2_X0P5M_A12TR u2326 ( .A(n3267), .B(n3265), .S0(n3235), .Y(n2710) );
  OAI221_X0P5M_A12TR u2327 ( .A0(n2486), .A1(n2903), .B0(n2904), .B1(n3268), 
        .C0(n3269), .Y(n2709) );
  NAND2_X0P5A_A12TR u2328 ( .A(datao[4]), .B(n2906), .Y(n3269) );
  MXIT2_X0P5M_A12TR u2329 ( .A(n3270), .B(n3271), .S0(n3235), .Y(n2708) );
  MXIT2_X0P5M_A12TR u2330 ( .A(n3272), .B(n3270), .S0(n3235), .Y(n2707) );
  OAI221_X0P5M_A12TR u2331 ( .A0(n2485), .A1(n2903), .B0(n2904), .B1(n3273), 
        .C0(n3274), .Y(n2706) );
  NAND2_X0P5A_A12TR u2332 ( .A(datao[5]), .B(n2906), .Y(n3274) );
  MXIT2_X0P5M_A12TR u2333 ( .A(n3275), .B(n3276), .S0(n3235), .Y(n2705) );
  MXIT2_X0P5M_A12TR u2334 ( .A(n3277), .B(n3275), .S0(n3235), .Y(n2704) );
  OAI221_X0P5M_A12TR u2335 ( .A0(n2484), .A1(n2903), .B0(n2904), .B1(n3278), 
        .C0(n3279), .Y(n2703) );
  NAND2_X0P5A_A12TR u2336 ( .A(datao[6]), .B(n2906), .Y(n3279) );
  INV_X0P5B_A12TR u2337 ( .A(n3280), .Y(n2906) );
  NAND2_X0P5A_A12TR u2338 ( .A(n2823), .B(n3280), .Y(n2904) );
  NAND2_X0P5A_A12TR u2339 ( .A(u3_u93_z_6), .B(n3280), .Y(n2903) );
  OAI31_X0P5M_A12TR u2340 ( .A0(n3166), .A1(reset), .A2(n30171), .B0(n3281), 
        .Y(n3280) );
  NAND3_X0P5A_A12TR u2341 ( .A(n3282), .B(n2894), .C(n30161), .Y(n3281) );
  MXIT2_X0P5M_A12TR u2342 ( .A(n3283), .B(n3284), .S0(n3235), .Y(n2702) );
  MXIT2_X0P5M_A12TR u2343 ( .A(n3285), .B(n3283), .S0(n3235), .Y(n2701) );
  MXIT2_X0P5M_A12TR u2344 ( .A(n3286), .B(n3252), .S0(n3287), .Y(n2700) );
  INV_X0P5B_A12TR u2345 ( .A(data_in[0]), .Y(n3252) );
  MXIT2_X0P5M_A12TR u2346 ( .A(n3288), .B(n3256), .S0(n3287), .Y(n2699) );
  INV_X0P5B_A12TR u2347 ( .A(data_in[1]), .Y(n3256) );
  MXIT2_X0P5M_A12TR u2348 ( .A(n3128), .B(n3261), .S0(n3287), .Y(n2698) );
  INV_X0P5B_A12TR u2349 ( .A(data_in[2]), .Y(n3261) );
  MXIT2_X0P5M_A12TR u2350 ( .A(n2828), .B(n3266), .S0(n3287), .Y(n2697) );
  INV_X0P5B_A12TR u2351 ( .A(data_in[3]), .Y(n3266) );
  MXIT2_X0P5M_A12TR u2352 ( .A(n3289), .B(n3271), .S0(n3287), .Y(n2696) );
  INV_X0P5B_A12TR u2353 ( .A(data_in[4]), .Y(n3271) );
  MXIT2_X0P5M_A12TR u2354 ( .A(n3290), .B(n3276), .S0(n3287), .Y(n2695) );
  INV_X0P5B_A12TR u2355 ( .A(data_in[5]), .Y(n3276) );
  MXIT2_X0P5M_A12TR u2356 ( .A(n3291), .B(n3284), .S0(n3287), .Y(n2694) );
  INV_X0P5B_A12TR u2357 ( .A(data_in[6]), .Y(n3284) );
  MXIT2_X0P5M_A12TR u2358 ( .A(n3292), .B(n3234), .S0(n3287), .Y(n2693) );
  AND4_X0P5M_A12TR u2359 ( .A(n30111), .B(n3233), .C(n2972), .D(n3293), .Y(
        n3287) );
  NOR3_X0P5A_A12TR u2360 ( .A(n3294), .B(reset), .C(n3295), .Y(n3293) );
  INV_X0P5B_A12TR u2361 ( .A(data_in[7]), .Y(n3234) );
  MXT2_X0P5M_A12TR u2362 ( .A(alucin), .B(carry), .S0(n3296), .Y(n2692) );
  AOI21_X0P5M_A12TR u2363 ( .A0(n3111), .A1(n3297), .B0(n3298), .Y(n3296) );
  AO22_X0P5M_A12TR u2364 ( .A0(alusel[0]), .A1(n3299), .B0(n3300), .B1(n236), 
        .Y(n2691) );
  AO1B2_X0P5M_A12TR u2365 ( .B0(n46), .B1(n3300), .A0N(n3301), .Y(n2690) );
  MXIT2_X0P5M_A12TR u2366 ( .A(alusel[1]), .B(n3302), .S0(n3303), .Y(n3301) );
  NOR2_X0P5A_A12TR u2367 ( .A(n3286), .B(n3036), .Y(n3302) );
  AO22_X0P5M_A12TR u2368 ( .A0(alusel[2]), .A1(n3299), .B0(n3300), .B1(n237), 
        .Y(n2689) );
  NOR2_X0P5A_A12TR u2369 ( .A(n3299), .B(n3227), .Y(n3300) );
  INV_X0P5B_A12TR u2370 ( .A(n3303), .Y(n3299) );
  MXIT2_X0P5M_A12TR u2371 ( .A(n3304), .B(n2828), .S0(n3305), .Y(n2688) );
  MXIT2_X0P5M_A12TR u2372 ( .A(n3306), .B(n3307), .S0(n3305), .Y(n2687) );
  NOR2_X0P5A_A12TR u2373 ( .A(n3308), .B(n46), .Y(n3307) );
  MXIT2_X0P5M_A12TR u2374 ( .A(n3309), .B(n3310), .S0(n3305), .Y(n2686) );
  OAI22_X0P5M_A12TR u2375 ( .A0(n3298), .A1(n3109), .B0(n3311), .B1(n3312), 
        .Y(n3305) );
  NOR2_X0P5A_A12TR u2376 ( .A(n3308), .B(n237), .Y(n3310) );
  MXIT2_X0P5M_A12TR u2377 ( .A(n3313), .B(n3289), .S0(n3314), .Y(n2685) );
  MXIT2_X0P5M_A12TR u2378 ( .A(n3315), .B(n3290), .S0(n3314), .Y(n2684) );
  NOR3_X0P5A_A12TR u2379 ( .A(n3316), .B(n3193), .C(n3298), .Y(n3314) );
  MXIT2_X0P5M_A12TR u2380 ( .A(n3317), .B(n3318), .S0(n3319), .Y(n2683) );
  AOI211_X0P5M_A12TR u2381 ( .A0(n3320), .A1(n3321), .B0(reset), .C0(n3322), 
        .Y(n3319) );
  MXIT2_X0P5M_A12TR u2382 ( .A(n3323), .B(n3324), .S0(n3325), .Y(n2682) );
  NOR3_X0P5A_A12TR u2383 ( .A(n3326), .B(reset), .C(n3327), .Y(n3325) );
  OAI22_X0P5M_A12TR u2384 ( .A0(n3318), .A1(n3328), .B0(n3329), .B1(n3330), 
        .Y(n3326) );
  INV_X0P5B_A12TR u2385 ( .A(eienb), .Y(n3318) );
  INV_X0P5B_A12TR u2386 ( .A(ei), .Y(n3324) );
  AOI21_X0P5M_A12TR u2387 ( .A0(eienb), .A1(n2972), .B0(reset), .Y(n3323) );
  OA21A1OI2_X0P5M_A12TR u2388 ( .A0(n3322), .A1(n3331), .B0(n3332), .C0(reset), 
        .Y(n2681) );
  MXIT2_X0P5M_A12TR u2389 ( .A(n3333), .B(n2461), .S0(n3334), .Y(n2680) );
  AOI211_X0P5M_A12TR u2390 ( .A0(n3322), .A1(n3134), .B0(n3335), .C0(n3336), 
        .Y(n3334) );
  NOR3_X0P5A_A12TR u2391 ( .A(n3210), .B(intcyc), .C(n3337), .Y(n3336) );
  OAI21_X0P5M_A12TR u2392 ( .A0(n3097), .A1(n3338), .B0(n3339), .Y(n2679) );
  AOI22_X0P5M_A12TR u2393 ( .A0(n3340), .A1(n3341), .B0(n35750), .B1(n3342), 
        .Y(n3339) );
  OAI21_X0P5M_A12TR u2394 ( .A0(n3036), .A1(n3343), .B0(n3227), .Y(n3341) );
  INV_X0P5B_A12TR u2395 ( .A(statesel[5]), .Y(n3097) );
  AO21A1AI2_X0P5M_A12TR u2396 ( .A0(n3344), .A1(n3345), .B0(n3346), .C0(n3347), 
        .Y(n2678) );
  MXIT2_X0P5M_A12TR u2397 ( .A(n3342), .B(n3348), .S0(statesel[0]), .Y(n3347)
         );
  NOR3_X0P5A_A12TR u2398 ( .A(n3349), .B(n3350), .C(n3351), .Y(n3345) );
  OAI31_X0P5M_A12TR u2399 ( .A0(n3352), .A1(n236), .A2(n3353), .B0(n3297), .Y(
        n3349) );
  AOI211_X0P5M_A12TR u2400 ( .A0(n3354), .A1(n237), .B0(n3355), .C0(n3124), 
        .Y(n3344) );
  OAI211_X0P5M_A12TR u2401 ( .A0(n3193), .A1(n3356), .B0(n3110), .C0(n3357), 
        .Y(n3124) );
  OAI21_X0P5M_A12TR u2402 ( .A0(n3051), .A1(n3338), .B0(n3358), .Y(n2677) );
  AOI22_X0P5M_A12TR u2403 ( .A0(n3340), .A1(n3359), .B0(n35710), .B1(n3342), 
        .Y(n3358) );
  NAND4B_X0P5M_A12TR u2404 ( .AN(n3360), .B(n3111), .C(n3361), .D(n3362), .Y(
        n3359) );
  AOI221_X0P5M_A12TR u2405 ( .A0(n3363), .A1(n3353), .B0(n3354), .B1(n3290), 
        .C0(n3355), .Y(n3362) );
  OAI31_X0P5M_A12TR u2406 ( .A0(n3192), .A1(n2984), .A2(n3036), .B0(n3364), 
        .Y(n3355) );
  NAND2_X0P5A_A12TR u2407 ( .A(n3365), .B(n3366), .Y(n3364) );
  INV_X0P5B_A12TR u2408 ( .A(n3352), .Y(n3363) );
  OAI31_X0P5M_A12TR u2409 ( .A0(n3289), .A1(n3286), .A2(n3367), .B0(n3109), 
        .Y(n3360) );
  INV_X0P5B_A12TR u2410 ( .A(statesel[1]), .Y(n3051) );
  OAI21_X0P5M_A12TR u2411 ( .A0(n31491), .A1(n3338), .B0(n3368), .Y(n2676) );
  AOI22_X0P5M_A12TR u2412 ( .A0(n3340), .A1(n3369), .B0(n35720), .B1(n3342), 
        .Y(n3368) );
  NAND4_X0P5A_A12TR u2413 ( .A(n3297), .B(n3361), .C(n3357), .D(n3370), .Y(
        n3369) );
  OA21A1OI2_X0P5M_A12TR u2414 ( .A0(n3371), .A1(n3372), .B0(n3127), .C0(n3373), 
        .Y(n3370) );
  AOI21_X0P5M_A12TR u2415 ( .A0(n3374), .A1(n3375), .B0(n3193), .Y(n3373) );
  INV_X0P5B_A12TR u2416 ( .A(n3376), .Y(n3361) );
  INV_X0P5B_A12TR u2417 ( .A(statesel[2]), .Y(n31491) );
  OAI21_X0P5M_A12TR u2418 ( .A0(n3057), .A1(n3338), .B0(n3377), .Y(n2675) );
  AOI22_X0P5M_A12TR u2419 ( .A0(n3340), .A1(n3378), .B0(n35730), .B1(n3342), 
        .Y(n3377) );
  NAND4_X0P5A_A12TR u2420 ( .A(n3379), .B(n3380), .C(n3381), .D(n3382), .Y(
        n3378) );
  AOI211_X0P5M_A12TR u2421 ( .A0(n3383), .A1(n3127), .B0(n3351), .C0(n3376), 
        .Y(n3382) );
  AOI21_X0P5M_A12TR u2422 ( .A0(n3384), .A1(n2867), .B0(n3193), .Y(n3376) );
  INV_X0P5B_A12TR u2423 ( .A(statesel[3]), .Y(n3057) );
  OAI21_X0P5M_A12TR u2424 ( .A0(n2997), .A1(n3338), .B0(n3385), .Y(n2674) );
  AOI22_X0P5M_A12TR u2425 ( .A0(n3340), .A1(n3386), .B0(n35740), .B1(n3342), 
        .Y(n3385) );
  AOI31_X0P5M_A12TR u2426 ( .A0(n30141), .A1(n30111), .A2(n3179), .B0(n3348), 
        .Y(n3342) );
  NAND3_X0P5A_A12TR u2427 ( .A(n3381), .B(n3380), .C(n3387), .Y(n3386) );
  AOI22_X0P5M_A12TR u2428 ( .A0(n3366), .A1(n3388), .B0(n3127), .B1(n3389), 
        .Y(n3387) );
  AOI211_X0P5M_A12TR u2429 ( .A0(n3390), .A1(n3127), .B0(n3391), .C0(n3030), 
        .Y(n3381) );
  INV_X0P5B_A12TR u2430 ( .A(n3392), .Y(n3030) );
  INV_X0P5B_A12TR u2431 ( .A(n3393), .Y(n3391) );
  NAND2_X0P5A_A12TR u2432 ( .A(n3394), .B(n3395), .Y(n3390) );
  INV_X0P5B_A12TR u2433 ( .A(n3346), .Y(n3340) );
  NAND3_X0P5A_A12TR u2434 ( .A(n3338), .B(n30111), .C(n30131), .Y(n3346) );
  INV_X0P5B_A12TR u2435 ( .A(n3348), .Y(n3338) );
  NOR3_X0P5A_A12TR u2436 ( .A(n3235), .B(n3396), .C(n3397), .Y(n3348) );
  OAI22_X0P5M_A12TR u2437 ( .A0(n3398), .A1(reset), .B0(n3298), .B1(n3399), 
        .Y(n3397) );
  AOI211_X0P5M_A12TR u2438 ( .A0(n2894), .A1(n3212), .B0(n3400), .C0(n3401), 
        .Y(n3398) );
  OAI211_X0P5M_A12TR u2439 ( .A0(n3086), .A1(n3166), .B0(n3165), .C0(n3402), 
        .Y(n3401) );
  AOI21_X0P5M_A12TR u2440 ( .A0(n3072), .A1(n3136), .B0(n3403), .Y(n3165) );
  OAI21_X0P5M_A12TR u2441 ( .A0(n2972), .A1(n3004), .B0(n2914), .Y(n3136) );
  OAI22_X0P5M_A12TR u2442 ( .A0(n3329), .A1(n3404), .B0(n3405), .B1(n3190), 
        .Y(n3400) );
  NOR3_X0P5A_A12TR u2443 ( .A(n3168), .B(reset), .C(n3242), .Y(n3235) );
  INV_X0P5B_A12TR u2444 ( .A(statesel[4]), .Y(n2997) );
  OAI21_X0P5M_A12TR u2445 ( .A0(n2877), .A1(n2884), .B0(n3406), .Y(n2673) );
  MXIT2_X0P5M_A12TR u2446 ( .A(n3407), .B(n3408), .S0(n2888), .Y(n3406) );
  OAI211_X0P5M_A12TR u2447 ( .A0(n3409), .A1(n2890), .B0(n3410), .C0(n3411), 
        .Y(n3408) );
  AOI222_X0P5M_A12TR u2448 ( .A0(rdatahold[0]), .A1(state[4]), .B0(n247), .B1(
        n2893), .C0(alures[0]), .C1(state[0]), .Y(n3411) );
  AOI21_X0P5M_A12TR u2449 ( .A0(n2894), .A1(n2874), .B0(n3412), .Y(n3410) );
  AOI31_X0P5M_A12TR u2450 ( .A0(n3413), .A1(n3414), .A2(n3415), .B0(n2900), 
        .Y(n3412) );
  AOI222_X0P5M_A12TR u2451 ( .A0(n2880), .A1(n1167), .B0(n2882), .B1(n1657), 
        .C0(n2902), .C1(carry), .Y(n3415) );
  MXIT2_X0P5M_A12TR u2452 ( .A(n2883), .B(n2881), .S0(pc[0]), .Y(n3414) );
  AOI22_X0P5M_A12TR u2453 ( .A0(n1150), .A1(n2901), .B0(n2825), .B1(n3416), 
        .Y(n3413) );
  INV_X0P5B_A12TR u2454 ( .A(n2498), .Y(n2874) );
  INV_X0P5B_A12TR u2455 ( .A(n2490), .Y(n3407) );
  OAI21_X0P5M_A12TR u2456 ( .A0(n2884), .A1(n3253), .B0(n3417), .Y(n26721) );
  MXIT2_X0P5M_A12TR u2457 ( .A(n3418), .B(n3419), .S0(n2888), .Y(n3417) );
  OAI211_X0P5M_A12TR u2458 ( .A0(n2890), .A1(n3420), .B0(n3421), .C0(n3422), 
        .Y(n3419) );
  AOI222_X0P5M_A12TR u2459 ( .A0(rdatahold[1]), .A1(state[4]), .B0(n246), .B1(
        n2893), .C0(alures[1]), .C1(state[0]), .Y(n3422) );
  AOI22_X0P5M_A12TR u2460 ( .A0(n3423), .A1(n3424), .B0(n2894), .B1(n3425), 
        .Y(n3421) );
  OAI211_X0P5M_A12TR u2461 ( .A0(n3426), .A1(n3427), .B0(n3428), .C0(n3429), 
        .Y(n3424) );
  AOI211_X0P5M_A12TR u2462 ( .A0(n1658), .A1(n2882), .B0(n3430), .C0(n2902), 
        .Y(n3429) );
  AO22_X0P5M_A12TR u2463 ( .A0(n2880), .A1(n1168), .B0(n2883), .B1(n30100), 
        .Y(n3430) );
  AOI22_X0P5M_A12TR u2464 ( .A0(pc[1]), .A1(n2881), .B0(n1151), .B1(n2901), 
        .Y(n3428) );
  INV_X0P5B_A12TR u2465 ( .A(r1226_sum_1_), .Y(n3427) );
  INV_X0P5B_A12TR u2466 ( .A(n2489), .Y(n3418) );
  OAI21_X0P5M_A12TR u2467 ( .A0(n2884), .A1(n3258), .B0(n3431), .Y(n26711) );
  MXIT2_X0P5M_A12TR u2468 ( .A(n3432), .B(n3433), .S0(n2888), .Y(n3431) );
  OAI211_X0P5M_A12TR u2469 ( .A0(n2890), .A1(n3434), .B0(n3435), .C0(n3436), 
        .Y(n3433) );
  AOI222_X0P5M_A12TR u2470 ( .A0(rdatahold[2]), .A1(state[4]), .B0(n245), .B1(
        n2893), .C0(alures[2]), .C1(state[0]), .Y(n3436) );
  AOI21_X0P5M_A12TR u2471 ( .A0(n2894), .A1(n3437), .B0(n3438), .Y(n3435) );
  AOI31_X0P5M_A12TR u2472 ( .A0(n3439), .A1(n3440), .A2(n3441), .B0(n2900), 
        .Y(n3438) );
  AOI222_X0P5M_A12TR u2473 ( .A0(r1226_sum_2_), .A1(n2825), .B0(pc[2]), .B1(
        n2881), .C0(n1152), .C1(n2901), .Y(n3441) );
  AOI22_X0P5M_A12TR u2474 ( .A0(n1659), .A1(n2882), .B0(n30110), .B1(n2883), 
        .Y(n3440) );
  AOI22_X0P5M_A12TR u2475 ( .A0(parity), .A1(n2902), .B0(n1169), .B1(n2880), 
        .Y(n3439) );
  INV_X0P5B_A12TR u2476 ( .A(n2488), .Y(n3432) );
  OAI221_X0P5M_A12TR u2477 ( .A0(n3442), .A1(n3443), .B0(n3263), .B1(n2884), 
        .C0(n3444), .Y(n26701) );
  MXIT2_X0P5M_A12TR u2478 ( .A(n3445), .B(n3446), .S0(n2888), .Y(n3444) );
  OAI221_X0P5M_A12TR u2479 ( .A0(n3004), .A1(n3447), .B0(n3179), .B1(n3265), 
        .C0(n3448), .Y(n3446) );
  AOI222_X0P5M_A12TR u2480 ( .A0(n244), .A1(n2893), .B0(n3423), .B1(n3449), 
        .C0(n2894), .C1(n3450), .Y(n3448) );
  OAI221_X0P5M_A12TR u2481 ( .A0(n3451), .A1(n3452), .B0(n3426), .B1(n3453), 
        .C0(n3454), .Y(n3449) );
  AOI222_X0P5M_A12TR u2482 ( .A0(n1170), .A1(n2880), .B0(n1660), .B1(n2882), 
        .C0(n30120), .C1(n2883), .Y(n3454) );
  INV_X0P5B_A12TR u2483 ( .A(r1226_sum_3_), .Y(n3453) );
  INV_X0P5B_A12TR u2484 ( .A(n2487), .Y(n3445) );
  OAI21_X0P5M_A12TR u2485 ( .A0(n2884), .A1(n3268), .B0(n3455), .Y(n26691) );
  MXIT2_X0P5M_A12TR u2486 ( .A(n3456), .B(n3457), .S0(n2888), .Y(n3455) );
  OAI211_X0P5M_A12TR u2487 ( .A0(n2890), .A1(n3458), .B0(n3459), .C0(n3460), 
        .Y(n3457) );
  AOI222_X0P5M_A12TR u2488 ( .A0(rdatahold[4]), .A1(state[4]), .B0(n243), .B1(
        n2893), .C0(alures[4]), .C1(state[0]), .Y(n3460) );
  AOI21_X0P5M_A12TR u2489 ( .A0(n2894), .A1(n3461), .B0(n3462), .Y(n3459) );
  AOI31_X0P5M_A12TR u2490 ( .A0(n3463), .A1(n3464), .A2(n3465), .B0(n2900), 
        .Y(n3462) );
  AOI222_X0P5M_A12TR u2491 ( .A0(r1226_sum_4_), .A1(n2825), .B0(pc[4]), .B1(
        n2881), .C0(n1154), .C1(n2901), .Y(n3465) );
  AOI22_X0P5M_A12TR u2492 ( .A0(n1661), .A1(n2882), .B0(n30130), .B1(n2883), 
        .Y(n3464) );
  AOI22_X0P5M_A12TR u2493 ( .A0(auxcar), .A1(n2902), .B0(n1171), .B1(n2880), 
        .Y(n3463) );
  INV_X0P5B_A12TR u2494 ( .A(n2486), .Y(n3456) );
  OAI221_X0P5M_A12TR u2495 ( .A0(n3442), .A1(n3466), .B0(n2884), .B1(n3273), 
        .C0(n3467), .Y(n26681) );
  MXIT2_X0P5M_A12TR u2496 ( .A(n3468), .B(n3469), .S0(n2888), .Y(n3467) );
  OAI221_X0P5M_A12TR u2497 ( .A0(n3004), .A1(n3470), .B0(n3179), .B1(n3275), 
        .C0(n3471), .Y(n3469) );
  AOI222_X0P5M_A12TR u2498 ( .A0(n242), .A1(n2893), .B0(n3423), .B1(n3472), 
        .C0(n2894), .C1(n3473), .Y(n3471) );
  OAI221_X0P5M_A12TR u2499 ( .A0(n3451), .A1(n3474), .B0(n3426), .B1(n3475), 
        .C0(n3476), .Y(n3472) );
  AOI222_X0P5M_A12TR u2500 ( .A0(n1172), .A1(n2880), .B0(n1662), .B1(n2882), 
        .C0(n30140), .C1(n2883), .Y(n3476) );
  INV_X0P5B_A12TR u2501 ( .A(r1226_sum_5_), .Y(n3475) );
  INV_X0P5B_A12TR u2502 ( .A(n2881), .Y(n3451) );
  INV_X0P5B_A12TR u2503 ( .A(n2485), .Y(n3468) );
  AO21A1AI2_X0P5M_A12TR u2504 ( .A0(n3423), .A1(n2901), .B0(n3477), .C0(n2888), 
        .Y(n3442) );
  INV_X0P5B_A12TR u2505 ( .A(n2900), .Y(n3423) );
  OAI21_X0P5M_A12TR u2506 ( .A0(n2884), .A1(n3278), .B0(n3478), .Y(n26671) );
  MXIT2_X0P5M_A12TR u2507 ( .A(n3479), .B(n3480), .S0(n2888), .Y(n3478) );
  OAI211_X0P5M_A12TR u2508 ( .A0(n2890), .A1(n3481), .B0(n3482), .C0(n3483), 
        .Y(n3480) );
  AOI222_X0P5M_A12TR u2509 ( .A0(rdatahold[6]), .A1(state[4]), .B0(n241), .B1(
        n2893), .C0(alures[6]), .C1(state[0]), .Y(n3483) );
  INV_X0P5B_A12TR u2510 ( .A(n3484), .Y(n2893) );
  AOI21_X0P5M_A12TR u2511 ( .A0(n2894), .A1(n3485), .B0(n3486), .Y(n3482) );
  AOI31_X0P5M_A12TR u2512 ( .A0(n3487), .A1(n3488), .A2(n3489), .B0(n2900), 
        .Y(n3486) );
  AOI222_X0P5M_A12TR u2513 ( .A0(r1226_sum_6_), .A1(n2825), .B0(pc[6]), .B1(
        n2881), .C0(n1156), .C1(n2901), .Y(n3489) );
  AOI22_X0P5M_A12TR u2514 ( .A0(n1663), .A1(n2882), .B0(n30150), .B1(n2883), 
        .Y(n3488) );
  AOI22_X0P5M_A12TR u2515 ( .A0(zero), .A1(n2902), .B0(n1173), .B1(n2880), .Y(
        n3487) );
  INV_X0P5B_A12TR u2516 ( .A(n2876), .Y(n2902) );
  INV_X0P5B_A12TR u2517 ( .A(n2484), .Y(n3479) );
  NAND3B_X0P5M_A12TR u2518 ( .AN(n3490), .B(n2826), .C(n2888), .Y(n2884) );
  OAI211_X0P5M_A12TR u2519 ( .A0(n3312), .A1(n3490), .B0(n2875), .C0(n3491), 
        .Y(n2888) );
  AOI2XB1_X0P5M_A12TR u2520 ( .A1N(n3492), .A0(n3493), .B0(n3396), .Y(n3491)
         );
  MXIT2_X0P5M_A12TR u2521 ( .A(n3494), .B(n3069), .S0(state[0]), .Y(n3493) );
  NAND2_X0P5A_A12TR u2522 ( .A(state[3]), .B(n30111), .Y(n3494) );
  NAND4_X0P5A_A12TR u2523 ( .A(n3495), .B(n3496), .C(n3497), .D(n3498), .Y(
        n26661) );
  AOI22_X0P5M_A12TR u2524 ( .A0(n2935), .A1(n1167), .B0(n2936), .B1(n3416), 
        .Y(n3498) );
  AOI22_X0P5M_A12TR u2525 ( .A0(n2937), .A1(n1657), .B0(n2938), .B1(n1150), 
        .Y(n3497) );
  AOI22_X0P5M_A12TR u2526 ( .A0(rdatahold2[0]), .A1(n2939), .B0(n31370), .B1(
        n2940), .Y(n3496) );
  AOI22_X0P5M_A12TR u2527 ( .A0(r201_sum_0_), .A1(n2941), .B0(raddrhold[0]), 
        .B1(n2942), .Y(n3495) );
  NAND4_X0P5A_A12TR u2528 ( .A(n3499), .B(n3500), .C(n3501), .D(n3502), .Y(
        n26651) );
  AOI22_X0P5M_A12TR u2529 ( .A0(n1168), .A1(n2935), .B0(r1226_sum_1_), .B1(
        n2936), .Y(n3502) );
  AOI22_X0P5M_A12TR u2530 ( .A0(n1658), .A1(n2937), .B0(n1151), .B1(n2938), 
        .Y(n3501) );
  AOI22_X0P5M_A12TR u2531 ( .A0(rdatahold2[1]), .A1(n2939), .B0(sp[1]), .B1(
        n2940), .Y(n3500) );
  AOI22_X0P5M_A12TR u2532 ( .A0(r201_sum_1_), .A1(n2941), .B0(raddrhold[1]), 
        .B1(n2942), .Y(n3499) );
  NAND4_X0P5A_A12TR u2533 ( .A(n3503), .B(n3504), .C(n3505), .D(n3506), .Y(
        n26641) );
  AOI22_X0P5M_A12TR u2534 ( .A0(n1169), .A1(n2935), .B0(r1226_sum_2_), .B1(
        n2936), .Y(n3506) );
  AOI22_X0P5M_A12TR u2535 ( .A0(n1659), .A1(n2937), .B0(n1152), .B1(n2938), 
        .Y(n3505) );
  AOI22_X0P5M_A12TR u2536 ( .A0(rdatahold2[2]), .A1(n2939), .B0(sp[2]), .B1(
        n2940), .Y(n3504) );
  AOI22_X0P5M_A12TR u2537 ( .A0(r201_sum_2_), .A1(n2941), .B0(raddrhold[2]), 
        .B1(n2942), .Y(n3503) );
  NAND4_X0P5A_A12TR u2538 ( .A(n3507), .B(n3508), .C(n3509), .D(n3510), .Y(
        n26631) );
  AOI22_X0P5M_A12TR u2539 ( .A0(n1170), .A1(n2935), .B0(r1226_sum_3_), .B1(
        n2936), .Y(n3510) );
  AOI22_X0P5M_A12TR u2540 ( .A0(n1660), .A1(n2937), .B0(n1153), .B1(n2938), 
        .Y(n3509) );
  AOI22_X0P5M_A12TR u2541 ( .A0(rdatahold2[3]), .A1(n2939), .B0(sp[3]), .B1(
        n2940), .Y(n3508) );
  AOI22_X0P5M_A12TR u2542 ( .A0(r201_sum_3_), .A1(n2941), .B0(raddrhold[3]), 
        .B1(n2942), .Y(n3507) );
  NAND4_X0P5A_A12TR u2543 ( .A(n3511), .B(n3512), .C(n3513), .D(n3514), .Y(
        n26621) );
  AOI22_X0P5M_A12TR u2544 ( .A0(n1171), .A1(n2935), .B0(r1226_sum_4_), .B1(
        n2936), .Y(n3514) );
  AOI22_X0P5M_A12TR u2545 ( .A0(n1661), .A1(n2937), .B0(n1154), .B1(n2938), 
        .Y(n3513) );
  AOI22_X0P5M_A12TR u2546 ( .A0(rdatahold2[4]), .A1(n2939), .B0(sp[4]), .B1(
        n2940), .Y(n3512) );
  AOI22_X0P5M_A12TR u2547 ( .A0(r201_sum_4_), .A1(n2941), .B0(raddrhold[4]), 
        .B1(n2942), .Y(n3511) );
  NAND4_X0P5A_A12TR u2548 ( .A(n3515), .B(n3516), .C(n3517), .D(n3518), .Y(
        n26611) );
  AOI22_X0P5M_A12TR u2549 ( .A0(n1172), .A1(n2935), .B0(r1226_sum_5_), .B1(
        n2936), .Y(n3518) );
  AOI22_X0P5M_A12TR u2550 ( .A0(n1662), .A1(n2937), .B0(n1155), .B1(n2938), 
        .Y(n3517) );
  AOI22_X0P5M_A12TR u2551 ( .A0(rdatahold2[5]), .A1(n2939), .B0(sp[5]), .B1(
        n2940), .Y(n3516) );
  AOI22_X0P5M_A12TR u2552 ( .A0(r201_sum_5_), .A1(n2941), .B0(raddrhold[5]), 
        .B1(n2942), .Y(n3515) );
  NAND4_X0P5A_A12TR u2553 ( .A(n3519), .B(n3520), .C(n3521), .D(n3522), .Y(
        n26601) );
  AOI22_X0P5M_A12TR u2554 ( .A0(n1173), .A1(n2935), .B0(r1226_sum_6_), .B1(
        n2936), .Y(n3522) );
  AOI22_X0P5M_A12TR u2555 ( .A0(n1663), .A1(n2937), .B0(n1156), .B1(n2938), 
        .Y(n3521) );
  AOI22_X0P5M_A12TR u2556 ( .A0(rdatahold2[6]), .A1(n2939), .B0(sp[6]), .B1(
        n2940), .Y(n3520) );
  AOI22_X0P5M_A12TR u2557 ( .A0(r201_sum_6_), .A1(n2941), .B0(raddrhold[6]), 
        .B1(n2942), .Y(n3519) );
  NAND4_X0P5A_A12TR u2558 ( .A(n3523), .B(n3524), .C(n3525), .D(n3526), .Y(
        n26591) );
  AOI22_X0P5M_A12TR u2559 ( .A0(n2935), .A1(n1174), .B0(n2936), .B1(
        r1226_sum_7_), .Y(n3526) );
  AOI22_X0P5M_A12TR u2560 ( .A0(n2937), .A1(n1664), .B0(n2938), .B1(n1157), 
        .Y(n3525) );
  AOI22_X0P5M_A12TR u2561 ( .A0(rdatahold2[7]), .A1(n2939), .B0(sp[7]), .B1(
        n2940), .Y(n3524) );
  AOI22_X0P5M_A12TR u2562 ( .A0(n2941), .A1(r201_sum_7_), .B0(raddrhold[7]), 
        .B1(n2942), .Y(n3523) );
  NAND4_X0P5A_A12TR u2563 ( .A(n3527), .B(n3528), .C(n3529), .D(n3530), .Y(
        n26581) );
  AOI22_X0P5M_A12TR u2564 ( .A0(n2935), .A1(n1175), .B0(n2936), .B1(
        r1226_sum_8_), .Y(n3530) );
  AOI22_X0P5M_A12TR u2565 ( .A0(n2937), .A1(regfil_2__0_), .B0(n2938), .B1(
        n1158), .Y(n3529) );
  AOI22_X0P5M_A12TR u2566 ( .A0(rdatahold[0]), .A1(n2939), .B0(sp[8]), .B1(
        n2940), .Y(n3528) );
  AOI22_X0P5M_A12TR u2567 ( .A0(r201_sum_8_), .A1(n2941), .B0(raddrhold[8]), 
        .B1(n2942), .Y(n3527) );
  NAND4_X0P5A_A12TR u2568 ( .A(n3531), .B(n3532), .C(n3533), .D(n3534), .Y(
        n2657) );
  AOI22_X0P5M_A12TR u2569 ( .A0(n2935), .A1(n1176), .B0(r1226_sum_9_), .B1(
        n2936), .Y(n3534) );
  AOI22_X0P5M_A12TR u2570 ( .A0(n2937), .A1(regfil_2__1_), .B0(n2938), .B1(
        n1159), .Y(n3533) );
  AOI22_X0P5M_A12TR u2571 ( .A0(rdatahold[1]), .A1(n2939), .B0(sp[9]), .B1(
        n2940), .Y(n3532) );
  AOI22_X0P5M_A12TR u2572 ( .A0(r201_sum_9_), .A1(n2941), .B0(raddrhold[9]), 
        .B1(n2942), .Y(n3531) );
  NAND4_X0P5A_A12TR u2573 ( .A(n3535), .B(n3536), .C(n3537), .D(n3538), .Y(
        n2656) );
  AOI22_X0P5M_A12TR u2574 ( .A0(n2935), .A1(n1177), .B0(r1226_sum_10_), .B1(
        n2936), .Y(n3538) );
  AOI22_X0P5M_A12TR u2575 ( .A0(n2937), .A1(regfil_2__2_), .B0(n2938), .B1(
        n1160), .Y(n3537) );
  AOI22_X0P5M_A12TR u2576 ( .A0(rdatahold[2]), .A1(n2939), .B0(sp[10]), .B1(
        n2940), .Y(n3536) );
  AOI22_X0P5M_A12TR u2577 ( .A0(r201_sum_10_), .A1(n2941), .B0(raddrhold[10]), 
        .B1(n2942), .Y(n3535) );
  NAND4_X0P5A_A12TR u2578 ( .A(n3539), .B(n3540), .C(n3541), .D(n3542), .Y(
        n2655) );
  AOI22_X0P5M_A12TR u2579 ( .A0(n2935), .A1(n1178), .B0(r1226_sum_11_), .B1(
        n2936), .Y(n3542) );
  AOI22_X0P5M_A12TR u2580 ( .A0(n2937), .A1(regfil_2__3_), .B0(n2938), .B1(
        n1161), .Y(n3541) );
  AOI22_X0P5M_A12TR u2581 ( .A0(rdatahold[3]), .A1(n2939), .B0(sp[11]), .B1(
        n2940), .Y(n3540) );
  AOI22_X0P5M_A12TR u2582 ( .A0(r201_sum_11_), .A1(n2941), .B0(raddrhold[11]), 
        .B1(n2942), .Y(n3539) );
  NAND4_X0P5A_A12TR u2583 ( .A(n3543), .B(n3544), .C(n3545), .D(n3546), .Y(
        n2654) );
  AOI22_X0P5M_A12TR u2584 ( .A0(n2935), .A1(n1179), .B0(r1226_sum_12_), .B1(
        n2936), .Y(n3546) );
  AOI22_X0P5M_A12TR u2585 ( .A0(n2937), .A1(regfil_2__4_), .B0(n2938), .B1(
        n1162), .Y(n3545) );
  AOI22_X0P5M_A12TR u2586 ( .A0(rdatahold[4]), .A1(n2939), .B0(sp[12]), .B1(
        n2940), .Y(n3544) );
  AOI22_X0P5M_A12TR u2587 ( .A0(r201_sum_12_), .A1(n2941), .B0(raddrhold[12]), 
        .B1(n2942), .Y(n3543) );
  NAND4_X0P5A_A12TR u2588 ( .A(n3547), .B(n3548), .C(n3549), .D(n3550), .Y(
        n2653) );
  AOI22_X0P5M_A12TR u2589 ( .A0(n2935), .A1(n1180), .B0(r1226_sum_13_), .B1(
        n2936), .Y(n3550) );
  AOI22_X0P5M_A12TR u2590 ( .A0(n2937), .A1(regfil_2__5_), .B0(n2938), .B1(
        n1163), .Y(n3549) );
  AOI22_X0P5M_A12TR u2591 ( .A0(rdatahold[5]), .A1(n2939), .B0(sp[13]), .B1(
        n2940), .Y(n3548) );
  AOI22_X0P5M_A12TR u2592 ( .A0(r201_sum_13_), .A1(n2941), .B0(raddrhold[13]), 
        .B1(n2942), .Y(n3547) );
  NAND4_X0P5A_A12TR u2593 ( .A(n3551), .B(n3552), .C(n3553), .D(n3554), .Y(
        n2652) );
  AOI22_X0P5M_A12TR u2594 ( .A0(n2935), .A1(n1181), .B0(r1226_sum_14_), .B1(
        n2936), .Y(n3554) );
  INV_X0P5B_A12TR u2595 ( .A(n3555), .Y(n2936) );
  AO21A1AI2_X0P5M_A12TR u2596 ( .A0(n3366), .A1(n3556), .B0(n3557), .C0(n3558), 
        .Y(n3555) );
  OAI21_X0P5M_A12TR u2597 ( .A0(n3286), .A1(n3367), .B0(n3559), .Y(n3557) );
  OAI21_X0P5M_A12TR u2598 ( .A0(n3560), .A1(n3045), .B0(n3127), .Y(n3559) );
  INV_X0P5B_A12TR u2599 ( .A(n3192), .Y(n3045) );
  AND3_X0P5M_A12TR u2600 ( .A(n3354), .B(n3203), .C(n3558), .Y(n2935) );
  AOI22_X0P5M_A12TR u2601 ( .A0(n2937), .A1(regfil_2__6_), .B0(n2938), .B1(
        n1164), .Y(n3553) );
  AOI21B_X0P5M_A12TR u2602 ( .A0(n3228), .A1(n3380), .B0N(n3558), .Y(n2938) );
  AND3_X0P5M_A12TR u2603 ( .A(n3354), .B(n3204), .C(n3558), .Y(n2937) );
  NOR2_X0P5A_A12TR u2604 ( .A(n3352), .B(n2828), .Y(n3354) );
  NAND2_X0P5A_A12TR u2605 ( .A(n3308), .B(n234), .Y(n3352) );
  INV_X0P5B_A12TR u2606 ( .A(n3367), .Y(n3308) );
  NAND2_X0P5A_A12TR u2607 ( .A(n3127), .B(n3128), .Y(n3367) );
  AOI22_X0P5M_A12TR u2608 ( .A0(rdatahold[6]), .A1(n2939), .B0(sp[14]), .B1(
        n2940), .Y(n3552) );
  AND3_X0P5M_A12TR u2609 ( .A(n3366), .B(n3561), .C(n3558), .Y(n2940) );
  NOR2_X0P5A_A12TR u2610 ( .A(n2942), .B(n2972), .Y(n3558) );
  NOR2_X0P5A_A12TR u2611 ( .A(n2942), .B(n30111), .Y(n2939) );
  AOI22_X0P5M_A12TR u2612 ( .A0(r201_sum_14_), .A1(n2941), .B0(raddrhold[14]), 
        .B1(n2942), .Y(n3551) );
  NOR2_X0P5A_A12TR u2613 ( .A(n2942), .B(n2823), .Y(n2941) );
  NAND2_X0P5A_A12TR u2614 ( .A(n3181), .B(n3562), .Y(n2942) );
  OAI211_X0P5M_A12TR u2615 ( .A0(n3399), .A1(n3229), .B0(n3402), .C0(n3563), 
        .Y(n3562) );
  NOR3_X0P5A_A12TR u2616 ( .A(n3564), .B(n3565), .C(n3403), .Y(n3563) );
  AND3_X0P5M_A12TR u2617 ( .A(n3076), .B(n3004), .C(n2918), .Y(n3403) );
  NOR3_X0P5A_A12TR u2618 ( .A(n3405), .B(n3189), .C(n3190), .Y(n3564) );
  OA21A1OI2_X0P5M_A12TR u2619 ( .A0(n3556), .A1(n3561), .B0(n3320), .C0(n3566), 
        .Y(n3402) );
  AND4_X0P5M_A12TR u2620 ( .A(n2989), .B(n2984), .C(n235), .D(n3286), .Y(n3566) );
  NAND4_X0P5A_A12TR u2621 ( .A(n3567), .B(n3393), .C(n3316), .D(n2869), .Y(
        n3561) );
  NAND4B_X0P5M_A12TR u2622 ( .AN(n3388), .B(n3384), .C(n2867), .D(n3123), .Y(
        n3556) );
  NAND3_X0P5A_A12TR u2623 ( .A(n3191), .B(n3568), .C(n3375), .Y(n3388) );
  INV_X0P5B_A12TR u2624 ( .A(n3188), .Y(n3399) );
  OAI211_X0P5M_A12TR u2625 ( .A0(n3123), .A1(n3111), .B0(n3569), .C0(n3109), 
        .Y(n3188) );
  NAND3_X0P5A_A12TR u2626 ( .A(n3570), .B(n3027), .C(n35711), .Y(n3109) );
  AO21A1AI2_X0P5M_A12TR u2627 ( .A0(n35721), .A1(n2984), .B0(n3365), .C0(n3127), .Y(n3569) );
  OAI221_X0P5M_A12TR u2628 ( .A0(n3251), .A1(n35731), .B0(n35741), .B1(n35751), 
        .C0(n3576), .Y(n2651) );
  MXIT2_X0P5M_A12TR u2629 ( .A(aluoprb_0_), .B(n3577), .S0(n3578), .Y(n3576)
         );
  NOR2_X0P5A_A12TR u2630 ( .A(state[5]), .B(n3036), .Y(n3577) );
  OAI222_X0P5M_A12TR u2631 ( .A0(n3579), .A1(n35751), .B0(n3255), .B1(n35731), 
        .C0(n2457), .C1(n3578), .Y(n2650) );
  OAI222_X0P5M_A12TR u2632 ( .A0(n3580), .A1(n35751), .B0(n3260), .B1(n35731), 
        .C0(n2458), .C1(n3578), .Y(n2649) );
  OAI222_X0P5M_A12TR u2633 ( .A0(n3581), .A1(n35751), .B0(n3265), .B1(n35731), 
        .C0(n2459), .C1(n3578), .Y(n2648) );
  OAI222_X0P5M_A12TR u2634 ( .A0(n3582), .A1(n35751), .B0(n3270), .B1(n35731), 
        .C0(n2463), .C1(n3578), .Y(n2647) );
  OAI222_X0P5M_A12TR u2635 ( .A0(n3583), .A1(n35751), .B0(n3275), .B1(n35731), 
        .C0(n2460), .C1(n3578), .Y(n2646) );
  OAI222_X0P5M_A12TR u2636 ( .A0(n3584), .A1(n35751), .B0(n3283), .B1(n35731), 
        .C0(n2464), .C1(n3578), .Y(n2645) );
  OAI222_X0P5M_A12TR u2637 ( .A0(n3585), .A1(n35751), .B0(n2912), .B1(n35731), 
        .C0(n2462), .C1(n3578), .Y(n2644) );
  OAI21_X0P5M_A12TR u2638 ( .A0(n3226), .A1(n2972), .B0(n3578), .Y(n35731) );
  NAND3_X0P5A_A12TR u2639 ( .A(n3578), .B(n30111), .C(n3122), .Y(n35751) );
  OAI21_X0P5M_A12TR u2640 ( .A0(n3380), .A1(n3298), .B0(n3586), .Y(n3578) );
  AOI32_X0P5M_A12TR u2641 ( .A0(n3282), .A1(n3226), .A2(n3076), .B0(n3587), 
        .B1(n3181), .Y(n3586) );
  INV_X0P5B_A12TR u2642 ( .A(n3133), .Y(n3587) );
  NAND3_X0P5A_A12TR u2643 ( .A(n3076), .B(n2972), .C(n3135), .Y(n3133) );
  MXIT2_X0P5M_A12TR u2644 ( .A(n3588), .B(n3589), .S0(n3590), .Y(n2643) );
  MXIT2_X0P5M_A12TR u2645 ( .A(rdatahold2[2]), .B(alupar), .S0(u3_u93_z_6), 
        .Y(n3589) );
  INV_X0P5B_A12TR u2646 ( .A(parity), .Y(n3588) );
  MXIT2_X0P5M_A12TR u2647 ( .A(n3591), .B(n3592), .S0(n3590), .Y(n2642) );
  MXIT2_X0P5M_A12TR u2648 ( .A(rdatahold2[6]), .B(aluzout), .S0(u3_u93_z_6), 
        .Y(n3592) );
  INV_X0P5B_A12TR u2649 ( .A(zero), .Y(n3591) );
  MXIT2_X0P5M_A12TR u2650 ( .A(n3201), .B(n3593), .S0(n3590), .Y(n2641) );
  AOI222_X0P5M_A12TR u2651 ( .A0(alusout), .A1(n3004), .B0(n3073), .B1(
        alures[7]), .C0(rdatahold2[7]), .C1(n2823), .Y(n3593) );
  INV_X0P5B_A12TR u2652 ( .A(sign), .Y(n3201) );
  MXIT2_X0P5M_A12TR u2653 ( .A(n3594), .B(n3595), .S0(n3596), .Y(n2640) );
  AOI211_X0P5M_A12TR u2654 ( .A0(n2928), .A1(r1606_sum_7_), .B0(n3597), .C0(
        n2930), .Y(n3595) );
  OAI22_X0P5M_A12TR u2655 ( .A0(n2823), .A1(n2915), .B0(n3585), .B1(n3598), 
        .Y(n2930) );
  MXIT2_X0P5M_A12TR u2656 ( .A(n3599), .B(n3600), .S0(n3601), .Y(n2639) );
  AOI31_X0P5M_A12TR u2657 ( .A0(n2865), .A1(n2866), .A2(n2968), .B0(n3590), 
        .Y(n3601) );
  OAI31_X0P5M_A12TR u2658 ( .A0(n3294), .A1(n3295), .A2(n3317), .B0(n3602), 
        .Y(n3590) );
  NAND2_X0P5A_A12TR u2659 ( .A(n3603), .B(n3181), .Y(n3602) );
  NOR3_X0P5A_A12TR u2660 ( .A(n3604), .B(reset), .C(n3605), .Y(n2968) );
  AOI21_X0P5M_A12TR u2661 ( .A0(rdatahold2[4]), .A1(state[4]), .B0(n3606), .Y(
        n3599) );
  MXT2_X0P5M_A12TR u2662 ( .A(n3607), .B(aluaxc), .S0(u3_u93_z_6), .Y(n3606)
         );
  NOR2B_X0P5M_A12TR u2663 ( .AN(r1606_sum_8_), .B(state[0]), .Y(n3607) );
  OAI21_X0P5M_A12TR u2664 ( .A0(n3608), .A1(n2908), .B0(n3609), .Y(n2638) );
  MXIT2_X0P5M_A12TR u2665 ( .A(n3610), .B(regfil_7__0_), .S0(n2911), .Y(n3609)
         );
  OAI221_X0P5M_A12TR u2666 ( .A0(n2913), .A1(n3251), .B0(n2914), .B1(n3611), 
        .C0(n3612), .Y(n3610) );
  AOI222_X0P5M_A12TR u2667 ( .A0(r1606_sum_0_), .A1(n2917), .B0(data_in[0]), .B1(
        n2918), .C0(n247), .C1(n2919), .Y(n3612) );
  AOI222_X0P5M_A12TR u2668 ( .A0(n2923), .A1(n2877), .B0(r201_sum_0_), .B1(
        n2924), .C0(n1102), .C1(n2982), .Y(n3608) );
  OAI21_X0P5M_A12TR u2669 ( .A0(n3613), .A1(n2908), .B0(n3614), .Y(n2637) );
  MXIT2_X0P5M_A12TR u2670 ( .A(n3615), .B(n1102), .S0(n2911), .Y(n3614) );
  OAI221_X0P5M_A12TR u2671 ( .A0(n2913), .A1(n3255), .B0(n2914), .B1(n3616), 
        .C0(n3617), .Y(n3615) );
  AOI222_X0P5M_A12TR u2672 ( .A0(r1606_sum_1_), .A1(n2917), .B0(data_in[1]), .B1(
        n2918), .C0(n246), .C1(n2919), .Y(n3617) );
  AOI222_X0P5M_A12TR u2673 ( .A0(n2923), .A1(n3253), .B0(r201_sum_1_), .B1(
        n2924), .C0(n1103), .C1(n2982), .Y(n3613) );
  OAI21_X0P5M_A12TR u2674 ( .A0(n3618), .A1(n2908), .B0(n3619), .Y(n2636) );
  MXIT2_X0P5M_A12TR u2675 ( .A(n3620), .B(n1103), .S0(n2911), .Y(n3619) );
  OAI221_X0P5M_A12TR u2676 ( .A0(n2913), .A1(n3260), .B0(n2914), .B1(n3621), 
        .C0(n3622), .Y(n3620) );
  AOI222_X0P5M_A12TR u2677 ( .A0(r1606_sum_2_), .A1(n2917), .B0(data_in[2]), .B1(
        n2918), .C0(n245), .C1(n2919), .Y(n3622) );
  AOI222_X0P5M_A12TR u2678 ( .A0(n2923), .A1(n3258), .B0(r201_sum_2_), .B1(
        n2924), .C0(n2982), .C1(n1104), .Y(n3618) );
  OAI21_X0P5M_A12TR u2679 ( .A0(n3623), .A1(n2908), .B0(n3624), .Y(n2635) );
  MXIT2_X0P5M_A12TR u2680 ( .A(n3625), .B(n1104), .S0(n2911), .Y(n3624) );
  OAI221_X0P5M_A12TR u2681 ( .A0(n2913), .A1(n3265), .B0(n2914), .B1(n3447), 
        .C0(n3626), .Y(n3625) );
  AOI222_X0P5M_A12TR u2682 ( .A0(r1606_sum_3_), .A1(n2917), .B0(data_in[3]), .B1(
        n2918), .C0(n244), .C1(n2919), .Y(n3626) );
  AOI222_X0P5M_A12TR u2683 ( .A0(n2923), .A1(n3263), .B0(r201_sum_3_), .B1(
        n2924), .C0(n1105), .C1(n2982), .Y(n3623) );
  OAI21_X0P5M_A12TR u2684 ( .A0(n3627), .A1(n2908), .B0(n3628), .Y(n2634) );
  MXIT2_X0P5M_A12TR u2685 ( .A(n3629), .B(n1105), .S0(n2911), .Y(n3628) );
  OAI221_X0P5M_A12TR u2686 ( .A0(n2913), .A1(n3270), .B0(n2914), .B1(n3630), 
        .C0(n3631), .Y(n3629) );
  AOI222_X0P5M_A12TR u2687 ( .A0(r1606_sum_4_), .A1(n2917), .B0(data_in[4]), .B1(
        n2918), .C0(n243), .C1(n2919), .Y(n3631) );
  AOI222_X0P5M_A12TR u2688 ( .A0(n2923), .A1(n3268), .B0(r201_sum_4_), .B1(
        n2924), .C0(n1106), .C1(n2982), .Y(n3627) );
  OAI21_X0P5M_A12TR u2689 ( .A0(n3632), .A1(n2908), .B0(n3633), .Y(n2633) );
  MXIT2_X0P5M_A12TR u2690 ( .A(n3634), .B(n1106), .S0(n2911), .Y(n3633) );
  OAI221_X0P5M_A12TR u2691 ( .A0(n2913), .A1(n3275), .B0(n2914), .B1(n3470), 
        .C0(n3635), .Y(n3634) );
  AOI222_X0P5M_A12TR u2692 ( .A0(r1606_sum_5_), .A1(n2917), .B0(data_in[5]), .B1(
        n2918), .C0(n242), .C1(n2919), .Y(n3635) );
  AOI222_X0P5M_A12TR u2693 ( .A0(n2923), .A1(n3273), .B0(r201_sum_5_), .B1(
        n2924), .C0(n1107), .C1(n2982), .Y(n3632) );
  OAI21_X0P5M_A12TR u2694 ( .A0(n3636), .A1(n2908), .B0(n3637), .Y(n2632) );
  MXIT2_X0P5M_A12TR u2695 ( .A(n3638), .B(n1107), .S0(n2911), .Y(n3637) );
  OAI221_X0P5M_A12TR u2696 ( .A0(n2913), .A1(n3283), .B0(n2914), .B1(n3639), 
        .C0(n3640), .Y(n3638) );
  AOI222_X0P5M_A12TR u2697 ( .A0(r1606_sum_6_), .A1(n2917), .B0(data_in[6]), .B1(
        n2918), .C0(n241), .C1(n2919), .Y(n3640) );
  NOR2_X0P5A_A12TR u2698 ( .A(n3484), .B(state[4]), .Y(n2919) );
  NOR2_X0P5A_A12TR u2699 ( .A(state[2]), .B(u3_u93_z_6), .Y(n2918) );
  OAI31_X0P5M_A12TR u2700 ( .A0(n3641), .A1(state[4]), .A2(n3642), .B0(n30111), 
        .Y(n2917) );
  NAND3B_X0P5M_A12TR u2701 ( .AN(n2911), .B(n2826), .C(n3179), .Y(n2908) );
  OAI21_X0P5M_A12TR u2702 ( .A0(n3643), .A1(n3644), .B0(n3181), .Y(n2911) );
  OAI31_X0P5M_A12TR u2703 ( .A0(n3026), .A1(n3200), .A2(n3229), .B0(n2970), 
        .Y(n3644) );
  AOI31_X0P5M_A12TR u2704 ( .A0(n3645), .A1(n3226), .A2(n3076), .B0(n3603), 
        .Y(n2970) );
  OAI21_X0P5M_A12TR u2705 ( .A0(n3604), .A1(n3646), .B0(n3647), .Y(n3603) );
  NAND3_X0P5A_A12TR u2706 ( .A(popdes[0]), .B(n3648), .C(popdes[1]), .Y(n3647)
         );
  AOI21_X0P5M_A12TR u2707 ( .A0(n2832), .A1(n3649), .B0(state[2]), .Y(n3645)
         );
  INV_X0P5B_A12TR u2708 ( .A(carry), .Y(n2832) );
  OAI31_X0P5M_A12TR u2709 ( .A0(n3405), .A1(n3650), .A2(n3426), .B0(n3651), 
        .Y(n3643) );
  AOI31_X0P5M_A12TR u2710 ( .A0(regd[2]), .A1(regd[1]), .A2(n3652), .B0(n3653), 
        .Y(n3651) );
  OA21A1OI2_X0P5M_A12TR u2711 ( .A0(n30171), .A1(n30211), .B0(n3654), .C0(
        n3304), .Y(n3652) );
  NAND2_X0P5A_A12TR u2712 ( .A(n3074), .B(u3_u93_z_6), .Y(n3654) );
  OA21A1OI2_X0P5M_A12TR u2713 ( .A0(n236), .A1(n2866), .B0(n3289), .C0(n3290), 
        .Y(n3650) );
  AOI222_X0P5M_A12TR u2714 ( .A0(n2923), .A1(n3278), .B0(r201_sum_6_), .B1(
        n2924), .C0(n2982), .C1(n1108), .Y(n3636) );
  INV_X0P5B_A12TR u2715 ( .A(n3655), .Y(n2923) );
  NAND2_X0P5A_A12TR u2716 ( .A(n3656), .B(n3657), .Y(n2631) );
  AOI22_X0P5M_A12TR u2717 ( .A0(n970), .A1(n3658), .B0(n3659), .B1(
        rdatahold[0]), .Y(n3657) );
  AOI22_X0P5M_A12TR u2718 ( .A0(n3660), .A1(regfil_7__0_), .B0(aluopra[0]), 
        .B1(n3661), .Y(n3656) );
  NAND2_X0P5A_A12TR u2719 ( .A(n3662), .B(n3663), .Y(n2630) );
  AOI22_X0P5M_A12TR u2720 ( .A0(n969), .A1(n3658), .B0(n3659), .B1(
        rdatahold[1]), .Y(n3663) );
  AOI22_X0P5M_A12TR u2721 ( .A0(n3660), .A1(n1102), .B0(aluopra[1]), .B1(n3661), .Y(n3662) );
  NAND2_X0P5A_A12TR u2722 ( .A(n3664), .B(n3665), .Y(n2629) );
  AOI22_X0P5M_A12TR u2723 ( .A0(n968), .A1(n3658), .B0(n3659), .B1(
        rdatahold[2]), .Y(n3665) );
  AOI22_X0P5M_A12TR u2724 ( .A0(n3660), .A1(n1103), .B0(aluopra[2]), .B1(n3661), .Y(n3664) );
  NAND2_X0P5A_A12TR u2725 ( .A(n3666), .B(n3667), .Y(n2628) );
  AOI22_X0P5M_A12TR u2726 ( .A0(n967), .A1(n3658), .B0(n3659), .B1(
        rdatahold[3]), .Y(n3667) );
  AOI22_X0P5M_A12TR u2727 ( .A0(n3660), .A1(n1104), .B0(aluopra[3]), .B1(n3661), .Y(n3666) );
  NAND2_X0P5A_A12TR u2728 ( .A(n3668), .B(n3669), .Y(n2627) );
  AOI22_X0P5M_A12TR u2729 ( .A0(n966), .A1(n3658), .B0(n3659), .B1(
        rdatahold[4]), .Y(n3669) );
  AOI22_X0P5M_A12TR u2730 ( .A0(n3660), .A1(n1105), .B0(aluopra[4]), .B1(n3661), .Y(n3668) );
  NAND2_X0P5A_A12TR u2731 ( .A(n3670), .B(n3671), .Y(n2626) );
  AOI22_X0P5M_A12TR u2732 ( .A0(n965), .A1(n3658), .B0(n3659), .B1(
        rdatahold[5]), .Y(n3671) );
  AOI22_X0P5M_A12TR u2733 ( .A0(n3660), .A1(n1106), .B0(aluopra[5]), .B1(n3661), .Y(n3670) );
  NAND2_X0P5A_A12TR u2734 ( .A(n3672), .B(n3673), .Y(n2625) );
  AOI22_X0P5M_A12TR u2735 ( .A0(n964), .A1(n3658), .B0(n3659), .B1(
        rdatahold[6]), .Y(n3673) );
  AOI22_X0P5M_A12TR u2736 ( .A0(n3660), .A1(n1107), .B0(aluopra[6]), .B1(n3661), .Y(n3672) );
  NAND2_X0P5A_A12TR u2737 ( .A(n3674), .B(n3675), .Y(n2624) );
  AOI22_X0P5M_A12TR u2738 ( .A0(n963), .A1(n3658), .B0(n3659), .B1(
        rdatahold[7]), .Y(n3675) );
  NOR2_X0P5A_A12TR u2739 ( .A(n3004), .B(n3661), .Y(n3659) );
  NOR2_X0P5A_A12TR u2740 ( .A(n3605), .B(n3661), .Y(n3658) );
  AOI22_X0P5M_A12TR u2741 ( .A0(n3660), .A1(n1108), .B0(aluopra[7]), .B1(n3661), .Y(n3674) );
  NOR3_X0P5A_A12TR u2742 ( .A(n3661), .B(state[0]), .C(n3227), .Y(n3660) );
  NOR2_X0P5A_A12TR u2743 ( .A(n3366), .B(n3122), .Y(n3227) );
  AOI31_X0P5M_A12TR u2744 ( .A0(n3135), .A1(n3282), .A2(n3076), .B0(n3303), 
        .Y(n3661) );
  AOI21_X0P5M_A12TR u2745 ( .A0(n3297), .A1(n3380), .B0(n3298), .Y(n3303) );
  AOI21_X0P5M_A12TR u2746 ( .A0(n3127), .A1(n3037), .B0(n3122), .Y(n3380) );
  INV_X0P5B_A12TR u2747 ( .A(n3111), .Y(n3122) );
  INV_X0P5B_A12TR u2748 ( .A(n3317), .Y(n3282) );
  NAND2_X0P5A_A12TR u2749 ( .A(state[2]), .B(n3181), .Y(n3317) );
  INV_X0P5B_A12TR u2750 ( .A(n2913), .Y(n3135) );
  OAI222_X0P5M_A12TR u2751 ( .A0(n3251), .A1(n3676), .B0(n3611), .B1(n3677), 
        .C0(n3678), .C1(n3679), .Y(n2623) );
  INV_X0P5B_A12TR u2752 ( .A(regfil_6__0_), .Y(n3679) );
  OAI222_X0P5M_A12TR u2753 ( .A0(n3255), .A1(n3676), .B0(n3616), .B1(n3677), 
        .C0(n3678), .C1(n3680), .Y(n2622) );
  INV_X0P5B_A12TR u2754 ( .A(regfil_6__1_), .Y(n3680) );
  OAI222_X0P5M_A12TR u2755 ( .A0(n3260), .A1(n3676), .B0(n3621), .B1(n3677), 
        .C0(n3678), .C1(n3681), .Y(n2621) );
  INV_X0P5B_A12TR u2756 ( .A(regfil_6__2_), .Y(n3681) );
  OAI222_X0P5M_A12TR u2757 ( .A0(n3265), .A1(n3676), .B0(n3447), .B1(n3677), 
        .C0(n3678), .C1(n3682), .Y(n2620) );
  INV_X0P5B_A12TR u2758 ( .A(regfil_6__3_), .Y(n3682) );
  OAI222_X0P5M_A12TR u2759 ( .A0(n3270), .A1(n3676), .B0(n3630), .B1(n3677), 
        .C0(n3678), .C1(n3683), .Y(n2619) );
  INV_X0P5B_A12TR u2760 ( .A(regfil_6__4_), .Y(n3683) );
  OAI222_X0P5M_A12TR u2761 ( .A0(n3275), .A1(n3676), .B0(n3470), .B1(n3677), 
        .C0(n3678), .C1(n3684), .Y(n2618) );
  INV_X0P5B_A12TR u2762 ( .A(regfil_6__5_), .Y(n3684) );
  OAI222_X0P5M_A12TR u2763 ( .A0(n3283), .A1(n3676), .B0(n3639), .B1(n3677), 
        .C0(n3678), .C1(n3685), .Y(n2617) );
  INV_X0P5B_A12TR u2764 ( .A(regfil_6__6_), .Y(n3685) );
  OAI222_X0P5M_A12TR u2765 ( .A0(n2912), .A1(n3676), .B0(n2915), .B1(n3677), 
        .C0(n3678), .C1(n3686), .Y(n2616) );
  INV_X0P5B_A12TR u2766 ( .A(regfil_6__7_), .Y(n3686) );
  NAND2_X0P5A_A12TR u2767 ( .A(n3678), .B(u3_u93_z_6), .Y(n3677) );
  NAND2_X0P5A_A12TR u2768 ( .A(n3678), .B(state[4]), .Y(n3676) );
  NOR3_X0P5A_A12TR u2769 ( .A(n3309), .B(reset), .C(n3687), .Y(n3678) );
  OAI221_X0P5M_A12TR u2770 ( .A0(n3611), .A1(n3688), .B0(n3689), .B1(n3690), 
        .C0(n3691), .Y(n2615) );
  MXIT2_X0P5M_A12TR u2771 ( .A(n1150), .B(n3692), .S0(n3693), .Y(n3691) );
  AOI221_X0P5M_A12TR u2772 ( .A0(n1318), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_0_), .C0(n3696), .Y(n3689) );
  OAI22_X0P5M_A12TR u2773 ( .A0(n3193), .A1(n3697), .B0(n3228), .B1(n35741), 
        .Y(n3696) );
  OAI221_X0P5M_A12TR u2774 ( .A0(n3616), .A1(n3688), .B0(n3698), .B1(n3690), 
        .C0(n3699), .Y(n2614) );
  MXIT2_X0P5M_A12TR u2775 ( .A(n1151), .B(n3700), .S0(n3693), .Y(n3699) );
  AOI221_X0P5M_A12TR u2776 ( .A0(n1319), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_1_), .C0(n3701), .Y(n3698) );
  OAI22_X0P5M_A12TR u2777 ( .A0(n3193), .A1(n3702), .B0(n3228), .B1(n3579), 
        .Y(n3701) );
  OAI221_X0P5M_A12TR u2778 ( .A0(n3621), .A1(n3688), .B0(n3703), .B1(n3690), 
        .C0(n3704), .Y(n2613) );
  MXIT2_X0P5M_A12TR u2779 ( .A(n1152), .B(n3705), .S0(n3693), .Y(n3704) );
  AOI221_X0P5M_A12TR u2780 ( .A0(n1320), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_2_), .C0(n3706), .Y(n3703) );
  OAI22_X0P5M_A12TR u2781 ( .A0(n3193), .A1(n3707), .B0(n3228), .B1(n3580), 
        .Y(n3706) );
  OAI221_X0P5M_A12TR u2782 ( .A0(n3447), .A1(n3688), .B0(n3708), .B1(n3690), 
        .C0(n3709), .Y(n2612) );
  MXIT2_X0P5M_A12TR u2783 ( .A(n1153), .B(n3710), .S0(n3693), .Y(n3709) );
  AOI221_X0P5M_A12TR u2784 ( .A0(n1321), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_3_), .C0(n3711), .Y(n3708) );
  OAI22_X0P5M_A12TR u2785 ( .A0(n3193), .A1(n3712), .B0(n3228), .B1(n3581), 
        .Y(n3711) );
  OAI221_X0P5M_A12TR u2786 ( .A0(n3630), .A1(n3688), .B0(n3713), .B1(n3690), 
        .C0(n3714), .Y(n2611) );
  MXIT2_X0P5M_A12TR u2787 ( .A(n1154), .B(n3715), .S0(n3693), .Y(n3714) );
  AOI221_X0P5M_A12TR u2788 ( .A0(n1322), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_4_), .C0(n3716), .Y(n3713) );
  OAI22_X0P5M_A12TR u2789 ( .A0(n3193), .A1(n3717), .B0(n3228), .B1(n3582), 
        .Y(n3716) );
  OAI221_X0P5M_A12TR u2790 ( .A0(n3470), .A1(n3688), .B0(n3718), .B1(n3690), 
        .C0(n3719), .Y(n2610) );
  MXIT2_X0P5M_A12TR u2791 ( .A(n1155), .B(n3720), .S0(n3693), .Y(n3719) );
  AOI221_X0P5M_A12TR u2792 ( .A0(n1323), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_5_), .C0(n3721), .Y(n3718) );
  OAI22_X0P5M_A12TR u2793 ( .A0(n3193), .A1(n3722), .B0(n3228), .B1(n3583), 
        .Y(n3721) );
  OAI221_X0P5M_A12TR u2794 ( .A0(n3639), .A1(n3688), .B0(n3723), .B1(n3690), 
        .C0(n3724), .Y(n2609) );
  MXIT2_X0P5M_A12TR u2795 ( .A(n1156), .B(n3725), .S0(n3693), .Y(n3724) );
  AOI221_X0P5M_A12TR u2796 ( .A0(n1324), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_6_), .C0(n3726), .Y(n3723) );
  OAI22_X0P5M_A12TR u2797 ( .A0(n3193), .A1(n3727), .B0(n3228), .B1(n3584), 
        .Y(n3726) );
  OAI221_X0P5M_A12TR u2798 ( .A0(n2915), .A1(n3688), .B0(n3728), .B1(n3690), 
        .C0(n3729), .Y(n2608) );
  MXIT2_X0P5M_A12TR u2799 ( .A(n1157), .B(n3597), .S0(n3693), .Y(n3729) );
  OAI22_X0P5M_A12TR u2800 ( .A0(n3167), .A1(n3236), .B0(n2912), .B1(n3730), 
        .Y(n3597) );
  INV_X0P5B_A12TR u2801 ( .A(rdatahold2[7]), .Y(n3236) );
  NAND3_X0P5A_A12TR u2802 ( .A(n3004), .B(n3153), .C(n3693), .Y(n3690) );
  AOI221_X0P5M_A12TR u2803 ( .A0(n1325), .A1(n3694), .B0(n3695), .B1(
        r1606_sum_7_), .C0(n3731), .Y(n3728) );
  OAI22_X0P5M_A12TR u2804 ( .A0(n3193), .A1(n3732), .B0(n3228), .B1(n3585), 
        .Y(n3731) );
  NAND2_X0P5A_A12TR u2805 ( .A(n3073), .B(n3693), .Y(n3688) );
  OAI21_X0P5M_A12TR u2806 ( .A0(reset), .A1(n3733), .B0(n3734), .Y(n3693) );
  AOI32_X0P5M_A12TR u2807 ( .A0(regd[2]), .A1(regd[0]), .A2(n3735), .B0(n3736), 
        .B1(n3196), .Y(n3734) );
  OAI221_X0P5M_A12TR u2808 ( .A0(n3737), .A1(n3738), .B0(n3611), .B1(n3739), 
        .C0(n3740), .Y(n2607) );
  AOI22_X0P5M_A12TR u2809 ( .A0(n3741), .A1(rdatahold[0]), .B0(n3742), .B1(
        n1158), .Y(n3740) );
  AOI221_X0P5M_A12TR u2810 ( .A0(n1326), .A1(n3694), .B0(n3695), .B1(
        r201_sum_8_), .C0(n3743), .Y(n3737) );
  AO22_X0P5M_A12TR u2811 ( .A0(n3366), .A1(regfil_2__0_), .B0(n35711), .B1(
        n247), .Y(n3743) );
  OAI221_X0P5M_A12TR u2812 ( .A0(n3744), .A1(n3738), .B0(n3616), .B1(n3739), 
        .C0(n3745), .Y(n2606) );
  AOI22_X0P5M_A12TR u2813 ( .A0(n3741), .A1(rdatahold[1]), .B0(n3742), .B1(
        n1159), .Y(n3745) );
  AOI221_X0P5M_A12TR u2814 ( .A0(n1327), .A1(n3694), .B0(n3695), .B1(
        r201_sum_9_), .C0(n3746), .Y(n3744) );
  AO22_X0P5M_A12TR u2815 ( .A0(n3366), .A1(regfil_2__1_), .B0(n35711), .B1(
        n246), .Y(n3746) );
  OAI221_X0P5M_A12TR u2816 ( .A0(n3747), .A1(n3738), .B0(n3621), .B1(n3739), 
        .C0(n3748), .Y(n2605) );
  AOI22_X0P5M_A12TR u2817 ( .A0(n3741), .A1(rdatahold[2]), .B0(n3742), .B1(
        n1160), .Y(n3748) );
  AOI221_X0P5M_A12TR u2818 ( .A0(n1328), .A1(n3694), .B0(n3695), .B1(
        r201_sum_10_), .C0(n3749), .Y(n3747) );
  AO22_X0P5M_A12TR u2819 ( .A0(n3366), .A1(regfil_2__2_), .B0(n35711), .B1(
        n245), .Y(n3749) );
  OAI221_X0P5M_A12TR u2820 ( .A0(n3750), .A1(n3738), .B0(n3447), .B1(n3739), 
        .C0(n3751), .Y(n2604) );
  AOI22_X0P5M_A12TR u2821 ( .A0(n3741), .A1(rdatahold[3]), .B0(n3742), .B1(
        n1161), .Y(n3751) );
  AOI221_X0P5M_A12TR u2822 ( .A0(n1329), .A1(n3694), .B0(n3695), .B1(
        r201_sum_11_), .C0(n3752), .Y(n3750) );
  AO22_X0P5M_A12TR u2823 ( .A0(n3366), .A1(regfil_2__3_), .B0(n35711), .B1(
        n244), .Y(n3752) );
  OAI221_X0P5M_A12TR u2824 ( .A0(n3753), .A1(n3738), .B0(n3630), .B1(n3739), 
        .C0(n3754), .Y(n2603) );
  AOI22_X0P5M_A12TR u2825 ( .A0(n3741), .A1(rdatahold[4]), .B0(n3742), .B1(
        n1162), .Y(n3754) );
  AOI221_X0P5M_A12TR u2826 ( .A0(n1330), .A1(n3694), .B0(n3695), .B1(
        r201_sum_12_), .C0(n3755), .Y(n3753) );
  AO22_X0P5M_A12TR u2827 ( .A0(n3366), .A1(regfil_2__4_), .B0(n35711), .B1(
        n243), .Y(n3755) );
  OAI221_X0P5M_A12TR u2828 ( .A0(n3756), .A1(n3738), .B0(n3470), .B1(n3739), 
        .C0(n3757), .Y(n2602) );
  AOI22_X0P5M_A12TR u2829 ( .A0(n3741), .A1(rdatahold[5]), .B0(n3742), .B1(
        n1163), .Y(n3757) );
  AOI221_X0P5M_A12TR u2830 ( .A0(n1331), .A1(n3694), .B0(n3695), .B1(
        r201_sum_13_), .C0(n3758), .Y(n3756) );
  AO22_X0P5M_A12TR u2831 ( .A0(n3366), .A1(regfil_2__5_), .B0(n35711), .B1(
        n242), .Y(n3758) );
  OAI221_X0P5M_A12TR u2832 ( .A0(n3759), .A1(n3738), .B0(n3639), .B1(n3739), 
        .C0(n3760), .Y(n2601) );
  AOI22_X0P5M_A12TR u2833 ( .A0(n3741), .A1(rdatahold[6]), .B0(n3742), .B1(
        n1164), .Y(n3760) );
  AOI221_X0P5M_A12TR u2834 ( .A0(n1332), .A1(n3694), .B0(n3695), .B1(
        r201_sum_14_), .C0(n3761), .Y(n3759) );
  AO22_X0P5M_A12TR u2835 ( .A0(n3366), .A1(regfil_2__6_), .B0(n35711), .B1(
        n241), .Y(n3761) );
  OAI221_X0P5M_A12TR u2836 ( .A0(n3762), .A1(n3738), .B0(n2915), .B1(n3739), 
        .C0(n3763), .Y(n2600) );
  AOI22_X0P5M_A12TR u2837 ( .A0(n3741), .A1(rdatahold[7]), .B0(n3742), .B1(
        n1165), .Y(n3763) );
  AOI21_X0P5M_A12TR u2838 ( .A0(n30141), .A1(n2913), .B0(n3742), .Y(n3741) );
  INV_X0P5B_A12TR u2839 ( .A(n3764), .Y(n3742) );
  NAND2_X0P5A_A12TR u2840 ( .A(state[0]), .B(n2823), .Y(n2913) );
  NAND2_X0P5A_A12TR u2841 ( .A(n3073), .B(n3764), .Y(n3739) );
  INV_X0P5B_A12TR u2842 ( .A(n3294), .Y(n3073) );
  NAND3_X0P5A_A12TR u2843 ( .A(n3004), .B(n3153), .C(n3764), .Y(n3738) );
  OAI21_X0P5M_A12TR u2844 ( .A0(reset), .A1(n3733), .B0(n3765), .Y(n3764) );
  AOI32_X0P5M_A12TR u2845 ( .A0(regd[2]), .A1(n3304), .A2(n3735), .B0(n3736), 
        .B1(n3766), .Y(n3765) );
  OA211_X0P5M_A12TR u2846 ( .A0(n3767), .A1(n3405), .B0(n3768), .C0(n3769), 
        .Y(n3733) );
  AOI31_X0P5M_A12TR u2847 ( .A0(n3648), .A1(n3313), .A2(popdes[1]), .B0(n3770), 
        .Y(n3769) );
  OAI21_X0P5M_A12TR u2848 ( .A0(n3078), .A1(n3212), .B0(n2894), .Y(n3768) );
  INV_X0P5B_A12TR u2849 ( .A(n3168), .Y(n3212) );
  NOR2_X0P5A_A12TR u2850 ( .A(n2981), .B(n3771), .Y(n3767) );
  AOI221_X0P5M_A12TR u2851 ( .A0(n1333), .A1(n3694), .B0(n3695), .B1(
        r201_sum_15_), .C0(n3772), .Y(n3762) );
  AO22_X0P5M_A12TR u2852 ( .A0(n3366), .A1(regfil_2__7_), .B0(n35711), .B1(
        n240), .Y(n3772) );
  INV_X0P5B_A12TR u2853 ( .A(n3773), .Y(n3695) );
  NOR2B_X0P5M_A12TR u2854 ( .AN(n2981), .B(n3036), .Y(n3694) );
  MXIT2_X0P5M_A12TR u2855 ( .A(n3774), .B(n3697), .S0(n3775), .Y(n2599) );
  INV_X0P5B_A12TR u2856 ( .A(n1657), .Y(n3697) );
  AOI211_X0P5M_A12TR u2857 ( .A0(rdatahold2[0]), .A1(n3087), .B0(n3776), .C0(
        n3777), .Y(n3774) );
  OAI222_X0P5M_A12TR u2858 ( .A0(n3605), .A1(n3778), .B0(n3251), .B1(n3230), 
        .C0(n3409), .C1(n2961), .Y(n3776) );
  INV_X0P5B_A12TR u2859 ( .A(r1606_sum_0_), .Y(n3778) );
  MXIT2_X0P5M_A12TR u2860 ( .A(n3779), .B(n3702), .S0(n3775), .Y(n2598) );
  INV_X0P5B_A12TR u2861 ( .A(n1658), .Y(n3702) );
  AOI211_X0P5M_A12TR u2862 ( .A0(rdatahold2[1]), .A1(n3087), .B0(n3780), .C0(
        n3781), .Y(n3779) );
  OAI222_X0P5M_A12TR u2863 ( .A0(n3605), .A1(n3782), .B0(n3255), .B1(n3230), 
        .C0(n2961), .C1(n3420), .Y(n3780) );
  INV_X0P5B_A12TR u2864 ( .A(r1606_sum_1_), .Y(n3782) );
  MXIT2_X0P5M_A12TR u2865 ( .A(n3783), .B(n3707), .S0(n3775), .Y(n2597) );
  INV_X0P5B_A12TR u2866 ( .A(n1659), .Y(n3707) );
  AOI211_X0P5M_A12TR u2867 ( .A0(rdatahold2[2]), .A1(n3087), .B0(n3784), .C0(
        n3785), .Y(n3783) );
  OAI222_X0P5M_A12TR u2868 ( .A0(n3605), .A1(n3786), .B0(n3260), .B1(n3230), 
        .C0(n2961), .C1(n3434), .Y(n3784) );
  INV_X0P5B_A12TR u2869 ( .A(r1606_sum_2_), .Y(n3786) );
  MXIT2_X0P5M_A12TR u2870 ( .A(n3787), .B(n3712), .S0(n3775), .Y(n2596) );
  INV_X0P5B_A12TR u2871 ( .A(n1660), .Y(n3712) );
  AOI211_X0P5M_A12TR u2872 ( .A0(rdatahold2[3]), .A1(n3087), .B0(n3788), .C0(
        n3789), .Y(n3787) );
  OAI222_X0P5M_A12TR u2873 ( .A0(n3605), .A1(n3790), .B0(n3265), .B1(n3230), 
        .C0(n2961), .C1(n3443), .Y(n3788) );
  INV_X0P5B_A12TR u2874 ( .A(r1606_sum_3_), .Y(n3790) );
  MXIT2_X0P5M_A12TR u2875 ( .A(n3791), .B(n3717), .S0(n3775), .Y(n2595) );
  INV_X0P5B_A12TR u2876 ( .A(n1661), .Y(n3717) );
  AOI211_X0P5M_A12TR u2877 ( .A0(rdatahold2[4]), .A1(n3087), .B0(n3792), .C0(
        n3793), .Y(n3791) );
  OAI222_X0P5M_A12TR u2878 ( .A0(n3605), .A1(n3794), .B0(n3270), .B1(n3230), 
        .C0(n2961), .C1(n3458), .Y(n3792) );
  INV_X0P5B_A12TR u2879 ( .A(r1606_sum_4_), .Y(n3794) );
  MXIT2_X0P5M_A12TR u2880 ( .A(n3795), .B(n3722), .S0(n3775), .Y(n2594) );
  INV_X0P5B_A12TR u2881 ( .A(n1662), .Y(n3722) );
  AOI211_X0P5M_A12TR u2882 ( .A0(rdatahold2[5]), .A1(n3087), .B0(n3796), .C0(
        n3797), .Y(n3795) );
  OAI222_X0P5M_A12TR u2883 ( .A0(n3605), .A1(n3798), .B0(n3275), .B1(n3230), 
        .C0(n2961), .C1(n3466), .Y(n3796) );
  INV_X0P5B_A12TR u2884 ( .A(r1606_sum_5_), .Y(n3798) );
  MXIT2_X0P5M_A12TR u2885 ( .A(n3799), .B(n3727), .S0(n3775), .Y(n2593) );
  INV_X0P5B_A12TR u2886 ( .A(n1663), .Y(n3727) );
  AOI211_X0P5M_A12TR u2887 ( .A0(rdatahold2[6]), .A1(n3087), .B0(n3800), .C0(
        n3801), .Y(n3799) );
  OAI222_X0P5M_A12TR u2888 ( .A0(n3605), .A1(n3802), .B0(n3283), .B1(n3230), 
        .C0(n2961), .C1(n3481), .Y(n3800) );
  INV_X0P5B_A12TR u2889 ( .A(r1606_sum_6_), .Y(n3802) );
  MXIT2_X0P5M_A12TR u2890 ( .A(n3803), .B(n3732), .S0(n3775), .Y(n2592) );
  OAI21_X0P5M_A12TR u2891 ( .A0(n3804), .A1(n3805), .B0(n3181), .Y(n3775) );
  OAI31_X0P5M_A12TR u2892 ( .A0(n3197), .A1(n3229), .A2(n3026), .B0(n3806), 
        .Y(n3805) );
  NAND4_X0P5A_A12TR u2893 ( .A(regd[1]), .B(regd[0]), .C(n3807), .D(n3309), 
        .Y(n3806) );
  INV_X0P5B_A12TR u2894 ( .A(n1664), .Y(n3732) );
  AOI211_X0P5M_A12TR u2895 ( .A0(rdatahold2[7]), .A1(n3087), .B0(n3808), .C0(
        n2964), .Y(n3803) );
  OAI22_X0P5M_A12TR u2896 ( .A0(n2823), .A1(n2915), .B0(n3585), .B1(n3809), 
        .Y(n2964) );
  INV_X0P5B_A12TR u2897 ( .A(n240), .Y(n3585) );
  INV_X0P5B_A12TR u2898 ( .A(alures[7]), .Y(n2915) );
  OAI222_X0P5M_A12TR u2899 ( .A0(n3810), .A1(n3605), .B0(n2912), .B1(n3230), 
        .C0(n2889), .C1(n2961), .Y(n3808) );
  NAND2_X0P5A_A12TR u2900 ( .A(state[3]), .B(state[2]), .Y(n3230) );
  INV_X0P5B_A12TR u2901 ( .A(r1606_sum_7_), .Y(n3810) );
  OAI221_X0P5M_A12TR u2902 ( .A0(n2954), .A1(n2978), .B0(n2956), .B1(n3811), 
        .C0(n3812), .Y(n2591) );
  MXIT2_X0P5M_A12TR u2903 ( .A(regfil_2__0_), .B(n3813), .S0(n2959), .Y(n3812)
         );
  OAI221_X0P5M_A12TR u2904 ( .A0(n2871), .A1(n2961), .B0(n2962), .B1(n3251), 
        .C0(n3814), .Y(n3813) );
  INV_X0P5B_A12TR u2905 ( .A(n3777), .Y(n3814) );
  OAI22_X0P5M_A12TR u2906 ( .A0(n2823), .A1(n3611), .B0(n3809), .B1(n35741), 
        .Y(n3777) );
  INV_X0P5B_A12TR u2907 ( .A(r194_sum_8_), .Y(n3811) );
  INV_X0P5B_A12TR u2908 ( .A(r201_sum_8_), .Y(n2978) );
  OAI221_X0P5M_A12TR u2909 ( .A0(n2954), .A1(n3815), .B0(n2956), .B1(n3816), 
        .C0(n3817), .Y(n2590) );
  MXIT2_X0P5M_A12TR u2910 ( .A(regfil_2__1_), .B(n3818), .S0(n2959), .Y(n3817)
         );
  OAI221_X0P5M_A12TR u2911 ( .A0(n3819), .A1(n2961), .B0(n2962), .B1(n3255), 
        .C0(n3820), .Y(n3818) );
  INV_X0P5B_A12TR u2912 ( .A(n3781), .Y(n3820) );
  OAI22_X0P5M_A12TR u2913 ( .A0(n2823), .A1(n3616), .B0(n3809), .B1(n3579), 
        .Y(n3781) );
  INV_X0P5B_A12TR u2914 ( .A(r194_sum_9_), .Y(n3816) );
  INV_X0P5B_A12TR u2915 ( .A(r201_sum_9_), .Y(n3815) );
  OAI221_X0P5M_A12TR u2916 ( .A0(n2954), .A1(n3821), .B0(n2956), .B1(n3822), 
        .C0(n3823), .Y(n2589) );
  MXIT2_X0P5M_A12TR u2917 ( .A(regfil_2__2_), .B(n3824), .S0(n2959), .Y(n3823)
         );
  OAI221_X0P5M_A12TR u2918 ( .A0(n3825), .A1(n2961), .B0(n2962), .B1(n3260), 
        .C0(n3826), .Y(n3824) );
  INV_X0P5B_A12TR u2919 ( .A(n3785), .Y(n3826) );
  OAI22_X0P5M_A12TR u2920 ( .A0(n2823), .A1(n3621), .B0(n3809), .B1(n3580), 
        .Y(n3785) );
  INV_X0P5B_A12TR u2921 ( .A(r194_sum_10_), .Y(n3822) );
  INV_X0P5B_A12TR u2922 ( .A(r201_sum_10_), .Y(n3821) );
  OAI221_X0P5M_A12TR u2923 ( .A0(n2954), .A1(n3827), .B0(n2956), .B1(n3828), 
        .C0(n3829), .Y(n2588) );
  MXIT2_X0P5M_A12TR u2924 ( .A(regfil_2__3_), .B(n3830), .S0(n2959), .Y(n3829)
         );
  OAI221_X0P5M_A12TR u2925 ( .A0(n3831), .A1(n2961), .B0(n2962), .B1(n3265), 
        .C0(n3832), .Y(n3830) );
  INV_X0P5B_A12TR u2926 ( .A(n3789), .Y(n3832) );
  OAI22_X0P5M_A12TR u2927 ( .A0(n2823), .A1(n3447), .B0(n3809), .B1(n3581), 
        .Y(n3789) );
  INV_X0P5B_A12TR u2928 ( .A(r194_sum_11_), .Y(n3828) );
  INV_X0P5B_A12TR u2929 ( .A(r201_sum_11_), .Y(n3827) );
  OAI221_X0P5M_A12TR u2930 ( .A0(n2954), .A1(n3833), .B0(n2956), .B1(n3834), 
        .C0(n3835), .Y(n2587) );
  MXIT2_X0P5M_A12TR u2931 ( .A(regfil_2__4_), .B(n3836), .S0(n2959), .Y(n3835)
         );
  OAI221_X0P5M_A12TR u2932 ( .A0(n3837), .A1(n2961), .B0(n2962), .B1(n3270), 
        .C0(n3838), .Y(n3836) );
  INV_X0P5B_A12TR u2933 ( .A(n3793), .Y(n3838) );
  OAI22_X0P5M_A12TR u2934 ( .A0(n2823), .A1(n3630), .B0(n3809), .B1(n3582), 
        .Y(n3793) );
  INV_X0P5B_A12TR u2935 ( .A(r194_sum_12_), .Y(n3834) );
  INV_X0P5B_A12TR u2936 ( .A(r201_sum_12_), .Y(n3833) );
  OAI221_X0P5M_A12TR u2937 ( .A0(n2954), .A1(n3839), .B0(n2956), .B1(n3840), 
        .C0(n3841), .Y(n2586) );
  MXIT2_X0P5M_A12TR u2938 ( .A(regfil_2__5_), .B(n3842), .S0(n2959), .Y(n3841)
         );
  OAI221_X0P5M_A12TR u2939 ( .A0(n3843), .A1(n2961), .B0(n2962), .B1(n3275), 
        .C0(n3844), .Y(n3842) );
  INV_X0P5B_A12TR u2940 ( .A(n3797), .Y(n3844) );
  OAI22_X0P5M_A12TR u2941 ( .A0(n2823), .A1(n3470), .B0(n3809), .B1(n3583), 
        .Y(n3797) );
  INV_X0P5B_A12TR u2942 ( .A(r194_sum_13_), .Y(n3840) );
  INV_X0P5B_A12TR u2943 ( .A(r201_sum_13_), .Y(n3839) );
  OAI221_X0P5M_A12TR u2944 ( .A0(n2954), .A1(n3845), .B0(n2956), .B1(n3846), 
        .C0(n3847), .Y(n2585) );
  MXIT2_X0P5M_A12TR u2945 ( .A(regfil_2__6_), .B(n3848), .S0(n2959), .Y(n3847)
         );
  OAI221_X0P5M_A12TR u2946 ( .A0(n3849), .A1(n2961), .B0(n2962), .B1(n3283), 
        .C0(n3850), .Y(n3848) );
  INV_X0P5B_A12TR u2947 ( .A(n3801), .Y(n3850) );
  OAI22_X0P5M_A12TR u2948 ( .A0(n2823), .A1(n3639), .B0(n3809), .B1(n3584), 
        .Y(n3801) );
  NAND2_X0P5A_A12TR u2949 ( .A(n35711), .B(n3004), .Y(n3809) );
  NOR2_X0P5A_A12TR u2950 ( .A(n2972), .B(state[4]), .Y(n2962) );
  NAND2_X0P5A_A12TR u2951 ( .A(n3366), .B(n3004), .Y(n2961) );
  INV_X0P5B_A12TR u2952 ( .A(r194_sum_14_), .Y(n3846) );
  NAND3_X0P5A_A12TR u2953 ( .A(n2959), .B(n3350), .C(n3851), .Y(n2956) );
  INV_X0P5B_A12TR u2954 ( .A(r201_sum_14_), .Y(n3845) );
  NAND3_X0P5A_A12TR u2955 ( .A(n2959), .B(n3852), .C(n3851), .Y(n2954) );
  INV_X0P5B_A12TR u2956 ( .A(n3605), .Y(n3851) );
  NAND2_X0P5A_A12TR u2957 ( .A(n3127), .B(n3004), .Y(n3605) );
  OA21_X0P5M_A12TR u2958 ( .A0(n3804), .A1(n3853), .B0(n3181), .Y(n2959) );
  OAI21_X0P5M_A12TR u2959 ( .A0(regd[2]), .A1(n3687), .B0(n3854), .Y(n3853) );
  NAND4B_X0P5M_A12TR u2960 ( .AN(n3026), .B(n3855), .C(n3204), .D(n2828), .Y(
        n3854) );
  NAND3_X0P5A_A12TR u2961 ( .A(n3807), .B(n3304), .C(regd[1]), .Y(n3687) );
  INV_X0P5B_A12TR u2962 ( .A(regd[0]), .Y(n3304) );
  OAI221_X0P5M_A12TR u2963 ( .A0(n3375), .A1(n3405), .B0(n30141), .B1(n3166), 
        .C0(n3856), .Y(n3804) );
  AOI31_X0P5M_A12TR u2964 ( .A0(n3648), .A1(n3315), .A2(popdes[0]), .B0(n3770), 
        .Y(n3856) );
  NOR3_X0P5A_A12TR u2965 ( .A(n3042), .B(n3857), .C(n3329), .Y(n3770) );
  MXIT2_X0P5M_A12TR u2966 ( .A(n3858), .B(n3859), .S0(n3596), .Y(n2584) );
  AOI211_X0P5M_A12TR u2967 ( .A0(r1606_sum_0_), .A1(n2928), .B0(n3692), .C0(
        n3860), .Y(n3859) );
  OAI22_X0P5M_A12TR u2968 ( .A0(n3167), .A1(n2975), .B0(n3251), .B1(n3730), 
        .Y(n3692) );
  MXIT2_X0P5M_A12TR u2969 ( .A(n3861), .B(n3862), .S0(n3596), .Y(n2583) );
  AOI211_X0P5M_A12TR u2970 ( .A0(r1606_sum_1_), .A1(n2928), .B0(n3700), .C0(
        n3863), .Y(n3862) );
  OAI22_X0P5M_A12TR u2971 ( .A0(n3167), .A1(n3257), .B0(n3255), .B1(n3730), 
        .Y(n3700) );
  INV_X0P5B_A12TR u2972 ( .A(rdatahold2[1]), .Y(n3257) );
  MXIT2_X0P5M_A12TR u2973 ( .A(n3864), .B(n3865), .S0(n3596), .Y(n2582) );
  AOI211_X0P5M_A12TR u2974 ( .A0(r1606_sum_2_), .A1(n2928), .B0(n3705), .C0(
        n3866), .Y(n3865) );
  OAI22_X0P5M_A12TR u2975 ( .A0(n3167), .A1(n3262), .B0(n3260), .B1(n3730), 
        .Y(n3705) );
  INV_X0P5B_A12TR u2976 ( .A(rdatahold2[2]), .Y(n3262) );
  MXIT2_X0P5M_A12TR u2977 ( .A(n3867), .B(n3868), .S0(n3596), .Y(n2581) );
  AOI211_X0P5M_A12TR u2978 ( .A0(r1606_sum_3_), .A1(n2928), .B0(n3710), .C0(
        n3869), .Y(n3868) );
  OAI22_X0P5M_A12TR u2979 ( .A0(n3167), .A1(n3267), .B0(n3265), .B1(n3730), 
        .Y(n3710) );
  INV_X0P5B_A12TR u2980 ( .A(rdatahold2[3]), .Y(n3267) );
  MXIT2_X0P5M_A12TR u2981 ( .A(n3870), .B(n3871), .S0(n3596), .Y(n2580) );
  AOI211_X0P5M_A12TR u2982 ( .A0(r1606_sum_4_), .A1(n2928), .B0(n3715), .C0(
        n3872), .Y(n3871) );
  OAI22_X0P5M_A12TR u2983 ( .A0(n3167), .A1(n3272), .B0(n3270), .B1(n3730), 
        .Y(n3715) );
  INV_X0P5B_A12TR u2984 ( .A(rdatahold2[4]), .Y(n3272) );
  MXIT2_X0P5M_A12TR u2985 ( .A(n3873), .B(n3874), .S0(n3596), .Y(n2579) );
  AOI211_X0P5M_A12TR u2986 ( .A0(r1606_sum_5_), .A1(n2928), .B0(n3720), .C0(
        n3875), .Y(n3874) );
  OAI22_X0P5M_A12TR u2987 ( .A0(n3167), .A1(n3277), .B0(n3275), .B1(n3730), 
        .Y(n3720) );
  INV_X0P5B_A12TR u2988 ( .A(rdatahold2[5]), .Y(n3277) );
  MXIT2_X0P5M_A12TR u2989 ( .A(n3876), .B(n3877), .S0(n3596), .Y(n2578) );
  OAI21_X0P5M_A12TR u2990 ( .A0(reset), .A1(n3878), .B0(n3879), .Y(n3596) );
  AOI32_X0P5M_A12TR u2991 ( .A0(regd[0]), .A1(n3309), .A2(n3735), .B0(n3736), 
        .B1(n2920), .Y(n3879) );
  INV_X0P5B_A12TR u2992 ( .A(n3880), .Y(n3735) );
  INV_X0P5B_A12TR u2993 ( .A(regd[2]), .Y(n3309) );
  AOI211_X0P5M_A12TR u2994 ( .A0(r1606_sum_6_), .A1(n2928), .B0(n3725), .C0(
        n3881), .Y(n3877) );
  OAI22_X0P5M_A12TR u2995 ( .A0(n3167), .A1(n3285), .B0(n3283), .B1(n3730), 
        .Y(n3725) );
  INV_X0P5B_A12TR u2996 ( .A(rdatahold2[6]), .Y(n3285) );
  INV_X0P5B_A12TR u2997 ( .A(n3087), .Y(n3167) );
  MXIT2_X0P5M_A12TR u2998 ( .A(n3882), .B(n3883), .S0(n2927), .Y(n2577) );
  AOI221_X0P5M_A12TR u2999 ( .A0(r201_sum_8_), .A1(n2928), .B0(rdatahold[0]), 
        .B1(n2929), .C0(n3860), .Y(n3883) );
  OAI22_X0P5M_A12TR u3000 ( .A0(n2823), .A1(n3611), .B0(n3598), .B1(n35741), 
        .Y(n3860) );
  INV_X0P5B_A12TR u3001 ( .A(n247), .Y(n35741) );
  INV_X0P5B_A12TR u3002 ( .A(alures[0]), .Y(n3611) );
  MXIT2_X0P5M_A12TR u3003 ( .A(n3884), .B(n3885), .S0(n2927), .Y(n2576) );
  AOI221_X0P5M_A12TR u3004 ( .A0(r201_sum_9_), .A1(n2928), .B0(rdatahold[1]), 
        .B1(n2929), .C0(n3863), .Y(n3885) );
  OAI22_X0P5M_A12TR u3005 ( .A0(n2823), .A1(n3616), .B0(n3598), .B1(n3579), 
        .Y(n3863) );
  INV_X0P5B_A12TR u3006 ( .A(n246), .Y(n3579) );
  INV_X0P5B_A12TR u3007 ( .A(alures[1]), .Y(n3616) );
  MXIT2_X0P5M_A12TR u3008 ( .A(n3886), .B(n3887), .S0(n2927), .Y(n2575) );
  AOI221_X0P5M_A12TR u3009 ( .A0(r201_sum_10_), .A1(n2928), .B0(rdatahold[2]), 
        .B1(n2929), .C0(n3866), .Y(n3887) );
  OAI22_X0P5M_A12TR u3010 ( .A0(n2823), .A1(n3621), .B0(n3598), .B1(n3580), 
        .Y(n3866) );
  INV_X0P5B_A12TR u3011 ( .A(n245), .Y(n3580) );
  INV_X0P5B_A12TR u3012 ( .A(alures[2]), .Y(n3621) );
  MXIT2_X0P5M_A12TR u3013 ( .A(n3888), .B(n3889), .S0(n2927), .Y(n2574) );
  AOI221_X0P5M_A12TR u3014 ( .A0(r201_sum_11_), .A1(n2928), .B0(rdatahold[3]), 
        .B1(n2929), .C0(n3869), .Y(n3889) );
  OAI22_X0P5M_A12TR u3015 ( .A0(n2823), .A1(n3447), .B0(n3598), .B1(n3581), 
        .Y(n3869) );
  INV_X0P5B_A12TR u3016 ( .A(n244), .Y(n3581) );
  INV_X0P5B_A12TR u3017 ( .A(alures[3]), .Y(n3447) );
  MXIT2_X0P5M_A12TR u3018 ( .A(n3890), .B(n3891), .S0(n2927), .Y(n2573) );
  AOI221_X0P5M_A12TR u3019 ( .A0(r201_sum_12_), .A1(n2928), .B0(rdatahold[4]), 
        .B1(n2929), .C0(n3872), .Y(n3891) );
  OAI22_X0P5M_A12TR u3020 ( .A0(n2823), .A1(n3630), .B0(n3598), .B1(n3582), 
        .Y(n3872) );
  INV_X0P5B_A12TR u3021 ( .A(n243), .Y(n3582) );
  INV_X0P5B_A12TR u3022 ( .A(alures[4]), .Y(n3630) );
  MXIT2_X0P5M_A12TR u3023 ( .A(n3892), .B(n3893), .S0(n2927), .Y(n2572) );
  AOI221_X0P5M_A12TR u3024 ( .A0(r201_sum_13_), .A1(n2928), .B0(rdatahold[5]), 
        .B1(n2929), .C0(n3875), .Y(n3893) );
  OAI22_X0P5M_A12TR u3025 ( .A0(n2823), .A1(n3470), .B0(n3598), .B1(n3583), 
        .Y(n3875) );
  INV_X0P5B_A12TR u3026 ( .A(n242), .Y(n3583) );
  INV_X0P5B_A12TR u3027 ( .A(alures[5]), .Y(n3470) );
  MXIT2_X0P5M_A12TR u3028 ( .A(n3894), .B(n3895), .S0(n2927), .Y(n2571) );
  OAI21_X0P5M_A12TR u3029 ( .A0(reset), .A1(n3878), .B0(n3896), .Y(n2927) );
  AOI31_X0P5M_A12TR u3030 ( .A0(n3203), .A1(n2828), .A2(n3736), .B0(n3897), 
        .Y(n3896) );
  NOR3_X0P5A_A12TR u3031 ( .A(n3880), .B(regd[2]), .C(regd[0]), .Y(n3897) );
  NAND3_X0P5A_A12TR u3032 ( .A(n3306), .B(n3181), .C(n3807), .Y(n3880) );
  OAI22_X0P5M_A12TR u3033 ( .A0(n30171), .A1(n30211), .B0(n3604), .B1(n3294), 
        .Y(n3807) );
  NAND2_X0P5A_A12TR u3034 ( .A(state[0]), .B(u3_u93_z_6), .Y(n3294) );
  INV_X0P5B_A12TR u3035 ( .A(regd[1]), .Y(n3306) );
  NOR2_X0P5A_A12TR u3036 ( .A(n3026), .B(n3298), .Y(n3736) );
  NAND3_X0P5A_A12TR u3037 ( .A(n3038), .B(n3123), .C(n35711), .Y(n3026) );
  AOI21B_X0P5M_A12TR u3038 ( .A0(n2894), .A1(n3241), .B0N(n3898), .Y(n3878) );
  AOI32_X0P5M_A12TR u3039 ( .A0(n3313), .A1(n3315), .A2(n3648), .B0(n2989), 
        .B1(n3899), .Y(n3898) );
  INV_X0P5B_A12TR u3040 ( .A(n3405), .Y(n2989) );
  NOR2_X0P5A_A12TR u3041 ( .A(n30211), .B(n3086), .Y(n3648) );
  INV_X0P5B_A12TR u3042 ( .A(popdes[1]), .Y(n3315) );
  INV_X0P5B_A12TR u3043 ( .A(popdes[0]), .Y(n3313) );
  AOI221_X0P5M_A12TR u3044 ( .A0(r201_sum_14_), .A1(n2928), .B0(rdatahold[6]), 
        .B1(n2929), .C0(n3881), .Y(n3895) );
  OAI22_X0P5M_A12TR u3045 ( .A0(n2823), .A1(n3639), .B0(n3598), .B1(n3584), 
        .Y(n3881) );
  INV_X0P5B_A12TR u3046 ( .A(n241), .Y(n3584) );
  NAND2_X0P5A_A12TR u3047 ( .A(n3088), .B(n35711), .Y(n3598) );
  INV_X0P5B_A12TR u3048 ( .A(alures[6]), .Y(n3639) );
  NAND2_X0P5A_A12TR u3049 ( .A(n3179), .B(n3070), .Y(n2929) );
  NOR2_X0P5A_A12TR u3050 ( .A(n30191), .B(n3036), .Y(n2928) );
  OAI211_X0P5M_A12TR u3051 ( .A0(n3409), .A1(n3900), .B0(n3901), .C0(n3902), 
        .Y(n2570) );
  AOI221_X0P5M_A12TR u3052 ( .A0(rdatahold2[0]), .A1(n2951), .B0(r194_sum_0_), 
        .B1(n2952), .C0(n3903), .Y(n3902) );
  MXIT2_X0P5M_A12TR u3053 ( .A(n3904), .B(n2943), .S0(pc[0]), .Y(n3903) );
  AOI22_X0P5M_A12TR u3054 ( .A0(r201_sum_0_), .A1(n2946), .B0(n2947), .B1(
        n3416), .Y(n3901) );
  INV_X0P5B_A12TR u3055 ( .A(n2950), .Y(n3900) );
  OAI211_X0P5M_A12TR u3056 ( .A0(n2943), .A1(n3905), .B0(n3906), .C0(n3907), 
        .Y(n2569) );
  AOI221_X0P5M_A12TR u3057 ( .A0(r201_sum_1_), .A1(n2946), .B0(r1226_sum_1_), 
        .B1(n2947), .C0(n3908), .Y(n3907) );
  AO22_X0P5M_A12TR u3058 ( .A0(n2949), .A1(n30100), .B0(n2950), .B1(n1151), 
        .Y(n3908) );
  AOI22_X0P5M_A12TR u3059 ( .A0(rdatahold2[1]), .A1(n2951), .B0(r194_sum_1_), 
        .B1(n2952), .Y(n3906) );
  OAI211_X0P5M_A12TR u3060 ( .A0(n2943), .A1(n3909), .B0(n3910), .C0(n3911), 
        .Y(n2568) );
  AOI221_X0P5M_A12TR u3061 ( .A0(r201_sum_2_), .A1(n2946), .B0(r1226_sum_2_), 
        .B1(n2947), .C0(n3912), .Y(n3911) );
  AO22_X0P5M_A12TR u3062 ( .A0(n2949), .A1(n30110), .B0(n2950), .B1(n1152), 
        .Y(n3912) );
  AOI22_X0P5M_A12TR u3063 ( .A0(rdatahold2[2]), .A1(n2951), .B0(r194_sum_2_), 
        .B1(n2952), .Y(n3910) );
  NAND4_X0P5A_A12TR u3064 ( .A(n3913), .B(n3914), .C(n3915), .D(n3916), .Y(
        n2567) );
  AOI32_X0P5M_A12TR u3065 ( .A0(n3917), .A1(n3918), .A2(r1226_sum_3_), .B0(
        n3919), .B1(n236), .Y(n3916) );
  AO21A1AI2_X0P5M_A12TR u3066 ( .A0(n3920), .A1(n3921), .B0(n3044), .C0(n3922), 
        .Y(n3918) );
  AOI22_X0P5M_A12TR u3067 ( .A0(r201_sum_3_), .A1(n2946), .B0(n1153), .B1(
        n2950), .Y(n3915) );
  AOI22_X0P5M_A12TR u3068 ( .A0(n30120), .A1(n2949), .B0(rdatahold2[3]), .B1(
        n2951), .Y(n3914) );
  AOI22_X0P5M_A12TR u3069 ( .A0(r194_sum_3_), .A1(n2952), .B0(pc[3]), .B1(
        n3923), .Y(n3913) );
  NAND4_X0P5A_A12TR u3070 ( .A(n3924), .B(n3925), .C(n3926), .D(n3927), .Y(
        n2566) );
  AOI32_X0P5M_A12TR u3071 ( .A0(n3917), .A1(n3928), .A2(r201_sum_4_), .B0(
        n3919), .B1(n46), .Y(n3927) );
  OAI31_X0P5M_A12TR u3072 ( .A0(n3044), .A1(n3288), .A2(n2831), .B0(n3379), 
        .Y(n3928) );
  AOI22_X0P5M_A12TR u3073 ( .A0(r1226_sum_4_), .A1(n2947), .B0(n1154), .B1(
        n2950), .Y(n3926) );
  AOI22_X0P5M_A12TR u3074 ( .A0(n30130), .A1(n2949), .B0(rdatahold2[4]), .B1(
        n2951), .Y(n3925) );
  AOI22_X0P5M_A12TR u3075 ( .A0(r194_sum_4_), .A1(n2952), .B0(pc[4]), .B1(
        n3923), .Y(n3924) );
  NAND4_X0P5A_A12TR u3076 ( .A(n3929), .B(n3930), .C(n3931), .D(n3932), .Y(
        n2565) );
  AOI22_X0P5M_A12TR u3077 ( .A0(n3933), .A1(r1226_sum_5_), .B0(n3919), .B1(
        n237), .Y(n3932) );
  NOR3_X0P5A_A12TR u3078 ( .A(n3934), .B(n3044), .C(n3192), .Y(n3919) );
  NAND2_X0P5A_A12TR u3079 ( .A(n235), .B(n234), .Y(n3192) );
  AOI21_X0P5M_A12TR u3080 ( .A0(n3922), .A1(n3935), .B0(n3934), .Y(n3933) );
  OAI31_X0P5M_A12TR u3081 ( .A0(n3936), .A1(n3560), .A2(n3937), .B0(n3112), 
        .Y(n3935) );
  INV_X0P5B_A12TR u3082 ( .A(n3938), .Y(n3937) );
  AOI22_X0P5M_A12TR u3083 ( .A0(r201_sum_5_), .A1(n2946), .B0(n1155), .B1(
        n2950), .Y(n3931) );
  AOI22_X0P5M_A12TR u3084 ( .A0(n30140), .A1(n2949), .B0(rdatahold2[5]), .B1(
        n2951), .Y(n3930) );
  AOI22_X0P5M_A12TR u3085 ( .A0(r194_sum_5_), .A1(n2952), .B0(pc[5]), .B1(
        n3923), .Y(n3929) );
  OAI211_X0P5M_A12TR u3086 ( .A0(n2943), .A1(n3939), .B0(n3940), .C0(n3941), 
        .Y(n2564) );
  AOI221_X0P5M_A12TR u3087 ( .A0(r201_sum_6_), .A1(n2946), .B0(r1226_sum_6_), 
        .B1(n2947), .C0(n3942), .Y(n3941) );
  AO22_X0P5M_A12TR u3088 ( .A0(n2949), .A1(n30150), .B0(n2950), .B1(n1156), 
        .Y(n3942) );
  AOI22_X0P5M_A12TR u3089 ( .A0(rdatahold2[6]), .A1(n2951), .B0(r194_sum_6_), 
        .B1(n2952), .Y(n3940) );
  OAI211_X0P5M_A12TR u3090 ( .A0(n3943), .A1(n2943), .B0(n3944), .C0(n3945), 
        .Y(n2563) );
  AOI221_X0P5M_A12TR u3091 ( .A0(n2946), .A1(r201_sum_7_), .B0(n2947), .B1(
        r1226_sum_7_), .C0(n3946), .Y(n3945) );
  AO22_X0P5M_A12TR u3092 ( .A0(n30160), .A1(n2949), .B0(n1157), .B1(n2950), 
        .Y(n3946) );
  AOI22_X0P5M_A12TR u3093 ( .A0(rdatahold2[7]), .A1(n2951), .B0(r194_sum_7_), 
        .B1(n2952), .Y(n3944) );
  OAI211_X0P5M_A12TR u3094 ( .A0(n3947), .A1(n2943), .B0(n3948), .C0(n3949), 
        .Y(n2562) );
  AOI221_X0P5M_A12TR u3095 ( .A0(r201_sum_8_), .A1(n2946), .B0(n2947), .B1(
        r1226_sum_8_), .C0(n3950), .Y(n3949) );
  AO22_X0P5M_A12TR u3096 ( .A0(n30170), .A1(n2949), .B0(n1158), .B1(n2950), 
        .Y(n3950) );
  AOI22_X0P5M_A12TR u3097 ( .A0(rdatahold[0]), .A1(n2951), .B0(r194_sum_8_), 
        .B1(n2952), .Y(n3948) );
  OAI211_X0P5M_A12TR u3098 ( .A0(n2834), .A1(n2943), .B0(n3951), .C0(n3952), 
        .Y(n2561) );
  AOI221_X0P5M_A12TR u3099 ( .A0(r201_sum_9_), .A1(n2946), .B0(r1226_sum_9_), 
        .B1(n2947), .C0(n3953), .Y(n3952) );
  AO22_X0P5M_A12TR u3100 ( .A0(n2949), .A1(n30180), .B0(n1159), .B1(n2950), 
        .Y(n3953) );
  AOI22_X0P5M_A12TR u3101 ( .A0(rdatahold[1]), .A1(n2951), .B0(r194_sum_9_), 
        .B1(n2952), .Y(n3951) );
  OAI211_X0P5M_A12TR u3102 ( .A0(n2852), .A1(n2943), .B0(n3954), .C0(n3955), 
        .Y(n2560) );
  AOI221_X0P5M_A12TR u3103 ( .A0(r201_sum_10_), .A1(n2946), .B0(r1226_sum_10_), 
        .B1(n2947), .C0(n3956), .Y(n3955) );
  AO22_X0P5M_A12TR u3104 ( .A0(n2949), .A1(n30190), .B0(n1160), .B1(n2950), 
        .Y(n3956) );
  AOI22_X0P5M_A12TR u3105 ( .A0(rdatahold[2]), .A1(n2951), .B0(r194_sum_10_), 
        .B1(n2952), .Y(n3954) );
  OAI211_X0P5M_A12TR u3106 ( .A0(n2849), .A1(n2943), .B0(n3957), .C0(n3958), 
        .Y(n2559) );
  AOI221_X0P5M_A12TR u3107 ( .A0(r201_sum_11_), .A1(n2946), .B0(r1226_sum_11_), 
        .B1(n2947), .C0(n3959), .Y(n3958) );
  AO22_X0P5M_A12TR u3108 ( .A0(n2949), .A1(n30200), .B0(n1161), .B1(n2950), 
        .Y(n3959) );
  AOI22_X0P5M_A12TR u3109 ( .A0(rdatahold[3]), .A1(n2951), .B0(r194_sum_11_), 
        .B1(n2952), .Y(n3957) );
  OAI211_X0P5M_A12TR u3110 ( .A0(n2846), .A1(n2943), .B0(n3960), .C0(n3961), 
        .Y(n2558) );
  AOI221_X0P5M_A12TR u3111 ( .A0(r201_sum_12_), .A1(n2946), .B0(r1226_sum_12_), 
        .B1(n2947), .C0(n3962), .Y(n3961) );
  AO22_X0P5M_A12TR u3112 ( .A0(n2949), .A1(n30210), .B0(n1162), .B1(n2950), 
        .Y(n3962) );
  AOI22_X0P5M_A12TR u3113 ( .A0(rdatahold[4]), .A1(n2951), .B0(r194_sum_12_), 
        .B1(n2952), .Y(n3960) );
  OAI211_X0P5M_A12TR u3114 ( .A0(n2843), .A1(n2943), .B0(n3963), .C0(n3964), 
        .Y(n2557) );
  AOI221_X0P5M_A12TR u3115 ( .A0(r201_sum_13_), .A1(n2946), .B0(r1226_sum_13_), 
        .B1(n2947), .C0(n3965), .Y(n3964) );
  AO22_X0P5M_A12TR u3116 ( .A0(n2949), .A1(n30220), .B0(n1163), .B1(n2950), 
        .Y(n3965) );
  AOI22_X0P5M_A12TR u3117 ( .A0(rdatahold[5]), .A1(n2951), .B0(r194_sum_13_), 
        .B1(n2952), .Y(n3963) );
  OAI211_X0P5M_A12TR u3118 ( .A0(n2840), .A1(n2943), .B0(n3966), .C0(n3967), 
        .Y(n2556) );
  AOI221_X0P5M_A12TR u3119 ( .A0(r201_sum_14_), .A1(n2946), .B0(r1226_sum_14_), 
        .B1(n2947), .C0(n3968), .Y(n3967) );
  AO22_X0P5M_A12TR u3120 ( .A0(n2949), .A1(n30230), .B0(n1164), .B1(n2950), 
        .Y(n3968) );
  NOR3_X0P5A_A12TR u3121 ( .A(n3044), .B(n3969), .C(n3934), .Y(n2950) );
  INV_X0P5B_A12TR u3122 ( .A(n3904), .Y(n2949) );
  NAND2_X0P5A_A12TR u3123 ( .A(n3031), .B(n3917), .Y(n3904) );
  AOI21_X0P5M_A12TR u3124 ( .A0(n3384), .A1(n3191), .B0(n3193), .Y(n3031) );
  NOR2B_X0P5M_A12TR u3125 ( .AN(n3970), .B(n3934), .Y(n2947) );
  AO21A1AI2_X0P5M_A12TR u3126 ( .A0(n3920), .A1(n3938), .B0(n3044), .C0(n3922), 
        .Y(n3970) );
  INV_X0P5B_A12TR u3127 ( .A(n3971), .Y(n3922) );
  NAND4B_X0P5M_A12TR u3128 ( .AN(n3972), .B(n3392), .C(n3773), .D(n3973), .Y(
        n3971) );
  OAI21_X0P5M_A12TR u3129 ( .A0(n3974), .A1(n3975), .B0(n3127), .Y(n3973) );
  NAND2_X0P5A_A12TR u3130 ( .A(n3127), .B(n3771), .Y(n3773) );
  NAND2_X0P5A_A12TR u3131 ( .A(n3040), .B(n3366), .Y(n3392) );
  NAND2_X0P5A_A12TR u3132 ( .A(n2920), .B(n3128), .Y(n3938) );
  AOI21_X0P5M_A12TR u3133 ( .A0(n3128), .A1(n3560), .B0(n3936), .Y(n3920) );
  AO21A1AI2_X0P5M_A12TR u3134 ( .A0(n236), .A1(n3289), .B0(n234), .C0(n3343), 
        .Y(n3936) );
  NOR2_X0P5A_A12TR u3135 ( .A(n3290), .B(n3288), .Y(n3560) );
  AOI21_X0P5M_A12TR u3136 ( .A0(n3379), .A1(n3976), .B0(n3934), .Y(n2946) );
  NAND4_X0P5A_A12TR u3137 ( .A(n3112), .B(n3204), .C(n234), .D(n3128), .Y(
        n3976) );
  INV_X0P5B_A12TR u3138 ( .A(n3044), .Y(n3112) );
  NAND2_X0P5A_A12TR u3139 ( .A(n3366), .B(n233), .Y(n3044) );
  NOR2_X0P5A_A12TR u3140 ( .A(n3977), .B(n3978), .Y(n3379) );
  AOI22_X0P5M_A12TR u3141 ( .A0(rdatahold[6]), .A1(n2951), .B0(r194_sum_14_), 
        .B1(n2952), .Y(n3966) );
  AND3_X0P5M_A12TR u3142 ( .A(n3127), .B(n2858), .C(n3917), .Y(n2952) );
  INV_X0P5B_A12TR u3143 ( .A(n3934), .Y(n3917) );
  NAND4_X0P5A_A12TR u3144 ( .A(n2943), .B(n3181), .C(n3153), .D(n30111), .Y(
        n3934) );
  AOI211_X0P5M_A12TR u3145 ( .A0(n3730), .A1(n30111), .B0(n3923), .C0(reset), 
        .Y(n2951) );
  INV_X0P5B_A12TR u3146 ( .A(n2943), .Y(n3923) );
  OAI211_X0P5M_A12TR u3147 ( .A0(n30141), .A1(n30211), .B0(n3221), .C0(n3979), 
        .Y(n2943) );
  AOI222_X0P5M_A12TR u3148 ( .A0(n3320), .A1(n3980), .B0(n3855), .B1(n3972), 
        .C0(n3076), .C1(n3981), .Y(n3979) );
  NAND2_X0P5A_A12TR u3149 ( .A(n3111), .B(n3228), .Y(n3972) );
  NAND4B_X0P5M_A12TR u3150 ( .AN(n3771), .B(n3404), .C(n3982), .D(n3983), .Y(
        n3980) );
  AND3_X0P5M_A12TR u3151 ( .A(n3969), .B(n3123), .C(n3191), .Y(n3983) );
  NOR2_X0P5A_A12TR u3152 ( .A(n3984), .B(n2825), .Y(n3404) );
  INV_X0P5B_A12TR u3153 ( .A(n3329), .Y(n3320) );
  INV_X0P5B_A12TR u3154 ( .A(n3985), .Y(n3221) );
  AO21A1AI2_X0P5M_A12TR u3155 ( .A0(n3986), .A1(n3987), .B0(n3405), .C0(n3181), 
        .Y(n3985) );
  NOR3_X0P5A_A12TR u3156 ( .A(n2967), .B(n3114), .C(n3974), .Y(n3987) );
  NAND3B_X0P5M_A12TR u3157 ( .AN(n3899), .B(n3375), .C(n2977), .Y(n3974) );
  INV_X0P5B_A12TR u3158 ( .A(n2924), .Y(n2977) );
  NAND4_X0P5A_A12TR u3159 ( .A(n3311), .B(n3988), .C(n3989), .D(n3641), .Y(
        n3114) );
  AND2_X0P5M_A12TR u3160 ( .A(n3490), .B(n3395), .Y(n3989) );
  OAI21_X0P5M_A12TR u3161 ( .A0(n3990), .A1(n2984), .B0(n3125), .Y(n3490) );
  AOI21_X0P5M_A12TR u3162 ( .A0(n3290), .A1(n3991), .B0(n3372), .Y(n3311) );
  NAND3_X0P5A_A12TR u3163 ( .A(n3992), .B(n3123), .C(n3343), .Y(n3372) );
  INV_X0P5B_A12TR u3164 ( .A(n3993), .Y(n2967) );
  NOR2_X0P5A_A12TR u3165 ( .A(n3994), .B(n3771), .Y(n3986) );
  NAND3_X0P5A_A12TR u3166 ( .A(state[2]), .B(n2859), .C(state[0]), .Y(n30211)
         );
  OAI211_X0P5M_A12TR u3167 ( .A0(n3995), .A1(n3996), .B0(n3997), .C0(n3998), 
        .Y(n2555) );
  AOI222_X0P5M_A12TR u3168 ( .A0(sp[15]), .A1(n3999), .B0(n4000), .B1(n1165), 
        .C0(n31520), .C1(n4001), .Y(n3998) );
  AOI22_X0P5M_A12TR u3169 ( .A0(n4002), .A1(rdatahold[7]), .B0(r194_sum_15_), 
        .B1(n4003), .Y(n3997) );
  INV_X0P5B_A12TR u3170 ( .A(n26720), .Y(n3996) );
  OAI211_X0P5M_A12TR u3171 ( .A0(n2975), .A1(n4004), .B0(n4005), .C0(n4006), 
        .Y(n2554) );
  AOI22_X0P5M_A12TR u3172 ( .A0(r194_sum_0_), .A1(n4003), .B0(n4000), .B1(
        n1150), .Y(n4006) );
  OAI31_X0P5M_A12TR u3173 ( .A0(n3999), .A1(n4007), .A2(n4001), .B0(n31370), 
        .Y(n4005) );
  INV_X0P5B_A12TR u3174 ( .A(n4002), .Y(n4004) );
  INV_X0P5B_A12TR u3175 ( .A(rdatahold2[0]), .Y(n2975) );
  OAI211_X0P5M_A12TR u3176 ( .A0(n3420), .A1(n4008), .B0(n4009), .C0(n4010), 
        .Y(n2553) );
  AOI222_X0P5M_A12TR u3177 ( .A0(n26580), .A1(n4007), .B0(n4002), .B1(
        rdatahold2[1]), .C0(r194_sum_1_), .C1(n4003), .Y(n4010) );
  MXIT2_X0P5M_A12TR u3178 ( .A(n4001), .B(n3999), .S0(sp[1]), .Y(n4009) );
  INV_X0P5B_A12TR u3179 ( .A(n4000), .Y(n4008) );
  OAI211_X0P5M_A12TR u3180 ( .A0(n3995), .A1(n4011), .B0(n4012), .C0(n4013), 
        .Y(n2552) );
  AOI222_X0P5M_A12TR u3181 ( .A0(sp[2]), .A1(n3999), .B0(n4000), .B1(n1152), 
        .C0(n31390), .C1(n4001), .Y(n4013) );
  AOI22_X0P5M_A12TR u3182 ( .A0(n4002), .A1(rdatahold2[2]), .B0(r194_sum_2_), 
        .B1(n4003), .Y(n4012) );
  INV_X0P5B_A12TR u3183 ( .A(n26590), .Y(n4011) );
  OAI211_X0P5M_A12TR u3184 ( .A0(n3995), .A1(n4014), .B0(n4015), .C0(n4016), 
        .Y(n2551) );
  AOI222_X0P5M_A12TR u3185 ( .A0(sp[3]), .A1(n3999), .B0(n4000), .B1(n1153), 
        .C0(n31400), .C1(n4001), .Y(n4016) );
  AOI22_X0P5M_A12TR u3186 ( .A0(n4002), .A1(rdatahold2[3]), .B0(r194_sum_3_), 
        .B1(n4003), .Y(n4015) );
  INV_X0P5B_A12TR u3187 ( .A(n26600), .Y(n4014) );
  OAI211_X0P5M_A12TR u3188 ( .A0(n3995), .A1(n4017), .B0(n4018), .C0(n4019), 
        .Y(n2550) );
  AOI222_X0P5M_A12TR u3189 ( .A0(sp[4]), .A1(n3999), .B0(n4000), .B1(n1154), 
        .C0(n31410), .C1(n4001), .Y(n4019) );
  AOI22_X0P5M_A12TR u3190 ( .A0(n4002), .A1(rdatahold2[4]), .B0(r194_sum_4_), 
        .B1(n4003), .Y(n4018) );
  INV_X0P5B_A12TR u3191 ( .A(n26610), .Y(n4017) );
  OAI211_X0P5M_A12TR u3192 ( .A0(n3995), .A1(n4020), .B0(n4021), .C0(n4022), 
        .Y(n2549) );
  AOI222_X0P5M_A12TR u3193 ( .A0(sp[5]), .A1(n3999), .B0(n4000), .B1(n1155), 
        .C0(n31420), .C1(n4001), .Y(n4022) );
  AOI22_X0P5M_A12TR u3194 ( .A0(n4002), .A1(rdatahold2[5]), .B0(r194_sum_5_), 
        .B1(n4003), .Y(n4021) );
  INV_X0P5B_A12TR u3195 ( .A(n26620), .Y(n4020) );
  OAI211_X0P5M_A12TR u3196 ( .A0(n3995), .A1(n4023), .B0(n4024), .C0(n4025), 
        .Y(n2548) );
  AOI222_X0P5M_A12TR u3197 ( .A0(sp[6]), .A1(n3999), .B0(n4000), .B1(n1156), 
        .C0(n31430), .C1(n4001), .Y(n4025) );
  AOI22_X0P5M_A12TR u3198 ( .A0(n4002), .A1(rdatahold2[6]), .B0(r194_sum_6_), 
        .B1(n4003), .Y(n4024) );
  INV_X0P5B_A12TR u3199 ( .A(n26630), .Y(n4023) );
  OAI211_X0P5M_A12TR u3200 ( .A0(n3995), .A1(n4026), .B0(n4027), .C0(n4028), 
        .Y(n2547) );
  AOI222_X0P5M_A12TR u3201 ( .A0(sp[7]), .A1(n3999), .B0(n4000), .B1(n1157), 
        .C0(n31440), .C1(n4001), .Y(n4028) );
  AOI22_X0P5M_A12TR u3202 ( .A0(n4002), .A1(rdatahold2[7]), .B0(r194_sum_7_), 
        .B1(n4003), .Y(n4027) );
  INV_X0P5B_A12TR u3203 ( .A(n26640), .Y(n4026) );
  OAI211_X0P5M_A12TR u3204 ( .A0(n3995), .A1(n4029), .B0(n4030), .C0(n4031), 
        .Y(n2546) );
  AOI222_X0P5M_A12TR u3205 ( .A0(sp[8]), .A1(n3999), .B0(n4000), .B1(n1158), 
        .C0(n31450), .C1(n4001), .Y(n4031) );
  AOI22_X0P5M_A12TR u3206 ( .A0(n4002), .A1(rdatahold[0]), .B0(r194_sum_8_), 
        .B1(n4003), .Y(n4030) );
  INV_X0P5B_A12TR u3207 ( .A(n26650), .Y(n4029) );
  OAI211_X0P5M_A12TR u3208 ( .A0(n3995), .A1(n4032), .B0(n4033), .C0(n4034), 
        .Y(n2545) );
  AOI222_X0P5M_A12TR u3209 ( .A0(sp[9]), .A1(n3999), .B0(n4000), .B1(n1159), 
        .C0(n31460), .C1(n4001), .Y(n4034) );
  AOI22_X0P5M_A12TR u3210 ( .A0(n4002), .A1(rdatahold[1]), .B0(r194_sum_9_), 
        .B1(n4003), .Y(n4033) );
  INV_X0P5B_A12TR u3211 ( .A(n26660), .Y(n4032) );
  OAI211_X0P5M_A12TR u3212 ( .A0(n3995), .A1(n4035), .B0(n4036), .C0(n4037), 
        .Y(n2544) );
  AOI222_X0P5M_A12TR u3213 ( .A0(sp[10]), .A1(n3999), .B0(n4000), .B1(n1160), 
        .C0(n31470), .C1(n4001), .Y(n4037) );
  AOI22_X0P5M_A12TR u3214 ( .A0(n4002), .A1(rdatahold[2]), .B0(r194_sum_10_), 
        .B1(n4003), .Y(n4036) );
  INV_X0P5B_A12TR u3215 ( .A(n26670), .Y(n4035) );
  OAI211_X0P5M_A12TR u3216 ( .A0(n3995), .A1(n4038), .B0(n4039), .C0(n4040), 
        .Y(n2543) );
  AOI222_X0P5M_A12TR u3217 ( .A0(sp[11]), .A1(n3999), .B0(n4000), .B1(n1161), 
        .C0(n31480), .C1(n4001), .Y(n4040) );
  AOI22_X0P5M_A12TR u3218 ( .A0(n4002), .A1(rdatahold[3]), .B0(r194_sum_11_), 
        .B1(n4003), .Y(n4039) );
  INV_X0P5B_A12TR u3219 ( .A(n26680), .Y(n4038) );
  OAI211_X0P5M_A12TR u3220 ( .A0(n3995), .A1(n4041), .B0(n4042), .C0(n4043), 
        .Y(n2542) );
  AOI222_X0P5M_A12TR u3221 ( .A0(sp[12]), .A1(n3999), .B0(n4000), .B1(n1162), 
        .C0(n31490), .C1(n4001), .Y(n4043) );
  AOI22_X0P5M_A12TR u3222 ( .A0(n4002), .A1(rdatahold[4]), .B0(r194_sum_12_), 
        .B1(n4003), .Y(n4042) );
  INV_X0P5B_A12TR u3223 ( .A(n26690), .Y(n4041) );
  OAI211_X0P5M_A12TR u3224 ( .A0(n3995), .A1(n4044), .B0(n4045), .C0(n4046), 
        .Y(n2541) );
  AOI222_X0P5M_A12TR u3225 ( .A0(sp[13]), .A1(n3999), .B0(n4000), .B1(n1163), 
        .C0(n31500), .C1(n4001), .Y(n4046) );
  AOI22_X0P5M_A12TR u3226 ( .A0(n4002), .A1(rdatahold[5]), .B0(r194_sum_13_), 
        .B1(n4003), .Y(n4045) );
  INV_X0P5B_A12TR u3227 ( .A(n26700), .Y(n4044) );
  OAI211_X0P5M_A12TR u3228 ( .A0(n3995), .A1(n4047), .B0(n4048), .C0(n4049), 
        .Y(n2540) );
  AOI222_X0P5M_A12TR u3229 ( .A0(sp[14]), .A1(n3999), .B0(n4000), .B1(n1164), 
        .C0(n31510), .C1(n4001), .Y(n4049) );
  NOR2_X0P5A_A12TR u3230 ( .A(n4050), .B(n3426), .Y(n4001) );
  NOR2_X0P5A_A12TR u3231 ( .A(n4051), .B(n4050), .Y(n4000) );
  AOI22_X0P5M_A12TR u3232 ( .A0(n4002), .A1(rdatahold[6]), .B0(r194_sum_14_), 
        .B1(n4003), .Y(n4048) );
  OAI22_X0P5M_A12TR u3233 ( .A0(n30111), .A1(n3999), .B0(n3036), .B1(n4050), 
        .Y(n4003) );
  NOR2_X0P5A_A12TR u3234 ( .A(n3999), .B(n3153), .Y(n4002) );
  INV_X0P5B_A12TR u3235 ( .A(n26710), .Y(n4047) );
  INV_X0P5B_A12TR u3236 ( .A(n4007), .Y(n3995) );
  NOR2_X0P5A_A12TR u3237 ( .A(n4050), .B(n3374), .Y(n4007) );
  NAND2B_X0P5M_A12TR u3238 ( .AN(n3999), .B(n2859), .Y(n4050) );
  NAND2_X0P5A_A12TR u3239 ( .A(n3181), .B(n4052), .Y(n3999) );
  OAI211_X0P5M_A12TR u3240 ( .A0(n2861), .A1(n3405), .B0(n4053), .C0(n4054), 
        .Y(n4052) );
  AOI22_X0P5M_A12TR u3241 ( .A0(n3076), .A1(n3981), .B0(n4055), .B1(n3855), 
        .Y(n4054) );
  OAI22_X0P5M_A12TR u3242 ( .A0(n3004), .A1(n3231), .B0(u3_u93_z_6), .B1(
        n30191), .Y(n3981) );
  INV_X0P5B_A12TR u3243 ( .A(n3069), .Y(n3076) );
  AOI31_X0P5M_A12TR u3244 ( .A0(n2894), .A1(state[0]), .A2(n3246), .B0(n4056), 
        .Y(n4053) );
  AOI21_X0P5M_A12TR u3245 ( .A0(n3374), .A1(n4051), .B0(n3329), .Y(n4056) );
  NAND2_X0P5A_A12TR u3246 ( .A(n3855), .B(n3366), .Y(n3329) );
  NOR2_X0P5A_A12TR u3247 ( .A(n3984), .B(n3365), .Y(n3374) );
  INV_X0P5B_A12TR u3248 ( .A(n3316), .Y(n3365) );
  INV_X0P5B_A12TR u3249 ( .A(n30141), .Y(n2894) );
  NAND2_X0P5A_A12TR u3250 ( .A(n3855), .B(n3127), .Y(n3405) );
  OAI211_X0P5M_A12TR u3251 ( .A0(n2482), .A1(n4057), .B0(n4058), .C0(n4059), 
        .Y(n2539) );
  OA211_X0P5M_A12TR u3252 ( .A0(n4060), .A1(n3858), .B0(n4061), .C0(n4062), 
        .Y(n4059) );
  OAI31_X0P5M_A12TR u3253 ( .A0(n4063), .A1(n4064), .A2(n4065), .B0(n31370), 
        .Y(n4062) );
  AOI22_X0P5M_A12TR u3254 ( .A0(n3416), .A1(n4066), .B0(n1657), .B1(n4067), 
        .Y(n4061) );
  INV_X0P5B_A12TR u3255 ( .A(u3_u84_z_0), .Y(n3416) );
  AOI22_X0P5M_A12TR u3256 ( .A0(n1150), .A1(n4068), .B0(n4069), .B1(
        rdatahold2[0]), .Y(n4058) );
  NAND4_X0P5A_A12TR u3257 ( .A(n4070), .B(n4071), .C(n4072), .D(n4073), .Y(
        n2538) );
  AOI22_X0P5M_A12TR u3258 ( .A0(n4065), .A1(n26580), .B0(n4074), .B1(n1168), 
        .Y(n4073) );
  AOI22_X0P5M_A12TR u3259 ( .A0(n4067), .A1(n1658), .B0(n4066), .B1(
        r1226_sum_1_), .Y(n4072) );
  AOI22_X0P5M_A12TR u3260 ( .A0(n1151), .A1(n4068), .B0(n4069), .B1(
        rdatahold2[1]), .Y(n4071) );
  AOI21_X0P5M_A12TR u3261 ( .A0(n4075), .A1(n4076), .B0(n4077), .Y(n4070) );
  MXT2_X0P5M_A12TR u3262 ( .A(n4064), .B(n4063), .S0(n4078), .Y(n4077) );
  NAND4_X0P5A_A12TR u3263 ( .A(n4079), .B(n4080), .C(n4081), .D(n4082), .Y(
        n2537) );
  AOI222_X0P5M_A12TR u3264 ( .A0(n4067), .A1(n1659), .B0(n4065), .B1(n26590), 
        .C0(n4074), .C1(n1169), .Y(n4082) );
  AOI22_X0P5M_A12TR u3265 ( .A0(n4063), .A1(n31390), .B0(n4064), .B1(sp[2]), 
        .Y(n4081) );
  AOI22_X0P5M_A12TR u3266 ( .A0(n4066), .A1(r1226_sum_2_), .B0(n1152), .B1(
        n4068), .Y(n4080) );
  AOI22_X0P5M_A12TR u3267 ( .A0(n4069), .A1(rdatahold2[2]), .B0(n4075), .B1(
        n4083), .Y(n4079) );
  NAND4_X0P5A_A12TR u3268 ( .A(n4084), .B(n4085), .C(n4086), .D(n4087), .Y(
        n2536) );
  AOI222_X0P5M_A12TR u3269 ( .A0(n4067), .A1(n1660), .B0(n4065), .B1(n26600), 
        .C0(n4074), .C1(n1170), .Y(n4087) );
  AOI22_X0P5M_A12TR u3270 ( .A0(n4063), .A1(n31400), .B0(n4064), .B1(sp[3]), 
        .Y(n4086) );
  AOI22_X0P5M_A12TR u3271 ( .A0(n4066), .A1(r1226_sum_3_), .B0(n1153), .B1(
        n4068), .Y(n4085) );
  AOI22_X0P5M_A12TR u3272 ( .A0(n4069), .A1(rdatahold2[3]), .B0(n4075), .B1(
        n4088), .Y(n4084) );
  NAND4_X0P5A_A12TR u3273 ( .A(n4089), .B(n4090), .C(n4091), .D(n4092), .Y(
        n2535) );
  AOI222_X0P5M_A12TR u3274 ( .A0(n4067), .A1(n1661), .B0(n4065), .B1(n26610), 
        .C0(n4074), .C1(n1171), .Y(n4092) );
  AOI22_X0P5M_A12TR u3275 ( .A0(n4063), .A1(n31410), .B0(n4064), .B1(sp[4]), 
        .Y(n4091) );
  AOI22_X0P5M_A12TR u3276 ( .A0(n4066), .A1(r1226_sum_4_), .B0(n1154), .B1(
        n4068), .Y(n4090) );
  AOI22_X0P5M_A12TR u3277 ( .A0(n4069), .A1(rdatahold2[4]), .B0(n4075), .B1(
        n4093), .Y(n4089) );
  NAND4_X0P5A_A12TR u3278 ( .A(n4094), .B(n4095), .C(n4096), .D(n4097), .Y(
        n2534) );
  AOI222_X0P5M_A12TR u3279 ( .A0(n4067), .A1(n1662), .B0(n4065), .B1(n26620), 
        .C0(n4074), .C1(n1172), .Y(n4097) );
  AOI22_X0P5M_A12TR u3280 ( .A0(n4063), .A1(n31420), .B0(n4064), .B1(sp[5]), 
        .Y(n4096) );
  AOI22_X0P5M_A12TR u3281 ( .A0(n4066), .A1(r1226_sum_5_), .B0(n1155), .B1(
        n4068), .Y(n4095) );
  AOI22_X0P5M_A12TR u3282 ( .A0(n4069), .A1(rdatahold2[5]), .B0(n4075), .B1(
        n4098), .Y(n4094) );
  NAND4_X0P5A_A12TR u3283 ( .A(n4099), .B(n4100), .C(n4101), .D(n4102), .Y(
        n2533) );
  AOI222_X0P5M_A12TR u3284 ( .A0(n4067), .A1(n1663), .B0(n4065), .B1(n26630), 
        .C0(n4074), .C1(n1173), .Y(n4102) );
  AOI22_X0P5M_A12TR u3285 ( .A0(n4063), .A1(n31430), .B0(n4064), .B1(sp[6]), 
        .Y(n4101) );
  AOI22_X0P5M_A12TR u3286 ( .A0(n4066), .A1(r1226_sum_6_), .B0(n1156), .B1(
        n4068), .Y(n4100) );
  AOI22_X0P5M_A12TR u3287 ( .A0(n4069), .A1(rdatahold2[6]), .B0(n4075), .B1(
        n4103), .Y(n4099) );
  NAND4_X0P5A_A12TR u3288 ( .A(n4104), .B(n4105), .C(n4106), .D(n4107), .Y(
        n2532) );
  AOI222_X0P5M_A12TR u3289 ( .A0(n4067), .A1(n1664), .B0(n4065), .B1(n26640), 
        .C0(n4074), .C1(n1174), .Y(n4107) );
  AOI22_X0P5M_A12TR u3290 ( .A0(n4063), .A1(n31440), .B0(n4064), .B1(sp[7]), 
        .Y(n4106) );
  AOI22_X0P5M_A12TR u3291 ( .A0(n4066), .A1(r1226_sum_7_), .B0(n1157), .B1(
        n4068), .Y(n4105) );
  AOI22_X0P5M_A12TR u3292 ( .A0(n4069), .A1(rdatahold2[7]), .B0(n4075), .B1(
        n4108), .Y(n4104) );
  NAND4_X0P5A_A12TR u3293 ( .A(n4109), .B(n4110), .C(n4111), .D(n4112), .Y(
        n2531) );
  AOI222_X0P5M_A12TR u3294 ( .A0(n4067), .A1(regfil_2__0_), .B0(n4065), .B1(
        n26650), .C0(n4074), .C1(n1175), .Y(n4112) );
  AOI22_X0P5M_A12TR u3295 ( .A0(n4063), .A1(n31450), .B0(n4064), .B1(sp[8]), 
        .Y(n4111) );
  AOI22_X0P5M_A12TR u3296 ( .A0(n4066), .A1(r1226_sum_8_), .B0(n1158), .B1(
        n4068), .Y(n4110) );
  AOI22_X0P5M_A12TR u3297 ( .A0(n4069), .A1(rdatahold[0]), .B0(n4075), .B1(
        n4113), .Y(n4109) );
  NAND4_X0P5A_A12TR u3298 ( .A(n4114), .B(n4115), .C(n4116), .D(n4117), .Y(
        n2530) );
  AOI222_X0P5M_A12TR u3299 ( .A0(n4067), .A1(regfil_2__1_), .B0(n4065), .B1(
        n26660), .C0(n4074), .C1(n1176), .Y(n4117) );
  AOI22_X0P5M_A12TR u3300 ( .A0(n4063), .A1(n31460), .B0(n4064), .B1(sp[9]), 
        .Y(n4116) );
  AOI22_X0P5M_A12TR u3301 ( .A0(n4066), .A1(r1226_sum_9_), .B0(n1159), .B1(
        n4068), .Y(n4115) );
  AOI22_X0P5M_A12TR u3302 ( .A0(n4069), .A1(rdatahold[1]), .B0(n4075), .B1(
        n4118), .Y(n4114) );
  NAND4_X0P5A_A12TR u3303 ( .A(n4119), .B(n4120), .C(n4121), .D(n4122), .Y(
        n2529) );
  AOI222_X0P5M_A12TR u3304 ( .A0(n4067), .A1(regfil_2__2_), .B0(n4065), .B1(
        n26670), .C0(n4074), .C1(n1177), .Y(n4122) );
  AOI22_X0P5M_A12TR u3305 ( .A0(n4063), .A1(n31470), .B0(n4064), .B1(sp[10]), 
        .Y(n4121) );
  AOI22_X0P5M_A12TR u3306 ( .A0(n4066), .A1(r1226_sum_10_), .B0(n1160), .B1(
        n4068), .Y(n4120) );
  AOI22_X0P5M_A12TR u3307 ( .A0(n4069), .A1(rdatahold[2]), .B0(n4075), .B1(
        n4123), .Y(n4119) );
  NAND4_X0P5A_A12TR u3308 ( .A(n4124), .B(n4125), .C(n4126), .D(n4127), .Y(
        n2528) );
  AOI222_X0P5M_A12TR u3309 ( .A0(n4067), .A1(regfil_2__3_), .B0(n4065), .B1(
        n26680), .C0(n4074), .C1(n1178), .Y(n4127) );
  AOI22_X0P5M_A12TR u3310 ( .A0(n4063), .A1(n31480), .B0(n4064), .B1(sp[11]), 
        .Y(n4126) );
  AOI22_X0P5M_A12TR u3311 ( .A0(n4066), .A1(r1226_sum_11_), .B0(n1161), .B1(
        n4068), .Y(n4125) );
  AOI22_X0P5M_A12TR u3312 ( .A0(n4069), .A1(rdatahold[3]), .B0(n4075), .B1(
        n4128), .Y(n4124) );
  NAND4_X0P5A_A12TR u3313 ( .A(n4129), .B(n4130), .C(n4131), .D(n4132), .Y(
        n2527) );
  AOI222_X0P5M_A12TR u3314 ( .A0(n4067), .A1(regfil_2__4_), .B0(n4065), .B1(
        n26690), .C0(n4074), .C1(n1179), .Y(n4132) );
  AOI22_X0P5M_A12TR u3315 ( .A0(n4063), .A1(n31490), .B0(n4064), .B1(sp[12]), 
        .Y(n4131) );
  AOI22_X0P5M_A12TR u3316 ( .A0(n4066), .A1(r1226_sum_12_), .B0(n1162), .B1(
        n4068), .Y(n4130) );
  AOI22_X0P5M_A12TR u3317 ( .A0(n4069), .A1(rdatahold[4]), .B0(n4075), .B1(
        n4133), .Y(n4129) );
  NAND4_X0P5A_A12TR u3318 ( .A(n4134), .B(n4135), .C(n4136), .D(n4137), .Y(
        n2526) );
  AOI222_X0P5M_A12TR u3319 ( .A0(n4067), .A1(regfil_2__5_), .B0(n4065), .B1(
        n26700), .C0(n4074), .C1(n1180), .Y(n4137) );
  AOI22_X0P5M_A12TR u3320 ( .A0(n4063), .A1(n31500), .B0(n4064), .B1(sp[13]), 
        .Y(n4136) );
  AOI22_X0P5M_A12TR u3321 ( .A0(n4066), .A1(r1226_sum_13_), .B0(n1163), .B1(
        n4068), .Y(n4135) );
  AOI22_X0P5M_A12TR u3322 ( .A0(n4069), .A1(rdatahold[5]), .B0(n4075), .B1(
        n4138), .Y(n4134) );
  NAND4_X0P5A_A12TR u3323 ( .A(n4139), .B(n4140), .C(n4141), .D(n4142), .Y(
        n2525) );
  AOI222_X0P5M_A12TR u3324 ( .A0(n4067), .A1(regfil_2__6_), .B0(n4065), .B1(
        n26710), .C0(n4074), .C1(n1181), .Y(n4142) );
  AOI22_X0P5M_A12TR u3325 ( .A0(n4063), .A1(n31510), .B0(n4064), .B1(sp[14]), 
        .Y(n4141) );
  AOI22_X0P5M_A12TR u3326 ( .A0(n4066), .A1(r1226_sum_14_), .B0(n1164), .B1(
        n4068), .Y(n4140) );
  AOI22_X0P5M_A12TR u3327 ( .A0(n4069), .A1(rdatahold[6]), .B0(n4075), .B1(
        n4143), .Y(n4139) );
  NAND4_X0P5A_A12TR u3328 ( .A(n4144), .B(n4145), .C(n4146), .D(n4147), .Y(
        n2524) );
  AOI222_X0P5M_A12TR u3329 ( .A0(n4067), .A1(regfil_2__7_), .B0(n4065), .B1(
        n26720), .C0(n4074), .C1(n1182), .Y(n4147) );
  INV_X0P5B_A12TR u3330 ( .A(n4060), .Y(n4074) );
  NAND3_X0P5A_A12TR u3331 ( .A(n4148), .B(n3289), .C(n3164), .Y(n4060) );
  NOR3_X0P5A_A12TR u3332 ( .A(n3193), .B(n4307), .C(n4149), .Y(n4065) );
  AND3_X0P5M_A12TR u3333 ( .A(n4148), .B(n46), .C(n3164), .Y(n4067) );
  AOI22_X0P5M_A12TR u3334 ( .A0(n4063), .A1(n31520), .B0(n4064), .B1(sp[15]), 
        .Y(n4146) );
  AND2_X0P5M_A12TR u3335 ( .A(n3351), .B(n4148), .Y(n4064) );
  INV_X0P5B_A12TR u3336 ( .A(n4149), .Y(n4148) );
  NOR2_X0P5A_A12TR u3337 ( .A(n4149), .B(n3357), .Y(n4063) );
  AOI22_X0P5M_A12TR u3338 ( .A0(n4066), .A1(r1226_sum_15_), .B0(n1165), .B1(
        n4068), .Y(n4145) );
  OAI22_X0P5M_A12TR u3339 ( .A0(n4075), .A1(n30111), .B0(n4150), .B1(n4149), 
        .Y(n4068) );
  NAND2_X0P5A_A12TR u3340 ( .A(n4057), .B(n2823), .Y(n4149) );
  NOR2_X0P5A_A12TR u3341 ( .A(n3978), .B(n35711), .Y(n4150) );
  NOR2_X0P5A_A12TR u3342 ( .A(n3646), .B(n4075), .Y(n4066) );
  AOI22_X0P5M_A12TR u3343 ( .A0(n4069), .A1(rdatahold[7]), .B0(n4075), .B1(
        n4151), .Y(n4144) );
  NOR2_X0P5A_A12TR u3344 ( .A(n3179), .B(n4075), .Y(n4069) );
  INV_X0P5B_A12TR u3345 ( .A(n4057), .Y(n4075) );
  OAI221_X0P5M_A12TR u3346 ( .A0(n3492), .A1(n4152), .B0(n4153), .B1(n3298), 
        .C0(n4154), .Y(n4057) );
  INV_X0P5B_A12TR u3347 ( .A(n3396), .Y(n4154) );
  NOR2_X0P5A_A12TR u3348 ( .A(n3110), .B(n3298), .Y(n3396) );
  NAND3_X0P5A_A12TR u3349 ( .A(n2984), .B(n3027), .C(n35711), .Y(n3110) );
  NAND3_X0P5A_A12TR u3350 ( .A(n2984), .B(n3570), .C(n35711), .Y(n3027) );
  AOI211_X0P5M_A12TR u3351 ( .A0(n3978), .A1(n2984), .B0(n4155), .C0(n3164), 
        .Y(n4153) );
  AND3_X0P5M_A12TR u3352 ( .A(n3990), .B(n3127), .C(n3125), .Y(n3164) );
  INV_X0P5B_A12TR u3353 ( .A(n4156), .Y(n4155) );
  NOR2_X0P5A_A12TR u3354 ( .A(n3123), .B(n3036), .Y(n3978) );
  INV_X0P5B_A12TR u3355 ( .A(n3570), .Y(n3123) );
  MXIT2_X0P5M_A12TR u3356 ( .A(n3239), .B(n3072), .S0(state[0]), .Y(n4152) );
  OAI21_X0P5M_A12TR u3357 ( .A0(state[5]), .A1(n30171), .B0(n3069), .Y(n3072)
         );
  NAND2_X0P5A_A12TR u3358 ( .A(state[5]), .B(n30131), .Y(n3069) );
  NOR2_X0P5A_A12TR u3359 ( .A(n30141), .B(state[5]), .Y(n3239) );
  OAI21_X0P5M_A12TR u3360 ( .A0(n3819), .A1(n2870), .B0(n4157), .Y(n2523) );
  MXIT2_X0P5M_A12TR u3361 ( .A(n4158), .B(n3425), .S0(n2875), .Y(n4157) );
  INV_X0P5B_A12TR u3362 ( .A(n2497), .Y(n3425) );
  OAI211_X0P5M_A12TR u3363 ( .A0(n2876), .A1(n3253), .B0(n4159), .C0(n4160), 
        .Y(n4158) );
  AOI222_X0P5M_A12TR u3364 ( .A0(r1226_sum_9_), .A1(n2825), .B0(n2880), .B1(
        n1176), .C0(n2881), .C1(pc[9]), .Y(n4160) );
  AOI22_X0P5M_A12TR u3365 ( .A0(n2882), .A1(regfil_2__1_), .B0(n30180), .B1(
        n2883), .Y(n4159) );
  OAI21_X0P5M_A12TR u3366 ( .A0(n3825), .A1(n2870), .B0(n4161), .Y(n2522) );
  MXIT2_X0P5M_A12TR u3367 ( .A(n4162), .B(n3437), .S0(n2875), .Y(n4161) );
  INV_X0P5B_A12TR u3368 ( .A(n2496), .Y(n3437) );
  OAI211_X0P5M_A12TR u3369 ( .A0(n2876), .A1(n3258), .B0(n4163), .C0(n4164), 
        .Y(n4162) );
  AOI222_X0P5M_A12TR u3370 ( .A0(r1226_sum_10_), .A1(n2825), .B0(n2880), .B1(
        n1177), .C0(n2881), .C1(pc[10]), .Y(n4164) );
  AOI22_X0P5M_A12TR u3371 ( .A0(n2882), .A1(regfil_2__2_), .B0(n30190), .B1(
        n2883), .Y(n4163) );
  OAI21_X0P5M_A12TR u3372 ( .A0(n3831), .A1(n2870), .B0(n4165), .Y(n2521) );
  MXIT2_X0P5M_A12TR u3373 ( .A(n4166), .B(n3450), .S0(n2875), .Y(n4165) );
  INV_X0P5B_A12TR u3374 ( .A(n2495), .Y(n3450) );
  OAI211_X0P5M_A12TR u3375 ( .A0(n3263), .A1(n2876), .B0(n4167), .C0(n4168), 
        .Y(n4166) );
  AOI222_X0P5M_A12TR u3376 ( .A0(r1226_sum_11_), .A1(n2825), .B0(n2880), .B1(
        n1178), .C0(n2881), .C1(pc[11]), .Y(n4168) );
  AOI22_X0P5M_A12TR u3377 ( .A0(n2882), .A1(regfil_2__3_), .B0(n30200), .B1(
        n2883), .Y(n4167) );
  OAI21_X0P5M_A12TR u3378 ( .A0(n3837), .A1(n2870), .B0(n4169), .Y(n2520) );
  MXIT2_X0P5M_A12TR u3379 ( .A(n4170), .B(n3461), .S0(n2875), .Y(n4169) );
  INV_X0P5B_A12TR u3380 ( .A(n2494), .Y(n3461) );
  OAI211_X0P5M_A12TR u3381 ( .A0(n2876), .A1(n3268), .B0(n4171), .C0(n4172), 
        .Y(n4170) );
  AOI222_X0P5M_A12TR u3382 ( .A0(r1226_sum_12_), .A1(n2825), .B0(n2880), .B1(
        n1179), .C0(n2881), .C1(pc[12]), .Y(n4172) );
  AOI22_X0P5M_A12TR u3383 ( .A0(n2882), .A1(regfil_2__4_), .B0(n30210), .B1(
        n2883), .Y(n4171) );
  OAI21_X0P5M_A12TR u3384 ( .A0(n3843), .A1(n2870), .B0(n4173), .Y(n2519) );
  MXIT2_X0P5M_A12TR u3385 ( .A(n4174), .B(n3473), .S0(n2875), .Y(n4173) );
  INV_X0P5B_A12TR u3386 ( .A(n2493), .Y(n3473) );
  OAI211_X0P5M_A12TR u3387 ( .A0(n2876), .A1(n3273), .B0(n4175), .C0(n4176), 
        .Y(n4174) );
  AOI222_X0P5M_A12TR u3388 ( .A0(r1226_sum_13_), .A1(n2825), .B0(n2880), .B1(
        n1180), .C0(n2881), .C1(pc[13]), .Y(n4176) );
  AOI22_X0P5M_A12TR u3389 ( .A0(n2882), .A1(regfil_2__5_), .B0(n30220), .B1(
        n2883), .Y(n4175) );
  OAI21_X0P5M_A12TR u3390 ( .A0(n3849), .A1(n2870), .B0(n4177), .Y(n2518) );
  MXIT2_X0P5M_A12TR u3391 ( .A(n4178), .B(n3485), .S0(n2875), .Y(n4177) );
  INV_X0P5B_A12TR u3392 ( .A(n2492), .Y(n3485) );
  OAI211_X0P5M_A12TR u3393 ( .A0(n2876), .A1(n3278), .B0(n4179), .C0(n4180), 
        .Y(n4178) );
  AOI222_X0P5M_A12TR u3394 ( .A0(r1226_sum_14_), .A1(n2825), .B0(n2880), .B1(
        n1181), .C0(n2881), .C1(pc[14]), .Y(n4180) );
  AOI22_X0P5M_A12TR u3395 ( .A0(n2882), .A1(regfil_2__6_), .B0(n30230), .B1(
        n2883), .Y(n4179) );
  OAI21_X0P5M_A12TR u3396 ( .A0(n2960), .A1(n2870), .B0(n4181), .Y(n2517) );
  MXIT2_X0P5M_A12TR u3397 ( .A(n4182), .B(n2895), .S0(n2875), .Y(n4181) );
  INV_X0P5B_A12TR u3398 ( .A(n4183), .Y(n2875) );
  INV_X0P5B_A12TR u3399 ( .A(n2491), .Y(n2895) );
  OAI211_X0P5M_A12TR u3400 ( .A0(n2830), .A1(n2876), .B0(n4184), .C0(n4185), 
        .Y(n4182) );
  AOI222_X0P5M_A12TR u3401 ( .A0(r1226_sum_15_), .A1(n2825), .B0(n2880), .B1(
        n1182), .C0(n2881), .C1(pc[15]), .Y(n4185) );
  NOR2_X0P5A_A12TR u3402 ( .A(n3331), .B(n3568), .Y(n2881) );
  NOR2_X0P5A_A12TR u3403 ( .A(n3356), .B(n2829), .Y(n2880) );
  AOI22_X0P5M_A12TR u3404 ( .A0(n2882), .A1(regfil_2__7_), .B0(n30240), .B1(
        n2883), .Y(n4184) );
  OAI21_X0P5M_A12TR u3405 ( .A0(intcyc), .A1(n3568), .B0(n3191), .Y(n2883) );
  NOR2_X0P5A_A12TR u3406 ( .A(n3356), .B(n2831), .Y(n2882) );
  NAND2_X0P5A_A12TR u3407 ( .A(n3984), .B(n2983), .Y(n2876) );
  INV_X0P5B_A12TR u3408 ( .A(n3356), .Y(n3984) );
  OAI21_X0P5M_A12TR u3409 ( .A0(n3127), .A1(n2901), .B0(n4183), .Y(n2870) );
  OAI22_X0P5M_A12TR u3410 ( .A0(n4156), .A1(n3298), .B0(n3395), .B1(n3312), 
        .Y(n4183) );
  NAND2B_X0P5M_A12TR u3411 ( .AN(n3298), .B(n3127), .Y(n3312) );
  NAND2_X0P5A_A12TR u3412 ( .A(n3855), .B(n3181), .Y(n3298) );
  INV_X0P5B_A12TR u3413 ( .A(n3229), .Y(n3855) );
  NAND3_X0P5A_A12TR u3414 ( .A(n2823), .B(n3004), .C(n3074), .Y(n3229) );
  INV_X0P5B_A12TR u3415 ( .A(n3604), .Y(n3074) );
  NAND3_X0P5A_A12TR u3416 ( .A(n30131), .B(n30111), .C(state[2]), .Y(n3604) );
  AOI211_X0P5M_A12TR u3417 ( .A0(r1298_carry_1_), .A1(n3366), .B0(n4055), .C0(
        n3351), .Y(n4156) );
  NOR2_X0P5A_A12TR u3418 ( .A(n2869), .B(n3193), .Y(n3351) );
  INV_X0P5B_A12TR u3419 ( .A(n3357), .Y(n4055) );
  OAI21_X0P5M_A12TR u3420 ( .A0(n3042), .A1(n3356), .B0(n2869), .Y(n2901) );
  OAI221_X0P5M_A12TR u3421 ( .A0(n2838), .A1(n4186), .B0(n2837), .B1(n4187), 
        .C0(n4188), .Y(n2516) );
  AOI22_X0P5M_A12TR u3422 ( .A0(n4189), .A1(n4151), .B0(addr[15]), .B1(n4190), 
        .Y(n4188) );
  INV_X0P5B_A12TR u3423 ( .A(n2467), .Y(n4151) );
  INV_X0P5B_A12TR u3424 ( .A(raddrhold[15]), .Y(n2838) );
  OAI221_X0P5M_A12TR u3425 ( .A0(n2841), .A1(n4186), .B0(n2840), .B1(n4187), 
        .C0(n4191), .Y(n2515) );
  AOI22_X0P5M_A12TR u3426 ( .A0(n4189), .A1(n4143), .B0(addr[14]), .B1(n4190), 
        .Y(n4191) );
  INV_X0P5B_A12TR u3427 ( .A(n2468), .Y(n4143) );
  INV_X0P5B_A12TR u3428 ( .A(raddrhold[14]), .Y(n2841) );
  OAI221_X0P5M_A12TR u3429 ( .A0(n2844), .A1(n4186), .B0(n2843), .B1(n4187), 
        .C0(n4192), .Y(n2514) );
  AOI22_X0P5M_A12TR u3430 ( .A0(n4189), .A1(n4138), .B0(addr[13]), .B1(n4190), 
        .Y(n4192) );
  INV_X0P5B_A12TR u3431 ( .A(n2469), .Y(n4138) );
  INV_X0P5B_A12TR u3432 ( .A(raddrhold[13]), .Y(n2844) );
  OAI221_X0P5M_A12TR u3433 ( .A0(n2847), .A1(n4186), .B0(n2846), .B1(n4187), 
        .C0(n4193), .Y(n2513) );
  AOI22_X0P5M_A12TR u3434 ( .A0(n4189), .A1(n4133), .B0(addr[12]), .B1(n4190), 
        .Y(n4193) );
  INV_X0P5B_A12TR u3435 ( .A(n2470), .Y(n4133) );
  INV_X0P5B_A12TR u3436 ( .A(raddrhold[12]), .Y(n2847) );
  OAI221_X0P5M_A12TR u3437 ( .A0(n2850), .A1(n4186), .B0(n2849), .B1(n4187), 
        .C0(n4194), .Y(n2512) );
  AOI22_X0P5M_A12TR u3438 ( .A0(n4189), .A1(n4128), .B0(addr[11]), .B1(n4190), 
        .Y(n4194) );
  INV_X0P5B_A12TR u3439 ( .A(n2471), .Y(n4128) );
  INV_X0P5B_A12TR u3440 ( .A(raddrhold[11]), .Y(n2850) );
  OAI221_X0P5M_A12TR u3441 ( .A0(n2853), .A1(n4186), .B0(n2852), .B1(n4187), 
        .C0(n4195), .Y(n2511) );
  AOI22_X0P5M_A12TR u3442 ( .A0(n4189), .A1(n4123), .B0(addr[10]), .B1(n4190), 
        .Y(n4195) );
  INV_X0P5B_A12TR u3443 ( .A(n2472), .Y(n4123) );
  INV_X0P5B_A12TR u3444 ( .A(raddrhold[10]), .Y(n2853) );
  OAI221_X0P5M_A12TR u3445 ( .A0(n2835), .A1(n4186), .B0(n2834), .B1(n4187), 
        .C0(n4196), .Y(n2510) );
  AOI22_X0P5M_A12TR u3446 ( .A0(n4189), .A1(n4118), .B0(addr[9]), .B1(n4190), 
        .Y(n4196) );
  INV_X0P5B_A12TR u3447 ( .A(n2473), .Y(n4118) );
  INV_X0P5B_A12TR u3448 ( .A(raddrhold[9]), .Y(n2835) );
  OAI221_X0P5M_A12TR u3449 ( .A0(n4197), .A1(n4186), .B0(n3947), .B1(n4187), 
        .C0(n4198), .Y(n2509) );
  AOI22_X0P5M_A12TR u3450 ( .A0(n4189), .A1(n4113), .B0(addr[8]), .B1(n4190), 
        .Y(n4198) );
  INV_X0P5B_A12TR u3451 ( .A(n2474), .Y(n4113) );
  INV_X0P5B_A12TR u3452 ( .A(n4199), .Y(n4187) );
  INV_X0P5B_A12TR u3453 ( .A(n4200), .Y(n4186) );
  OAI211_X0P5M_A12TR u3454 ( .A0(n2912), .A1(n4201), .B0(n4202), .C0(n4203), 
        .Y(n2508) );
  AOI22_X0P5M_A12TR u3455 ( .A0(n4189), .A1(n4108), .B0(addr[7]), .B1(n4190), 
        .Y(n4203) );
  INV_X0P5B_A12TR u3456 ( .A(n2475), .Y(n4108) );
  AOI22_X0P5M_A12TR u3457 ( .A0(n4200), .A1(raddrhold[7]), .B0(n4199), .B1(
        pc[7]), .Y(n4202) );
  INV_X0P5B_A12TR u3458 ( .A(rdatahold[7]), .Y(n2912) );
  OAI211_X0P5M_A12TR u3459 ( .A0(n3283), .A1(n4201), .B0(n4204), .C0(n4205), 
        .Y(n2507) );
  AOI22_X0P5M_A12TR u3460 ( .A0(n4189), .A1(n4103), .B0(addr[6]), .B1(n4190), 
        .Y(n4205) );
  INV_X0P5B_A12TR u3461 ( .A(n2476), .Y(n4103) );
  AOI22_X0P5M_A12TR u3462 ( .A0(n4200), .A1(raddrhold[6]), .B0(n4199), .B1(
        pc[6]), .Y(n4204) );
  INV_X0P5B_A12TR u3463 ( .A(rdatahold[6]), .Y(n3283) );
  OAI211_X0P5M_A12TR u3464 ( .A0(n3275), .A1(n4201), .B0(n4206), .C0(n4207), 
        .Y(n2506) );
  AOI22_X0P5M_A12TR u3465 ( .A0(n4189), .A1(n4098), .B0(addr[5]), .B1(n4190), 
        .Y(n4207) );
  INV_X0P5B_A12TR u3466 ( .A(n2477), .Y(n4098) );
  AOI22_X0P5M_A12TR u3467 ( .A0(n4200), .A1(raddrhold[5]), .B0(n4199), .B1(
        pc[5]), .Y(n4206) );
  INV_X0P5B_A12TR u3468 ( .A(rdatahold[5]), .Y(n3275) );
  OAI211_X0P5M_A12TR u3469 ( .A0(n3270), .A1(n4201), .B0(n4208), .C0(n4209), 
        .Y(n2505) );
  AOI22_X0P5M_A12TR u3470 ( .A0(n4189), .A1(n4093), .B0(addr[4]), .B1(n4190), 
        .Y(n4209) );
  INV_X0P5B_A12TR u3471 ( .A(n2478), .Y(n4093) );
  AOI22_X0P5M_A12TR u3472 ( .A0(n4200), .A1(raddrhold[4]), .B0(n4199), .B1(
        pc[4]), .Y(n4208) );
  INV_X0P5B_A12TR u3473 ( .A(rdatahold[4]), .Y(n3270) );
  OAI211_X0P5M_A12TR u3474 ( .A0(n3265), .A1(n4201), .B0(n4210), .C0(n4211), 
        .Y(n2504) );
  AOI22_X0P5M_A12TR u3475 ( .A0(n4189), .A1(n4088), .B0(addr[3]), .B1(n4190), 
        .Y(n4211) );
  INV_X0P5B_A12TR u3476 ( .A(n2479), .Y(n4088) );
  AOI22_X0P5M_A12TR u3477 ( .A0(n4200), .A1(raddrhold[3]), .B0(n4199), .B1(
        pc[3]), .Y(n4210) );
  INV_X0P5B_A12TR u3478 ( .A(rdatahold[3]), .Y(n3265) );
  OAI211_X0P5M_A12TR u3479 ( .A0(n3260), .A1(n4201), .B0(n4212), .C0(n4213), 
        .Y(n2503) );
  AOI22_X0P5M_A12TR u3480 ( .A0(n4189), .A1(n4083), .B0(addr[2]), .B1(n4190), 
        .Y(n4213) );
  INV_X0P5B_A12TR u3481 ( .A(n2480), .Y(n4083) );
  AOI22_X0P5M_A12TR u3482 ( .A0(n4200), .A1(raddrhold[2]), .B0(n4199), .B1(
        pc[2]), .Y(n4212) );
  INV_X0P5B_A12TR u3483 ( .A(rdatahold[2]), .Y(n3260) );
  OAI211_X0P5M_A12TR u3484 ( .A0(n3255), .A1(n4201), .B0(n4214), .C0(n4215), 
        .Y(n2502) );
  AOI22_X0P5M_A12TR u3485 ( .A0(n4189), .A1(n4076), .B0(addr[1]), .B1(n4190), 
        .Y(n4215) );
  INV_X0P5B_A12TR u3486 ( .A(n2481), .Y(n4076) );
  AOI22_X0P5M_A12TR u3487 ( .A0(n4200), .A1(raddrhold[1]), .B0(n4199), .B1(
        pc[1]), .Y(n4214) );
  INV_X0P5B_A12TR u3488 ( .A(rdatahold[1]), .Y(n3255) );
  OAI211_X0P5M_A12TR u3489 ( .A0(n3251), .A1(n4201), .B0(n4216), .C0(n4217), 
        .Y(n2501) );
  AOI22_X0P5M_A12TR u3490 ( .A0(n4189), .A1(n4218), .B0(addr[0]), .B1(n4190), 
        .Y(n4217) );
  INV_X0P5B_A12TR u3491 ( .A(n2482), .Y(n4218) );
  NOR3_X0P5A_A12TR u3492 ( .A(n3153), .B(n2823), .C(n4190), .Y(n4189) );
  AOI22_X0P5M_A12TR u3493 ( .A0(n4200), .A1(raddrhold[0]), .B0(n4199), .B1(
        pc[0]), .Y(n4216) );
  NOR3_X0P5A_A12TR u3494 ( .A(u3_u93_z_6), .B(state[3]), .C(n4190), .Y(n4199)
         );
  NOR2_X0P5A_A12TR u3495 ( .A(n4190), .B(n3231), .Y(n4200) );
  INV_X0P5B_A12TR u3496 ( .A(n4219), .Y(n4201) );
  OA21A1OI2_X0P5M_A12TR u3497 ( .A0(n2972), .A1(state[3]), .B0(n3730), .C0(
        n4190), .Y(n4219) );
  OAI31_X0P5M_A12TR u3498 ( .A0(n4220), .A1(n4221), .A2(n3565), .B0(n3181), 
        .Y(n4190) );
  NOR2B_X0P5M_A12TR u3499 ( .AN(n3078), .B(n3086), .Y(n3565) );
  NOR2_X0P5A_A12TR u3500 ( .A(n4222), .B(state[2]), .Y(n3078) );
  INV_X0P5B_A12TR u3501 ( .A(n3084), .Y(n4221) );
  NAND3_X0P5A_A12TR u3502 ( .A(state[2]), .B(n3087), .C(n30161), .Y(n3084) );
  INV_X0P5B_A12TR u3503 ( .A(n4222), .Y(n30161) );
  NOR2_X0P5A_A12TR u3504 ( .A(n3166), .B(n3087), .Y(n4220) );
  NAND2_X0P5A_A12TR u3505 ( .A(n3086), .B(n30141), .Y(n3087) );
  NAND2_X0P5A_A12TR u3506 ( .A(state[3]), .B(n3179), .Y(n30141) );
  NAND2_X0P5A_A12TR u3507 ( .A(state[0]), .B(state[3]), .Y(n3730) );
  INV_X0P5B_A12TR u3508 ( .A(rdatahold[0]), .Y(n3251) );
  OAI31_X0P5M_A12TR u3509 ( .A0(n3086), .A1(n3492), .A2(n4222), .B0(n4223), 
        .Y(n2500) );
  NAND3B_X0P5M_A12TR u3510 ( .AN(n3653), .B(n3181), .C(readio), .Y(n4223) );
  AND3_X0P5M_A12TR u3511 ( .A(n3155), .B(n3233), .C(n3241), .Y(n3653) );
  NOR2B_X0P5M_A12TR u3512 ( .AN(n2859), .B(n3070), .Y(n3241) );
  NAND2_X0P5A_A12TR u3513 ( .A(n3004), .B(n2972), .Y(n3070) );
  INV_X0P5B_A12TR u3514 ( .A(n30171), .Y(n3155) );
  NAND2_X0P5A_A12TR u3515 ( .A(state[4]), .B(state[3]), .Y(n30171) );
  NAND2_X0P5A_A12TR u3516 ( .A(n3226), .B(n30111), .Y(n4222) );
  NAND2_X0P5A_A12TR u3517 ( .A(n2971), .B(n3181), .Y(n3492) );
  INV_X0P5B_A12TR u3518 ( .A(n2914), .Y(n2971) );
  NAND2_X0P5A_A12TR u3519 ( .A(state[2]), .B(u3_u93_z_6), .Y(n2914) );
  MXIT2_X0P5M_A12TR u3520 ( .A(n3333), .B(n2456), .S0(n4224), .Y(n2499) );
  NOR2_X0P5A_A12TR u3521 ( .A(n3335), .B(n4225), .Y(n4224) );
  OAI31_X0P5M_A12TR u3522 ( .A0(n3210), .A1(n3331), .A2(n3337), .B0(n3332), 
        .Y(n4225) );
  INV_X0P5B_A12TR u3523 ( .A(n3327), .Y(n3332) );
  NOR2_X0P5A_A12TR u3524 ( .A(n3134), .B(n3328), .Y(n3327) );
  INV_X0P5B_A12TR u3525 ( .A(n3322), .Y(n3328) );
  NOR2_X0P5A_A12TR u3526 ( .A(n3166), .B(n3295), .Y(n3322) );
  NAND3_X0P5A_A12TR u3527 ( .A(n2859), .B(n2972), .C(state[0]), .Y(n3166) );
  NAND2_X0P5A_A12TR u3528 ( .A(intr), .B(ei), .Y(n3134) );
  INV_X0P5B_A12TR u3529 ( .A(intcyc), .Y(n3331) );
  NAND2_X0P5A_A12TR u3530 ( .A(n31401), .B(n3004), .Y(n3210) );
  OAI211_X0P5M_A12TR u3531 ( .A0(n3168), .A1(n3242), .B0(n4226), .C0(n3181), 
        .Y(n3335) );
  NAND4_X0P5A_A12TR u3532 ( .A(n3246), .B(state[0]), .C(n30131), .D(n3233), 
        .Y(n4226) );
  INV_X0P5B_A12TR u3533 ( .A(n3295), .Y(n30131) );
  NAND2_X0P5A_A12TR u3534 ( .A(n3179), .B(n3153), .Y(n3295) );
  INV_X0P5B_A12TR u3535 ( .A(n3337), .Y(n3246) );
  NAND2_X0P5A_A12TR u3536 ( .A(n3075), .B(n30111), .Y(n3337) );
  INV_X0P5B_A12TR u3537 ( .A(n3231), .Y(n3075) );
  NAND2_X0P5A_A12TR u3538 ( .A(u3_u93_z_6), .B(n2972), .Y(n3231) );
  INV_X0P5B_A12TR u3539 ( .A(state[2]), .Y(n2972) );
  NAND2_X0P5A_A12TR u3540 ( .A(n31401), .B(n3233), .Y(n3242) );
  INV_X0P5B_A12TR u3541 ( .A(waitr), .Y(n3233) );
  INV_X0P5B_A12TR u3542 ( .A(n3086), .Y(n31401) );
  NAND2_X0P5A_A12TR u3543 ( .A(state[4]), .B(n3153), .Y(n3086) );
  INV_X0P5B_A12TR u3544 ( .A(state[3]), .Y(n3153) );
  NAND2_X0P5A_A12TR u3545 ( .A(n3088), .B(n2859), .Y(n3168) );
  INV_X0P5B_A12TR u3546 ( .A(n30191), .Y(n3088) );
  NAND2_X0P5A_A12TR u3547 ( .A(state[2]), .B(n3004), .Y(n30191) );
  AO21A1AI2_X0P5M_A12TR u3548 ( .A0(n3179), .A1(n2823), .B0(n3226), .C0(n3181), 
        .Y(n3333) );
  INV_X0P5B_A12TR u3549 ( .A(reset), .Y(n3181) );
  INV_X0P5B_A12TR u3550 ( .A(n3646), .Y(n3226) );
  NAND2_X0P5A_A12TR u3551 ( .A(u3_u93_z_6), .B(n3004), .Y(n3646) );
  INV_X0P5B_A12TR u3552 ( .A(state[0]), .Y(n3004) );
  INV_X0P5B_A12TR u3553 ( .A(state[4]), .Y(n3179) );
  OAI211_X0P5M_A12TR u3554 ( .A0(n4227), .A1(n2829), .B0(n4228), .C0(n4229), 
        .Y(u3_u94_z_0) );
  OAI221_X0P5M_A12TR u3555 ( .A0(n4230), .A1(n2830), .B0(n3594), .B1(n4231), 
        .C0(n4232), .Y(u3_u92_z_7) );
  AOI22_X0P5M_A12TR u3556 ( .A0(n1157), .A1(n4233), .B0(n1664), .B1(n4234), 
        .Y(n4232) );
  OAI221_X0P5M_A12TR u3557 ( .A0(n4230), .A1(n3278), .B0(n3876), .B1(n4231), 
        .C0(n4235), .Y(u3_u92_z_6) );
  AOI22_X0P5M_A12TR u3558 ( .A0(n1156), .A1(n4233), .B0(n1663), .B1(n4234), 
        .Y(n4235) );
  OAI221_X0P5M_A12TR u3559 ( .A0(n4230), .A1(n3273), .B0(n3873), .B1(n4231), 
        .C0(n4236), .Y(u3_u92_z_5) );
  AOI22_X0P5M_A12TR u3560 ( .A0(n1155), .A1(n4233), .B0(n1662), .B1(n4234), 
        .Y(n4236) );
  OAI221_X0P5M_A12TR u3561 ( .A0(n4230), .A1(n3268), .B0(n3870), .B1(n4231), 
        .C0(n4237), .Y(u3_u92_z_4) );
  AOI22_X0P5M_A12TR u3562 ( .A0(n1154), .A1(n4233), .B0(n1661), .B1(n4234), 
        .Y(n4237) );
  OAI221_X0P5M_A12TR u3563 ( .A0(n4230), .A1(n3263), .B0(n3867), .B1(n4231), 
        .C0(n4238), .Y(u3_u92_z_3) );
  AOI22_X0P5M_A12TR u3564 ( .A0(n1153), .A1(n4233), .B0(n1660), .B1(n4234), 
        .Y(n4238) );
  OAI221_X0P5M_A12TR u3565 ( .A0(n4230), .A1(n3258), .B0(n3864), .B1(n4231), 
        .C0(n4239), .Y(u3_u92_z_2) );
  AOI22_X0P5M_A12TR u3566 ( .A0(n1152), .A1(n4233), .B0(n1659), .B1(n4234), 
        .Y(n4239) );
  OAI221_X0P5M_A12TR u3567 ( .A0(n4230), .A1(n3253), .B0(n3861), .B1(n4231), 
        .C0(n4240), .Y(u3_u92_z_1) );
  AOI22_X0P5M_A12TR u3568 ( .A0(n1151), .A1(n4233), .B0(n1658), .B1(n4234), 
        .Y(n4240) );
  OAI221_X0P5M_A12TR u3569 ( .A0(n4230), .A1(n2877), .B0(n3858), .B1(n4231), 
        .C0(n4241), .Y(u3_u92_z_0) );
  AOI22_X0P5M_A12TR u3570 ( .A0(n1150), .A1(n4233), .B0(n1657), .B1(n4234), 
        .Y(n4241) );
  NAND2_X0P5A_A12TR u3571 ( .A(n2823), .B(n3899), .Y(n4231) );
  AOI21_X0P5M_A12TR u3572 ( .A0(n2866), .A1(n2865), .B0(u3_u93_z_6), .Y(n4230)
         );
  NAND2_X0P5A_A12TR u3573 ( .A(n3649), .B(n3600), .Y(n2866) );
  INV_X0P5B_A12TR u3574 ( .A(auxcar), .Y(n3600) );
  MXT2_X0P5M_A12TR u3575 ( .A(n4242), .B(n4243), .S0(n2823), .Y(n3649) );
  OAI21_X0P5M_A12TR u3576 ( .A0(n1103), .A1(n1102), .B0(n1104), .Y(n4243) );
  OAI21_X0P5M_A12TR u3577 ( .A0(n1107), .A1(n1106), .B0(n1108), .Y(n4242) );
  OAI222_X0P5M_A12TR u3578 ( .A0(n2833), .A1(n2862), .B0(n2834), .B1(n2863), 
        .C0(n4244), .C1(n4245), .Y(u3_u88_z_9) );
  OAI222_X0P5M_A12TR u3579 ( .A0(n4246), .A1(n2862), .B0(n3947), .B1(n2863), 
        .C0(n4244), .C1(n4247), .Y(u3_u88_z_8) );
  OAI222_X0P5M_A12TR u3580 ( .A0(n4248), .A1(n2862), .B0(n3943), .B1(n2863), 
        .C0(n4244), .C1(n4249), .Y(u3_u88_z_7) );
  OAI222_X0P5M_A12TR u3581 ( .A0(n4250), .A1(n2862), .B0(n3939), .B1(n2863), 
        .C0(n4244), .C1(n4251), .Y(u3_u88_z_6) );
  OAI222_X0P5M_A12TR u3582 ( .A0(n4252), .A1(n2862), .B0(n3474), .B1(n2863), 
        .C0(n4244), .C1(n4253), .Y(u3_u88_z_5) );
  OAI222_X0P5M_A12TR u3583 ( .A0(n4254), .A1(n2862), .B0(n4255), .B1(n2863), 
        .C0(n4244), .C1(n4256), .Y(u3_u88_z_4) );
  OAI222_X0P5M_A12TR u3584 ( .A0(n4257), .A1(n2862), .B0(n3452), .B1(n2863), 
        .C0(n4244), .C1(n4258), .Y(u3_u88_z_3) );
  OAI222_X0P5M_A12TR u3585 ( .A0(n4259), .A1(n2862), .B0(n3909), .B1(n2863), 
        .C0(n4244), .C1(n4260), .Y(u3_u88_z_2) );
  OAI222_X0P5M_A12TR u3586 ( .A0(n2836), .A1(n2862), .B0(n2837), .B1(n2863), 
        .C0(n4244), .C1(n4261), .Y(u3_u88_z_15) );
  OAI222_X0P5M_A12TR u3587 ( .A0(n2839), .A1(n2862), .B0(n2840), .B1(n2863), 
        .C0(n4244), .C1(n4262), .Y(u3_u88_z_14) );
  OAI222_X0P5M_A12TR u3588 ( .A0(n2842), .A1(n2862), .B0(n2843), .B1(n2863), 
        .C0(n4244), .C1(n4263), .Y(u3_u88_z_13) );
  OAI222_X0P5M_A12TR u3589 ( .A0(n2845), .A1(n2862), .B0(n2846), .B1(n2863), 
        .C0(n4244), .C1(n4264), .Y(u3_u88_z_12) );
  OAI222_X0P5M_A12TR u3590 ( .A0(n2848), .A1(n2862), .B0(n2849), .B1(n2863), 
        .C0(n4244), .C1(n4265), .Y(u3_u88_z_11) );
  OAI222_X0P5M_A12TR u3591 ( .A0(n2851), .A1(n2862), .B0(n2852), .B1(n2863), 
        .C0(n4244), .C1(n4266), .Y(u3_u88_z_10) );
  OAI222_X0P5M_A12TR u3592 ( .A0(n4267), .A1(n2862), .B0(n3905), .B1(n2863), 
        .C0(n4244), .C1(n4078), .Y(u3_u88_z_1) );
  OAI222_X0P5M_A12TR u3593 ( .A0(n2854), .A1(n2862), .B0(n2855), .B1(n2863), 
        .C0(n4244), .C1(n4268), .Y(u3_u88_z_0) );
  AND2_X0P5M_A12TR u3594 ( .A(n2859), .B(n2861), .Y(n4244) );
  NOR2_X0P5A_A12TR u3595 ( .A(state[5]), .B(u3_u93_z_6), .Y(n2859) );
  NAND2_X0P5A_A12TR u3596 ( .A(n30111), .B(n2858), .Y(n2863) );
  NAND3_X0P5A_A12TR u3597 ( .A(n3988), .B(n3395), .C(n4269), .Y(n2858) );
  NAND2_X0P5A_A12TR u3598 ( .A(n3350), .B(n30111), .Y(n2862) );
  INV_X0P5B_A12TR u3599 ( .A(state[5]), .Y(n30111) );
  OAI221_X0P5M_A12TR u3600 ( .A0(n2820), .A1(n3947), .B0(n2830), .B1(n4270), 
        .C0(n4271), .Y(u3_u85_z_8) );
  OA22_X0P5M_A12TR u3601 ( .A0(n4246), .A1(n2824), .B0(n4197), .B1(n2823), .Y(
        n4271) );
  INV_X0P5B_A12TR u3602 ( .A(raddrhold[8]), .Y(n4197) );
  INV_X0P5B_A12TR u3603 ( .A(n1108), .Y(n2830) );
  OAI221_X0P5M_A12TR u3604 ( .A0(n2820), .A1(n3943), .B0(n3278), .B1(n4270), 
        .C0(n4272), .Y(u3_u85_z_7) );
  AOI22_X0P5M_A12TR u3605 ( .A0(n4273), .A1(n4274), .B0(raddrhold[7]), .B1(
        u3_u93_z_6), .Y(n4272) );
  INV_X0P5B_A12TR u3606 ( .A(n4248), .Y(n4273) );
  INV_X0P5B_A12TR u3607 ( .A(n1107), .Y(n3278) );
  OAI221_X0P5M_A12TR u3608 ( .A0(n2820), .A1(n3939), .B0(n3273), .B1(n4270), 
        .C0(n4275), .Y(u3_u85_z_6) );
  AOI22_X0P5M_A12TR u3609 ( .A0(n4276), .A1(n4274), .B0(raddrhold[6]), .B1(
        u3_u93_z_6), .Y(n4275) );
  INV_X0P5B_A12TR u3610 ( .A(n4250), .Y(n4276) );
  INV_X0P5B_A12TR u3611 ( .A(n1106), .Y(n3273) );
  OAI221_X0P5M_A12TR u3612 ( .A0(n2820), .A1(n3474), .B0(n3268), .B1(n4270), 
        .C0(n4277), .Y(u3_u85_z_5) );
  AOI22_X0P5M_A12TR u3613 ( .A0(n4278), .A1(n4274), .B0(raddrhold[5]), .B1(
        u3_u93_z_6), .Y(n4277) );
  INV_X0P5B_A12TR u3614 ( .A(n4252), .Y(n4278) );
  INV_X0P5B_A12TR u3615 ( .A(n1105), .Y(n3268) );
  OAI221_X0P5M_A12TR u3616 ( .A0(n2820), .A1(n4255), .B0(n3263), .B1(n4270), 
        .C0(n4279), .Y(u3_u85_z_4) );
  AOI22_X0P5M_A12TR u3617 ( .A0(n4280), .A1(n4274), .B0(raddrhold[4]), .B1(
        u3_u93_z_6), .Y(n4279) );
  INV_X0P5B_A12TR u3618 ( .A(n4254), .Y(n4280) );
  INV_X0P5B_A12TR u3619 ( .A(n1104), .Y(n3263) );
  OAI221_X0P5M_A12TR u3620 ( .A0(n2820), .A1(n3452), .B0(n3258), .B1(n4270), 
        .C0(n4281), .Y(u3_u85_z_3) );
  AOI22_X0P5M_A12TR u3621 ( .A0(n4282), .A1(n4274), .B0(raddrhold[3]), .B1(
        u3_u93_z_6), .Y(n4281) );
  INV_X0P5B_A12TR u3622 ( .A(n4257), .Y(n4282) );
  INV_X0P5B_A12TR u3623 ( .A(n1103), .Y(n3258) );
  OAI221_X0P5M_A12TR u3624 ( .A0(n2820), .A1(n3909), .B0(n3253), .B1(n4270), 
        .C0(n4283), .Y(u3_u85_z_2) );
  AOI22_X0P5M_A12TR u3625 ( .A0(n4284), .A1(n4274), .B0(raddrhold[2]), .B1(
        u3_u93_z_6), .Y(n4283) );
  INV_X0P5B_A12TR u3626 ( .A(n4259), .Y(n4284) );
  INV_X0P5B_A12TR u3627 ( .A(n1102), .Y(n3253) );
  OAI221_X0P5M_A12TR u3628 ( .A0(n2820), .A1(n3905), .B0(n2877), .B1(n4270), 
        .C0(n4285), .Y(u3_u85_z_1) );
  AOI22_X0P5M_A12TR u3629 ( .A0(n4286), .A1(n4274), .B0(raddrhold[1]), .B1(
        u3_u93_z_6), .Y(n4285) );
  INV_X0P5B_A12TR u3630 ( .A(n4267), .Y(n4286) );
  INV_X0P5B_A12TR u3631 ( .A(regfil_7__0_), .Y(n2877) );
  OAI22_X0P5M_A12TR u3632 ( .A0(n2473), .A1(n2823), .B0(n4287), .B1(n2834), 
        .Y(u3_u84_z_9) );
  INV_X0P5B_A12TR u3633 ( .A(pc[9]), .Y(n2834) );
  OAI22_X0P5M_A12TR u3634 ( .A0(n2474), .A1(n2823), .B0(n4287), .B1(n3947), 
        .Y(u3_u84_z_8) );
  INV_X0P5B_A12TR u3635 ( .A(pc[8]), .Y(n3947) );
  OAI22_X0P5M_A12TR u3636 ( .A0(n2475), .A1(n2823), .B0(n4287), .B1(n3943), 
        .Y(u3_u84_z_7) );
  INV_X0P5B_A12TR u3637 ( .A(pc[7]), .Y(n3943) );
  OAI22_X0P5M_A12TR u3638 ( .A0(n2476), .A1(n2823), .B0(n4287), .B1(n3939), 
        .Y(u3_u84_z_6) );
  INV_X0P5B_A12TR u3639 ( .A(pc[6]), .Y(n3939) );
  OAI22_X0P5M_A12TR u3640 ( .A0(n2477), .A1(n2823), .B0(n4287), .B1(n3474), 
        .Y(u3_u84_z_5) );
  INV_X0P5B_A12TR u3641 ( .A(pc[5]), .Y(n3474) );
  OAI22_X0P5M_A12TR u3642 ( .A0(n2478), .A1(n2823), .B0(n4287), .B1(n4255), 
        .Y(u3_u84_z_4) );
  INV_X0P5B_A12TR u3643 ( .A(pc[4]), .Y(n4255) );
  OAI22_X0P5M_A12TR u3644 ( .A0(n2479), .A1(n2823), .B0(n4287), .B1(n3452), 
        .Y(u3_u84_z_3) );
  INV_X0P5B_A12TR u3645 ( .A(pc[3]), .Y(n3452) );
  OAI22_X0P5M_A12TR u3646 ( .A0(n2480), .A1(n2823), .B0(n4287), .B1(n3909), 
        .Y(u3_u84_z_2) );
  INV_X0P5B_A12TR u3647 ( .A(pc[2]), .Y(n3909) );
  OAI22_X0P5M_A12TR u3648 ( .A0(n2467), .A1(n2823), .B0(n4287), .B1(n2837), 
        .Y(u3_u84_z_15) );
  INV_X0P5B_A12TR u3649 ( .A(pc[15]), .Y(n2837) );
  OAI22_X0P5M_A12TR u3650 ( .A0(n2468), .A1(n2823), .B0(n4287), .B1(n2840), 
        .Y(u3_u84_z_14) );
  INV_X0P5B_A12TR u3651 ( .A(pc[14]), .Y(n2840) );
  OAI22_X0P5M_A12TR u3652 ( .A0(n2469), .A1(n2823), .B0(n4287), .B1(n2843), 
        .Y(u3_u84_z_13) );
  INV_X0P5B_A12TR u3653 ( .A(pc[13]), .Y(n2843) );
  OAI22_X0P5M_A12TR u3654 ( .A0(n2470), .A1(n2823), .B0(n4287), .B1(n2846), 
        .Y(u3_u84_z_12) );
  INV_X0P5B_A12TR u3655 ( .A(pc[12]), .Y(n2846) );
  OAI22_X0P5M_A12TR u3656 ( .A0(n2471), .A1(n2823), .B0(n4287), .B1(n2849), 
        .Y(u3_u84_z_11) );
  INV_X0P5B_A12TR u3657 ( .A(pc[11]), .Y(n2849) );
  OAI22_X0P5M_A12TR u3658 ( .A0(n2472), .A1(n2823), .B0(n4287), .B1(n2852), 
        .Y(u3_u84_z_10) );
  INV_X0P5B_A12TR u3659 ( .A(pc[10]), .Y(n2852) );
  OAI22_X0P5M_A12TR u3660 ( .A0(n2481), .A1(n2823), .B0(n4287), .B1(n3905), 
        .Y(u3_u84_z_1) );
  INV_X0P5B_A12TR u3661 ( .A(pc[1]), .Y(n3905) );
  OAI22_X0P5M_A12TR u3662 ( .A0(n2482), .A1(n2823), .B0(n4287), .B1(n2855), 
        .Y(u3_u84_z_0) );
  INV_X0P5B_A12TR u3663 ( .A(pc[0]), .Y(n2855) );
  AND4_X0P5M_A12TR u3664 ( .A(n2824), .B(n2820), .C(n4288), .D(n4289), .Y(
        n4287) );
  AOI211_X0P5M_A12TR u3665 ( .A0(n2826), .A1(n4290), .B0(n4291), .C0(n4292), 
        .Y(n4289) );
  AOI21_X0P5M_A12TR u3666 ( .A0(n3357), .A1(n3111), .B0(u3_u93_z_6), .Y(n4292)
         );
  NAND2_X0P5A_A12TR u3667 ( .A(opcode[7]), .B(n3291), .Y(n3111) );
  NAND2_X0P5A_A12TR u3668 ( .A(n2825), .B(n3366), .Y(n3357) );
  NAND3_X0P5A_A12TR u3669 ( .A(n3484), .B(n4270), .C(n2890), .Y(n4291) );
  INV_X0P5B_A12TR u3670 ( .A(n3477), .Y(n2890) );
  NOR2_X0P5A_A12TR u3671 ( .A(n3395), .B(n3642), .Y(n3477) );
  NAND2_X0P5A_A12TR u3672 ( .A(n3125), .B(n3766), .Y(n3395) );
  NAND2_X0P5A_A12TR u3673 ( .A(n2924), .B(n2826), .Y(n4270) );
  NOR3_X0P5A_A12TR u3674 ( .A(n4293), .B(n236), .C(n3426), .Y(n2924) );
  NAND2_X0P5A_A12TR u3675 ( .A(n35711), .B(n2823), .Y(n3484) );
  INV_X0P5B_A12TR u3676 ( .A(n3228), .Y(n35711) );
  NAND2_X0P5A_A12TR u3677 ( .A(opcode[6]), .B(n3292), .Y(n3228) );
  NAND4B_X0P5M_A12TR u3678 ( .AN(n3975), .B(n4269), .C(n3988), .D(n2868), .Y(
        n4290) );
  NOR2_X0P5A_A12TR u3679 ( .A(n3371), .B(n3383), .Y(n3988) );
  AOI21_X0P5M_A12TR u3680 ( .A0(n3042), .A1(n3200), .B0(n3316), .Y(n3383) );
  OAI21_X0P5M_A12TR u3681 ( .A0(n4293), .A1(n3316), .B0(n3394), .Y(n3371) );
  NAND2_X0P5A_A12TR u3682 ( .A(n3196), .B(n3125), .Y(n3394) );
  INV_X0P5B_A12TR u3683 ( .A(n3389), .Y(n4269) );
  OAI21_X0P5M_A12TR u3684 ( .A0(n3384), .A1(n3038), .B0(n3992), .Y(n3389) );
  NAND2_X0P5A_A12TR u3685 ( .A(n3991), .B(n2983), .Y(n3992) );
  NAND3B_X0P5M_A12TR u3686 ( .AN(n3994), .B(n3993), .C(n4294), .Y(n3975) );
  AOI211_X0P5M_A12TR u3687 ( .A0(n3991), .A1(n3290), .B0(n2865), .C0(n3037), 
        .Y(n4294) );
  INV_X0P5B_A12TR u3688 ( .A(n3641), .Y(n2865) );
  NAND2_X0P5A_A12TR u3689 ( .A(n2825), .B(n3766), .Y(n3641) );
  NOR2_X0P5A_A12TR u3690 ( .A(n3384), .B(n2828), .Y(n3991) );
  AOI211_X0P5M_A12TR u3691 ( .A0(n2825), .A1(n2983), .B0(n2982), .C0(n2981), 
        .Y(n3993) );
  NAND2_X0P5A_A12TR u3692 ( .A(n4295), .B(n4296), .Y(n2981) );
  AOI21_X0P5M_A12TR u3693 ( .A0(n3197), .A1(n3921), .B0(n3426), .Y(n2982) );
  NAND2_X0P5A_A12TR u3694 ( .A(n3204), .B(n236), .Y(n3197) );
  NAND4_X0P5A_A12TR u3695 ( .A(n2861), .B(n4297), .C(n4298), .D(n3655), .Y(
        n3994) );
  NAND2_X0P5A_A12TR u3696 ( .A(n3196), .B(n2825), .Y(n3655) );
  INV_X0P5B_A12TR u3697 ( .A(n3426), .Y(n2825) );
  NAND2_X0P5A_A12TR u3698 ( .A(n235), .B(n3041), .Y(n3426) );
  OAI31_X0P5M_A12TR u3699 ( .A0(n3289), .A1(n3204), .A2(n2828), .B0(n3040), 
        .Y(n4298) );
  INV_X0P5B_A12TR u3700 ( .A(n3567), .Y(n3040) );
  NAND2_X0P5A_A12TR u3701 ( .A(n3189), .B(n3286), .Y(n4297) );
  AOI21_X0P5M_A12TR u3702 ( .A0(n3366), .A1(n4233), .B0(n4299), .Y(n4288) );
  AOI31_X0P5M_A12TR u3703 ( .A0(n2867), .A1(n4307), .A2(n3982), .B0(n2900), 
        .Y(n4299) );
  NAND2_X0P5A_A12TR u3704 ( .A(n3366), .B(n2823), .Y(n2900) );
  AND4_X0P5M_A12TR u3705 ( .A(n4300), .B(n4051), .C(n3567), .D(n4301), .Y(
        n3982) );
  AND4_X0P5M_A12TR u3706 ( .A(n3316), .B(n3384), .C(n2831), .D(n3857), .Y(
        n4301) );
  INV_X0P5B_A12TR u3707 ( .A(n3125), .Y(n3384) );
  NOR2_X0P5A_A12TR u3708 ( .A(n3190), .B(n235), .Y(n3125) );
  NAND3_X0P5A_A12TR u3709 ( .A(n233), .B(n2828), .C(n4302), .Y(n3316) );
  NAND2_X0P5A_A12TR u3710 ( .A(n4302), .B(n3286), .Y(n3567) );
  AOI21B_X0P5M_A12TR u3711 ( .A0(n3037), .A1(n237), .B0N(n2861), .Y(n4300) );
  NOR2B_X0P5M_A12TR u3712 ( .AN(n3330), .B(n3321), .Y(n2861) );
  NOR2_X0P5A_A12TR u3713 ( .A(n3200), .B(n3857), .Y(n3321) );
  NAND2_X0P5A_A12TR u3714 ( .A(n2984), .B(n3039), .Y(n3330) );
  INV_X0P5B_A12TR u3715 ( .A(n3038), .Y(n2984) );
  NAND2_X0P5A_A12TR u3716 ( .A(n2983), .B(n2828), .Y(n3038) );
  INV_X0P5B_A12TR u3717 ( .A(r1298_carry_1_), .Y(n4307) );
  OAI21_X0P5M_A12TR u3718 ( .A0(u3_u93_z_6), .A1(n2869), .B0(n4228), .Y(n4233)
         );
  NAND2_X0P5A_A12TR u3719 ( .A(n3353), .B(n4303), .Y(n4228) );
  INV_X0P5B_A12TR u3720 ( .A(n3042), .Y(n3353) );
  AOI222_X0P5M_A12TR u3721 ( .A0(n2823), .A1(n3977), .B0(n4234), .B1(n3366), 
        .C0(n2826), .C1(n3570), .Y(n2820) );
  INV_X0P5B_A12TR u3722 ( .A(n3642), .Y(n2826) );
  OAI21_X0P5M_A12TR u3723 ( .A0(u3_u93_z_6), .A1(n2868), .B0(n4229), .Y(n4234)
         );
  NAND2_X0P5A_A12TR u3724 ( .A(n4303), .B(n3204), .Y(n4229) );
  INV_X0P5B_A12TR u3725 ( .A(n4227), .Y(n4303) );
  NAND2_X0P5A_A12TR u3726 ( .A(n3852), .B(n2823), .Y(n4227) );
  INV_X0P5B_A12TR u3727 ( .A(n3297), .Y(n3977) );
  NAND2_X0P5A_A12TR u3728 ( .A(n3570), .B(n3366), .Y(n3297) );
  INV_X0P5B_A12TR u3729 ( .A(n3193), .Y(n3366) );
  NAND2_X0P5A_A12TR u3730 ( .A(opcode[7]), .B(opcode[6]), .Y(n3193) );
  NOR2_X0P5A_A12TR u3731 ( .A(n3128), .B(n3190), .Y(n3570) );
  NAND2_X0P5A_A12TR u3732 ( .A(n234), .B(n3286), .Y(n3190) );
  INV_X0P5B_A12TR u3733 ( .A(n4274), .Y(n2824) );
  AO21A1AI2_X0P5M_A12TR u3734 ( .A0(n2869), .A1(n2867), .B0(n3642), .C0(n2821), 
        .Y(n4274) );
  INV_X0P5B_A12TR u3735 ( .A(u3_u87_z_0), .Y(n2821) );
  NOR2_X0P5A_A12TR u3736 ( .A(n3203), .B(n3204), .Y(n4293) );
  NAND2_X0P5A_A12TR u3737 ( .A(n3127), .B(n2823), .Y(n3642) );
  INV_X0P5B_A12TR u3738 ( .A(n3036), .Y(n3127) );
  NAND2_X0P5A_A12TR u3739 ( .A(n3292), .B(n3291), .Y(n3036) );
  INV_X0P5B_A12TR u3740 ( .A(opcode[6]), .Y(n3291) );
  INV_X0P5B_A12TR u3741 ( .A(opcode[7]), .Y(n3292) );
  NAND2_X0P5A_A12TR u3742 ( .A(n3037), .B(n3286), .Y(n3191) );
  INV_X0P5B_A12TR u3743 ( .A(n3343), .Y(n3037) );
  NAND2_X0P5A_A12TR u3744 ( .A(n35721), .B(n2828), .Y(n3356) );
  NAND2_X0P5A_A12TR u3745 ( .A(n2920), .B(n35721), .Y(n3568) );
  NOR2_X0P5A_A12TR u3746 ( .A(n3343), .B(n3286), .Y(n35721) );
  NAND2_X0P5A_A12TR u3747 ( .A(n235), .B(n3288), .Y(n3343) );
  INV_X0P5B_A12TR u3748 ( .A(n3921), .Y(n2920) );
  NAND2_X0P5A_A12TR u3749 ( .A(n3203), .B(n236), .Y(n3921) );
  OAI222_X0P5M_A12TR u3750 ( .A0(n4245), .A1(n4051), .B0(n4304), .B1(n3819), 
        .C0(n3884), .C1(n3393), .Y(u3_u80_z_9) );
  INV_X0P5B_A12TR u3751 ( .A(n1176), .Y(n3884) );
  INV_X0P5B_A12TR u3752 ( .A(sp[9]), .Y(n4245) );
  OAI222_X0P5M_A12TR u3753 ( .A0(n4247), .A1(n4051), .B0(n4304), .B1(n2871), 
        .C0(n3882), .C1(n3393), .Y(u3_u80_z_8) );
  INV_X0P5B_A12TR u3754 ( .A(n1175), .Y(n3882) );
  INV_X0P5B_A12TR u3755 ( .A(sp[8]), .Y(n4247) );
  OAI222_X0P5M_A12TR u3756 ( .A0(n4249), .A1(n4051), .B0(n4304), .B1(n2889), 
        .C0(n3594), .C1(n3393), .Y(u3_u80_z_7) );
  INV_X0P5B_A12TR u3757 ( .A(n1174), .Y(n3594) );
  INV_X0P5B_A12TR u3758 ( .A(sp[7]), .Y(n4249) );
  OAI222_X0P5M_A12TR u3759 ( .A0(n4251), .A1(n4051), .B0(n4304), .B1(n3481), 
        .C0(n3876), .C1(n3393), .Y(u3_u80_z_6) );
  INV_X0P5B_A12TR u3760 ( .A(n1173), .Y(n3876) );
  INV_X0P5B_A12TR u3761 ( .A(sp[6]), .Y(n4251) );
  OAI222_X0P5M_A12TR u3762 ( .A0(n4253), .A1(n4051), .B0(n4304), .B1(n3466), 
        .C0(n3873), .C1(n3393), .Y(u3_u80_z_5) );
  INV_X0P5B_A12TR u3763 ( .A(n1172), .Y(n3873) );
  INV_X0P5B_A12TR u3764 ( .A(sp[5]), .Y(n4253) );
  OAI222_X0P5M_A12TR u3765 ( .A0(n4256), .A1(n4051), .B0(n4304), .B1(n3458), 
        .C0(n3870), .C1(n3393), .Y(u3_u80_z_4) );
  INV_X0P5B_A12TR u3766 ( .A(n1171), .Y(n3870) );
  INV_X0P5B_A12TR u3767 ( .A(sp[4]), .Y(n4256) );
  OAI222_X0P5M_A12TR u3768 ( .A0(n4258), .A1(n4051), .B0(n4304), .B1(n3443), 
        .C0(n3867), .C1(n3393), .Y(u3_u80_z_3) );
  INV_X0P5B_A12TR u3769 ( .A(n1170), .Y(n3867) );
  INV_X0P5B_A12TR u3770 ( .A(sp[3]), .Y(n4258) );
  OAI222_X0P5M_A12TR u3771 ( .A0(n4260), .A1(n4051), .B0(n4304), .B1(n3434), 
        .C0(n3864), .C1(n3393), .Y(u3_u80_z_2) );
  INV_X0P5B_A12TR u3772 ( .A(n1169), .Y(n3864) );
  INV_X0P5B_A12TR u3773 ( .A(sp[2]), .Y(n4260) );
  OAI222_X0P5M_A12TR u3774 ( .A0(n4261), .A1(n4051), .B0(n4304), .B1(n2960), 
        .C0(n2925), .C1(n3393), .Y(u3_u80_z_15) );
  INV_X0P5B_A12TR u3775 ( .A(n1182), .Y(n2925) );
  INV_X0P5B_A12TR u3776 ( .A(sp[15]), .Y(n4261) );
  OAI222_X0P5M_A12TR u3777 ( .A0(n4262), .A1(n4051), .B0(n4304), .B1(n3849), 
        .C0(n3894), .C1(n3393), .Y(u3_u80_z_14) );
  INV_X0P5B_A12TR u3778 ( .A(n1181), .Y(n3894) );
  INV_X0P5B_A12TR u3779 ( .A(sp[14]), .Y(n4262) );
  OAI222_X0P5M_A12TR u3780 ( .A0(n4263), .A1(n4051), .B0(n4304), .B1(n3843), 
        .C0(n3892), .C1(n3393), .Y(u3_u80_z_13) );
  INV_X0P5B_A12TR u3781 ( .A(n1180), .Y(n3892) );
  INV_X0P5B_A12TR u3782 ( .A(sp[13]), .Y(n4263) );
  OAI222_X0P5M_A12TR u3783 ( .A0(n4264), .A1(n4051), .B0(n4304), .B1(n3837), 
        .C0(n3890), .C1(n3393), .Y(u3_u80_z_12) );
  INV_X0P5B_A12TR u3784 ( .A(n1179), .Y(n3890) );
  INV_X0P5B_A12TR u3785 ( .A(sp[12]), .Y(n4264) );
  OAI222_X0P5M_A12TR u3786 ( .A0(n4265), .A1(n4051), .B0(n4304), .B1(n3831), 
        .C0(n3888), .C1(n3393), .Y(u3_u80_z_11) );
  INV_X0P5B_A12TR u3787 ( .A(n1178), .Y(n3888) );
  INV_X0P5B_A12TR u3788 ( .A(sp[11]), .Y(n4265) );
  OAI222_X0P5M_A12TR u3789 ( .A0(n4266), .A1(n4051), .B0(n4304), .B1(n3825), 
        .C0(n3886), .C1(n3393), .Y(u3_u80_z_10) );
  INV_X0P5B_A12TR u3790 ( .A(n1177), .Y(n3886) );
  INV_X0P5B_A12TR u3791 ( .A(sp[10]), .Y(n4266) );
  OAI222_X0P5M_A12TR u3792 ( .A0(n4078), .A1(n4051), .B0(n4304), .B1(n3420), 
        .C0(n3861), .C1(n3393), .Y(u3_u80_z_1) );
  INV_X0P5B_A12TR u3793 ( .A(n1168), .Y(n3861) );
  INV_X0P5B_A12TR u3794 ( .A(sp[1]), .Y(n4078) );
  OAI222_X0P5M_A12TR u3795 ( .A0(n4268), .A1(n4051), .B0(n4304), .B1(n3409), 
        .C0(n3858), .C1(n3393), .Y(u3_u80_z_0) );
  INV_X0P5B_A12TR u3796 ( .A(n1167), .Y(n3858) );
  OA21_X0P5M_A12TR u3797 ( .A0(n3286), .A1(n3969), .B0(n4296), .Y(n4304) );
  INV_X0P5B_A12TR u3798 ( .A(n31370), .Y(n4268) );
  OAI22_X0P5M_A12TR u3799 ( .A0(n4295), .A1(n3819), .B0(n2833), .B1(n4296), 
        .Y(u3_u79_z_9) );
  AOI222_X0P5M_A12TR u3800 ( .A0(n3771), .A1(n1159), .B0(n4305), .B1(
        regfil_2__1_), .C0(n3899), .C1(n1176), .Y(n2833) );
  INV_X0P5B_A12TR u3801 ( .A(n1159), .Y(n3819) );
  OAI22_X0P5M_A12TR u3802 ( .A0(n4295), .A1(n2871), .B0(n4246), .B1(n4296), 
        .Y(u3_u79_z_8) );
  AOI222_X0P5M_A12TR u3803 ( .A0(n3771), .A1(n1158), .B0(n4305), .B1(
        regfil_2__0_), .C0(n3899), .C1(n1175), .Y(n4246) );
  INV_X0P5B_A12TR u3804 ( .A(n1158), .Y(n2871) );
  OAI22_X0P5M_A12TR u3805 ( .A0(n4295), .A1(n2889), .B0(n4248), .B1(n4296), 
        .Y(u3_u79_z_7) );
  AOI222_X0P5M_A12TR u3806 ( .A0(n3771), .A1(n1157), .B0(n4305), .B1(n1664), 
        .C0(n3899), .C1(n1174), .Y(n4248) );
  INV_X0P5B_A12TR u3807 ( .A(n1157), .Y(n2889) );
  OAI22_X0P5M_A12TR u3808 ( .A0(n4295), .A1(n3481), .B0(n4250), .B1(n4296), 
        .Y(u3_u79_z_6) );
  AOI222_X0P5M_A12TR u3809 ( .A0(n3771), .A1(n1156), .B0(n4305), .B1(n1663), 
        .C0(n3899), .C1(n1173), .Y(n4250) );
  INV_X0P5B_A12TR u3810 ( .A(n1156), .Y(n3481) );
  OAI22_X0P5M_A12TR u3811 ( .A0(n4295), .A1(n3466), .B0(n4252), .B1(n4296), 
        .Y(u3_u79_z_5) );
  AOI222_X0P5M_A12TR u3812 ( .A0(n3771), .A1(n1155), .B0(n4305), .B1(n1662), 
        .C0(n3899), .C1(n1172), .Y(n4252) );
  INV_X0P5B_A12TR u3813 ( .A(n1155), .Y(n3466) );
  OAI22_X0P5M_A12TR u3814 ( .A0(n4295), .A1(n3458), .B0(n4254), .B1(n4296), 
        .Y(u3_u79_z_4) );
  AOI222_X0P5M_A12TR u3815 ( .A0(n3771), .A1(n1154), .B0(n4305), .B1(n1661), 
        .C0(n3899), .C1(n1171), .Y(n4254) );
  INV_X0P5B_A12TR u3816 ( .A(n1154), .Y(n3458) );
  OAI22_X0P5M_A12TR u3817 ( .A0(n4295), .A1(n3443), .B0(n4257), .B1(n4296), 
        .Y(u3_u79_z_3) );
  AOI222_X0P5M_A12TR u3818 ( .A0(n3771), .A1(n1153), .B0(n4305), .B1(n1660), 
        .C0(n3899), .C1(n1170), .Y(n4257) );
  INV_X0P5B_A12TR u3819 ( .A(n1153), .Y(n3443) );
  OAI22_X0P5M_A12TR u3820 ( .A0(n4295), .A1(n3434), .B0(n4259), .B1(n4296), 
        .Y(u3_u79_z_2) );
  AOI222_X0P5M_A12TR u3821 ( .A0(n3771), .A1(n1152), .B0(n4305), .B1(n1659), 
        .C0(n3899), .C1(n1169), .Y(n4259) );
  INV_X0P5B_A12TR u3822 ( .A(n1152), .Y(n3434) );
  OAI22_X0P5M_A12TR u3823 ( .A0(n4295), .A1(n2960), .B0(n2836), .B1(n4296), 
        .Y(u3_u79_z_15) );
  AOI222_X0P5M_A12TR u3824 ( .A0(n3771), .A1(n1165), .B0(n4305), .B1(
        regfil_2__7_), .C0(n3899), .C1(n1182), .Y(n2836) );
  INV_X0P5B_A12TR u3825 ( .A(n1165), .Y(n2960) );
  OAI22_X0P5M_A12TR u3826 ( .A0(n4295), .A1(n3849), .B0(n2839), .B1(n4296), 
        .Y(u3_u79_z_14) );
  AOI222_X0P5M_A12TR u3827 ( .A0(n3771), .A1(n1164), .B0(n4305), .B1(
        regfil_2__6_), .C0(n3899), .C1(n1181), .Y(n2839) );
  INV_X0P5B_A12TR u3828 ( .A(n1164), .Y(n3849) );
  OAI22_X0P5M_A12TR u3829 ( .A0(n4295), .A1(n3843), .B0(n2842), .B1(n4296), 
        .Y(u3_u79_z_13) );
  AOI222_X0P5M_A12TR u3830 ( .A0(n3771), .A1(n1163), .B0(n4305), .B1(
        regfil_2__5_), .C0(n3899), .C1(n1180), .Y(n2842) );
  INV_X0P5B_A12TR u3831 ( .A(n1163), .Y(n3843) );
  OAI22_X0P5M_A12TR u3832 ( .A0(n4295), .A1(n3837), .B0(n2845), .B1(n4296), 
        .Y(u3_u79_z_12) );
  AOI222_X0P5M_A12TR u3833 ( .A0(n3771), .A1(n1162), .B0(n4305), .B1(
        regfil_2__4_), .C0(n3899), .C1(n1179), .Y(n2845) );
  INV_X0P5B_A12TR u3834 ( .A(n1162), .Y(n3837) );
  OAI22_X0P5M_A12TR u3835 ( .A0(n4295), .A1(n3831), .B0(n2848), .B1(n4296), 
        .Y(u3_u79_z_11) );
  AOI222_X0P5M_A12TR u3836 ( .A0(n3771), .A1(n1161), .B0(n4305), .B1(
        regfil_2__3_), .C0(n3899), .C1(n1178), .Y(n2848) );
  INV_X0P5B_A12TR u3837 ( .A(n1161), .Y(n3831) );
  OAI22_X0P5M_A12TR u3838 ( .A0(n4295), .A1(n3825), .B0(n2851), .B1(n4296), 
        .Y(u3_u79_z_10) );
  AOI222_X0P5M_A12TR u3839 ( .A0(n3771), .A1(n1160), .B0(n4305), .B1(
        regfil_2__2_), .C0(n3899), .C1(n1177), .Y(n2851) );
  INV_X0P5B_A12TR u3840 ( .A(n1160), .Y(n3825) );
  OAI22_X0P5M_A12TR u3841 ( .A0(n4295), .A1(n3420), .B0(n4267), .B1(n4296), 
        .Y(u3_u79_z_1) );
  AOI222_X0P5M_A12TR u3842 ( .A0(n3771), .A1(n1151), .B0(n4305), .B1(n1658), 
        .C0(n3899), .C1(n1168), .Y(n4267) );
  INV_X0P5B_A12TR u3843 ( .A(n1151), .Y(n3420) );
  OAI22_X0P5M_A12TR u3844 ( .A0(n2854), .A1(n4296), .B0(n4295), .B1(n3409), 
        .Y(u3_u79_z_0) );
  INV_X0P5B_A12TR u3845 ( .A(n1150), .Y(n3409) );
  OA211_X0P5M_A12TR u3846 ( .A0(n3286), .A1(n3969), .B0(n4051), .C0(n3393), 
        .Y(n4295) );
  NAND2_X0P5A_A12TR u3847 ( .A(n4306), .B(n3203), .Y(n3393) );
  INV_X0P5B_A12TR u3848 ( .A(n2829), .Y(n3203) );
  NAND2_X0P5A_A12TR u3849 ( .A(n2983), .B(n4306), .Y(n4051) );
  INV_X0P5B_A12TR u3850 ( .A(n3200), .Y(n2983) );
  NAND2_X0P5A_A12TR u3851 ( .A(n46), .B(n237), .Y(n3200) );
  NAND2_X0P5A_A12TR u3852 ( .A(n3196), .B(n4302), .Y(n3969) );
  NOR2_X0P5A_A12TR u3853 ( .A(n3042), .B(n2828), .Y(n3196) );
  INV_X0P5B_A12TR u3854 ( .A(n236), .Y(n2828) );
  AOI222_X0P5M_A12TR u3855 ( .A0(n3771), .A1(n1150), .B0(n4305), .B1(n1657), 
        .C0(n3899), .C1(n1167), .Y(n2854) );
  OAI21_X0P5M_A12TR u3856 ( .A0(n3857), .A1(n2829), .B0(n2867), .Y(n3899) );
  NAND3_X0P5A_A12TR u3857 ( .A(n3041), .B(n3289), .C(n3189), .Y(n2867) );
  NAND2_X0P5A_A12TR u3858 ( .A(n3289), .B(n3290), .Y(n2829) );
  NAND2_X0P5A_A12TR u3859 ( .A(n3375), .B(n4296), .Y(n4305) );
  NAND2_X0P5A_A12TR u3860 ( .A(n4306), .B(n3204), .Y(n4296) );
  AND3_X0P5M_A12TR u3861 ( .A(n236), .B(n233), .C(n4302), .Y(n4306) );
  NOR2_X0P5A_A12TR u3862 ( .A(n235), .B(n234), .Y(n4302) );
  AOI21_X0P5M_A12TR u3863 ( .A0(n3852), .A1(n3204), .B0(n3350), .Y(n3375) );
  INV_X0P5B_A12TR u3864 ( .A(n2868), .Y(n3350) );
  NAND3_X0P5A_A12TR u3865 ( .A(n46), .B(n3041), .C(n3189), .Y(n2868) );
  INV_X0P5B_A12TR u3866 ( .A(n3129), .Y(n3189) );
  NAND2_X0P5A_A12TR u3867 ( .A(n3990), .B(n3128), .Y(n3129) );
  INV_X0P5B_A12TR u3868 ( .A(n235), .Y(n3128) );
  NOR2_X0P5A_A12TR u3869 ( .A(n236), .B(n237), .Y(n3990) );
  INV_X0P5B_A12TR u3870 ( .A(n2831), .Y(n3204) );
  NAND2_X0P5A_A12TR u3871 ( .A(n46), .B(n3290), .Y(n2831) );
  INV_X0P5B_A12TR u3872 ( .A(n237), .Y(n3290) );
  INV_X0P5B_A12TR u3873 ( .A(n3857), .Y(n3852) );
  OAI21_X0P5M_A12TR u3874 ( .A0(n3857), .A1(n3042), .B0(n2869), .Y(n3771) );
  NAND2_X0P5A_A12TR u3875 ( .A(n3766), .B(n3039), .Y(n2869) );
  NOR2_X0P5A_A12TR u3876 ( .A(n3042), .B(n236), .Y(n3766) );
  NAND2_X0P5A_A12TR u3877 ( .A(n237), .B(n3289), .Y(n3042) );
  INV_X0P5B_A12TR u3878 ( .A(n46), .Y(n3289) );
  NAND2_X0P5A_A12TR u3879 ( .A(n236), .B(n3039), .Y(n3857) );
  NOR2B_X0P5M_A12TR u3880 ( .AN(n3041), .B(n235), .Y(n3039) );
  NOR2_X0P5A_A12TR u3881 ( .A(n3288), .B(n3286), .Y(n3041) );
  INV_X0P5B_A12TR u3882 ( .A(n233), .Y(n3286) );
  INV_X0P5B_A12TR u3883 ( .A(n234), .Y(n3288) );
  INV_X0P5B_A12TR alu_u87 ( .A(aluopra[7]), .Y(alu_n20) );
  INV_X0P5B_A12TR alu_u86 ( .A(n4311), .Y(alu_n42) );
  NOR2_X0P5A_A12TR alu_u85 ( .A(alu_n20), .B(alu_n42), .Y(alu_n101) );
  INV_X0P5B_A12TR alu_u84 ( .A(aluopra[6]), .Y(alu_n22) );
  INV_X0P5B_A12TR alu_u83 ( .A(n4308), .Y(alu_n41) );
  NOR2_X0P5A_A12TR alu_u82 ( .A(alu_n22), .B(alu_n41), .Y(alu_n110) );
  INV_X0P5B_A12TR alu_u81 ( .A(aluopra[5]), .Y(alu_n23) );
  INV_X0P5B_A12TR alu_u80 ( .A(n4313), .Y(alu_n40) );
  NOR2_X0P5A_A12TR alu_u79 ( .A(alu_n23), .B(alu_n40), .Y(alu_n120) );
  INV_X0P5B_A12TR alu_u78 ( .A(aluopra[4]), .Y(alu_n24) );
  INV_X0P5B_A12TR alu_u77 ( .A(n4309), .Y(alu_n39) );
  NOR2_X0P5A_A12TR alu_u76 ( .A(alu_n24), .B(alu_n39), .Y(alu_n130) );
  INV_X0P5B_A12TR alu_u75 ( .A(aluopra[3]), .Y(alu_n25) );
  INV_X0P5B_A12TR alu_u74 ( .A(n4314), .Y(alu_n38) );
  NOR2_X0P5A_A12TR alu_u73 ( .A(alu_n25), .B(alu_n38), .Y(alu_n140) );
  INV_X0P5B_A12TR alu_u72 ( .A(aluopra[2]), .Y(alu_n26) );
  INV_X0P5B_A12TR alu_u71 ( .A(n4315), .Y(alu_n37) );
  NOR2_X0P5A_A12TR alu_u70 ( .A(alu_n26), .B(alu_n37), .Y(alu_n150) );
  INV_X0P5B_A12TR alu_u69 ( .A(aluopra[1]), .Y(alu_n27) );
  INV_X0P5B_A12TR alu_u68 ( .A(n4316), .Y(alu_n35) );
  NOR2_X0P5A_A12TR alu_u67 ( .A(alu_n27), .B(alu_n35), .Y(alu_n160) );
  INV_X0P5B_A12TR alu_u66 ( .A(aluopra[0]), .Y(alu_n28) );
  INV_X0P5B_A12TR alu_u65 ( .A(aluoprb_0_), .Y(alu_n34) );
  NOR2_X0P5A_A12TR alu_u64 ( .A(alu_n28), .B(alu_n34), .Y(alu_n170) );
  XNOR2_X0P5M_A12TR alu_u63 ( .A(alu_n42), .B(aluopra[7]), .Y(alu_n180) );
  XNOR2_X0P5M_A12TR alu_u62 ( .A(alu_n41), .B(aluopra[6]), .Y(alu_n190) );
  XNOR2_X0P5M_A12TR alu_u61 ( .A(alu_n40), .B(aluopra[5]), .Y(alu_n200) );
  XNOR2_X0P5M_A12TR alu_u60 ( .A(alu_n39), .B(aluopra[4]), .Y(alu_n210) );
  XNOR2_X0P5M_A12TR alu_u59 ( .A(alu_n38), .B(aluopra[3]), .Y(alu_n220) );
  XNOR2_X0P5M_A12TR alu_u58 ( .A(alu_n37), .B(aluopra[2]), .Y(alu_n230) );
  XNOR2_X0P5M_A12TR alu_u57 ( .A(alu_n35), .B(aluopra[1]), .Y(alu_n240) );
  XNOR2_X0P5M_A12TR alu_u56 ( .A(alu_n34), .B(aluopra[0]), .Y(alu_n250) );
  NAND2_X0P5A_A12TR alu_u55 ( .A(alu_n42), .B(alu_n20), .Y(alu_n260) );
  NAND2_X0P5A_A12TR alu_u54 ( .A(alu_n41), .B(alu_n22), .Y(alu_n270) );
  NAND2_X0P5A_A12TR alu_u53 ( .A(alu_n40), .B(alu_n23), .Y(alu_n280) );
  NAND2_X0P5A_A12TR alu_u52 ( .A(alu_n39), .B(alu_n24), .Y(alu_n290) );
  NAND2_X0P5A_A12TR alu_u51 ( .A(alu_n38), .B(alu_n25), .Y(alu_n300) );
  NAND2_X0P5A_A12TR alu_u50 ( .A(alu_n37), .B(alu_n26), .Y(alu_n310) );
  NAND2_X0P5A_A12TR alu_u49 ( .A(alu_n35), .B(alu_n27), .Y(alu_n320) );
  NAND2_X0P5A_A12TR alu_u48 ( .A(alu_n34), .B(alu_n28), .Y(alu_n330) );
  INV_X0P5B_A12TR alu_u47 ( .A(alusel[2]), .Y(alu_n33) );
  AND3_X0P5M_A12TR alu_u46 ( .A(alusel[0]), .B(alu_n33), .C(alucin), .Y(
        alu_u2_u3_z_0) );
  NAND3_X0P5A_A12TR alu_u45 ( .A(alusel[1]), .B(alusel[0]), .C(alusel[2]), .Y(
        alu_n21) );
  AO1B2_X0P5M_A12TR alu_u44 ( .B0(alu_n33), .B1(alusel[1]), .A0N(alu_n21), .Y(
        alu_u2_u4_z_0) );
  XNOR2_X0P5M_A12TR alu_u43 ( .A(alu_n1), .B(alu_resi_2_), .Y(alu_n32) );
  XNOR3_X0P5M_A12TR alu_u42 ( .A(alu_n32), .B(alu_resi_1_), .C(alu_resi_0_), 
        .Y(alu_n29) );
  INV_X0P5B_A12TR alu_u41 ( .A(alusout), .Y(alu_n19) );
  XNOR2_X0P5M_A12TR alu_u40 ( .A(alu_n19), .B(alu_resi_6_), .Y(alu_n31) );
  XNOR3_X0P5M_A12TR alu_u39 ( .A(alu_n2), .B(alu_n31), .C(alu_resi_4_), .Y(
        alu_n30) );
  XOR2_X0P5M_A12TR alu_u38 ( .A(alu_n29), .B(alu_n30), .Y(alupar) );
  INV_X0P5B_A12TR alu_u37 ( .A(alu_resi_0_), .Y(alu_n14) );
  MXIT2_X0P5M_A12TR alu_u36 ( .A(alu_n28), .B(alu_n14), .S0(alu_n21), .Y(
        alures[0]) );
  INV_X0P5B_A12TR alu_u35 ( .A(alu_resi_1_), .Y(alu_n15) );
  MXIT2_X0P5M_A12TR alu_u34 ( .A(alu_n27), .B(alu_n15), .S0(alu_n21), .Y(
        alures[1]) );
  INV_X0P5B_A12TR alu_u33 ( .A(alu_resi_2_), .Y(alu_n16) );
  MXIT2_X0P5M_A12TR alu_u32 ( .A(alu_n26), .B(alu_n16), .S0(alu_n21), .Y(
        alures[2]) );
  MXIT2_X0P5M_A12TR alu_u31 ( .A(alu_n25), .B(alu_n1), .S0(alu_n21), .Y(
        alures[3]) );
  INV_X0P5B_A12TR alu_u30 ( .A(alu_resi_4_), .Y(alu_n17) );
  MXIT2_X0P5M_A12TR alu_u29 ( .A(alu_n24), .B(alu_n17), .S0(alu_n21), .Y(
        alures[4]) );
  MXIT2_X0P5M_A12TR alu_u28 ( .A(alu_n23), .B(alu_n2), .S0(alu_n21), .Y(
        alures[5]) );
  INV_X0P5B_A12TR alu_u27 ( .A(alu_resi_6_), .Y(alu_n18) );
  MXIT2_X0P5M_A12TR alu_u26 ( .A(alu_n22), .B(alu_n18), .S0(alu_n21), .Y(
        alures[6]) );
  MXIT2_X0P5M_A12TR alu_u25 ( .A(alu_n20), .B(alu_n19), .S0(alu_n21), .Y(
        alures[7]) );
  NAND4_X0P5A_A12TR alu_u24 ( .A(alu_n17), .B(alu_n2), .C(alu_n18), .D(alu_n19), .Y(alu_n12) );
  NAND4_X0P5A_A12TR alu_u23 ( .A(alu_n14), .B(alu_n15), .C(alu_n16), .D(alu_n1), .Y(alu_n13) );
  NOR2_X0P5A_A12TR alu_u22 ( .A(alu_n12), .B(alu_n13), .Y(aluzout) );
  TIELO_X1M_A12TR alu_u21 ( .Y(alu_n36) );
  NOR2XB_X1M_A12TR alu_u20 ( .BN(alu_n100), .A(alu_n3), .Y(aluaxc) );
  MXT4_X1M_A12TR alu_u19 ( .A(alu_n170), .B(alu_n330), .C(alu_n250), .D(
        alu_n91), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n11) );
  MXT2_X1M_A12TR alu_u18 ( .A(alu_n91), .B(alu_n11), .S0(alusel[2]), .Y(
        alu_resi_0_) );
  MXT4_X1M_A12TR alu_u17 ( .A(alu_n130), .B(alu_n290), .C(alu_n210), .D(
        alu_n95), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n10) );
  MXT2_X1M_A12TR alu_u16 ( .A(alu_n95), .B(alu_n10), .S0(alusel[2]), .Y(
        alu_resi_4_) );
  MXT4_X1M_A12TR alu_u15 ( .A(alu_n101), .B(alu_n260), .C(alu_n180), .D(
        alu_n98), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n9) );
  MXT2_X1M_A12TR alu_u14 ( .A(alu_n98), .B(alu_n9), .S0(alusel[2]), .Y(alusout) );
  MXT4_X1M_A12TR alu_u13 ( .A(alu_n110), .B(alu_n270), .C(alu_n190), .D(
        alu_n97), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n8) );
  MXT2_X1M_A12TR alu_u12 ( .A(alu_n97), .B(alu_n8), .S0(alusel[2]), .Y(
        alu_resi_6_) );
  MXT4_X1M_A12TR alu_u11 ( .A(alu_n150), .B(alu_n310), .C(alu_n230), .D(
        alu_n93), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n7) );
  MXT2_X1M_A12TR alu_u10 ( .A(alu_n93), .B(alu_n7), .S0(alusel[2]), .Y(
        alu_resi_2_) );
  MXT4_X1M_A12TR alu_u9 ( .A(alu_n160), .B(alu_n320), .C(alu_n240), .D(alu_n92), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n6) );
  MXT2_X1M_A12TR alu_u8 ( .A(alu_n92), .B(alu_n6), .S0(alusel[2]), .Y(
        alu_resi_1_) );
  MXT4_X1M_A12TR alu_u7 ( .A(alu_n120), .B(alu_n280), .C(alu_n200), .D(alu_n96), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n5) );
  MXT4_X1M_A12TR alu_u6 ( .A(alu_n140), .B(alu_n300), .C(alu_n220), .D(alu_n94), .S0(alusel[1]), .S1(alusel[0]), .Y(alu_n4) );
  AOI21B_X1M_A12TR alu_u5 ( .A0(alusel[0]), .A1(alusel[1]), .B0N(alusel[2]), 
        .Y(alu_n3) );
  NOR2XB_X1M_A12TR alu_u4 ( .BN(alu_n99), .A(alu_n3), .Y(alucout) );
  MXIT2_X0P7M_A12TR alu_u3 ( .A(alu_n96), .B(alu_n5), .S0(alusel[2]), .Y(
        alu_n2) );
  MXIT2_X0P7M_A12TR alu_u2 ( .A(alu_n94), .B(alu_n4), .S0(alusel[2]), .Y(
        alu_n1) );
  XOR2_X0P5M_A12TR alu_r24_u10 ( .A(aluoprb_0_), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_0_) );
  XOR2_X0P5M_A12TR alu_r24_u9 ( .A(n4316), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_1_) );
  XOR2_X0P5M_A12TR alu_r24_u8 ( .A(n4315), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_2_) );
  XOR2_X0P5M_A12TR alu_r24_u7 ( .A(n4314), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_3_) );
  XOR2_X0P5M_A12TR alu_r24_u6 ( .A(n4309), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_4_) );
  XOR2_X0P5M_A12TR alu_r24_u5 ( .A(n4313), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_5_) );
  XOR2_X0P5M_A12TR alu_r24_u4 ( .A(n4308), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_6_) );
  XOR2_X0P5M_A12TR alu_r24_u3 ( .A(n4311), .B(alu_u2_u4_z_0), .Y(
        alu_r24_b_as_7_) );
  XOR2_X0P5M_A12TR alu_r24_u2 ( .A(alu_u2_u3_z_0), .B(alu_u2_u4_z_0), .Y(
        alu_r24_carry[0]) );
  XOR2_X1M_A12TR alu_r24_u1 ( .A(alu_u2_u4_z_0), .B(alu_r24_carry[8]), .Y(
        alu_n99) );
  ADDF_X1M_A12TR alu_r24_u1_0 ( .A(aluopra[0]), .B(alu_r24_b_as_0_), .CI(
        alu_r24_carry[0]), .CO(alu_r24_carry[1]), .S(alu_n91) );
  ADDF_X1M_A12TR alu_r24_u1_1 ( .A(aluopra[1]), .B(alu_r24_b_as_1_), .CI(
        alu_r24_carry[1]), .CO(alu_r24_carry[2]), .S(alu_n92) );
  ADDF_X1M_A12TR alu_r24_u1_2 ( .A(aluopra[2]), .B(alu_r24_b_as_2_), .CI(
        alu_r24_carry[2]), .CO(alu_r24_carry[3]), .S(alu_n93) );
  ADDF_X1M_A12TR alu_r24_u1_3 ( .A(aluopra[3]), .B(alu_r24_b_as_3_), .CI(
        alu_r24_carry[3]), .CO(alu_r24_carry[4]), .S(alu_n94) );
  ADDF_X1M_A12TR alu_r24_u1_4 ( .A(aluopra[4]), .B(alu_r24_b_as_4_), .CI(
        alu_r24_carry[4]), .CO(alu_r24_carry[5]), .S(alu_n95) );
  ADDF_X1M_A12TR alu_r24_u1_5 ( .A(aluopra[5]), .B(alu_r24_b_as_5_), .CI(
        alu_r24_carry[5]), .CO(alu_r24_carry[6]), .S(alu_n96) );
  ADDF_X1M_A12TR alu_r24_u1_6 ( .A(aluopra[6]), .B(alu_r24_b_as_6_), .CI(
        alu_r24_carry[6]), .CO(alu_r24_carry[7]), .S(alu_n97) );
  ADDF_X1M_A12TR alu_r24_u1_7 ( .A(aluopra[7]), .B(alu_r24_b_as_7_), .CI(
        alu_r24_carry[7]), .CO(alu_r24_carry[8]), .S(alu_n98) );
  XOR2_X0P5M_A12TR alu_r373_u15 ( .A(aluoprb_0_), .B(alu_u2_u4_z_0), .Y(
        alu_r373_n12) );
  XOR2_X0P5M_A12TR alu_r373_u14 ( .A(alu_u2_u3_z_0), .B(alu_u2_u4_z_0), .Y(
        alu_r373_n13) );
  CGENI_X1M_A12TR alu_r373_u13 ( .A(aluopra[0]), .B(alu_r373_n12), .CI(
        alu_r373_n13), .CON(alu_r373_n9) );
  NOR2B_X0P5M_A12TR alu_r373_u12 ( .AN(alu_r373_n9), .B(aluopra[1]), .Y(
        alu_r373_n10) );
  XNOR2_X0P5M_A12TR alu_r373_u11 ( .A(alu_u2_u4_z_0), .B(n4316), .Y(
        alu_r373_n11) );
  OAI22_X0P5M_A12TR alu_r373_u10 ( .A0(alu_r373_n9), .A1(alu_r373_n2), .B0(
        alu_r373_n10), .B1(alu_r373_n11), .Y(alu_r373_n6) );
  OR2_X0P5M_A12TR alu_r373_u9 ( .A(aluopra[2]), .B(alu_r373_n6), .Y(
        alu_r373_n7) );
  XOR2_X0P5M_A12TR alu_r373_u8 ( .A(alu_u2_u4_z_0), .B(n4315), .Y(alu_r373_n8)
         );
  AOI22_X0P5M_A12TR alu_r373_u7 ( .A0(alu_r373_n6), .A1(aluopra[2]), .B0(
        alu_r373_n7), .B1(alu_r373_n8), .Y(alu_r373_n3) );
  NOR2B_X0P5M_A12TR alu_r373_u6 ( .AN(alu_r373_n3), .B(aluopra[3]), .Y(
        alu_r373_n4) );
  XNOR2_X0P5M_A12TR alu_r373_u5 ( .A(alu_u2_u4_z_0), .B(n4314), .Y(alu_r373_n5) );
  OAI22_X0P5M_A12TR alu_r373_u4 ( .A0(alu_r373_n3), .A1(alu_r373_n1), .B0(
        alu_r373_n4), .B1(alu_r373_n5), .Y(alu_r373_carry_4_) );
  INV_X1M_A12TR alu_r373_u3 ( .A(aluopra[1]), .Y(alu_r373_n2) );
  INV_X1M_A12TR alu_r373_u2 ( .A(aluopra[3]), .Y(alu_r373_n1) );
  XOR2_X1M_A12TR alu_r373_u1 ( .A(alu_u2_u4_z_0), .B(alu_r373_carry_4_), .Y(
        alu_n100) );
  XOR2_X1M_A12TR r1610_u2 ( .A(u3_u80_z_0), .B(u3_u79_z_0), .Y(n1318) );
  AND2_X1M_A12TR r1610_u1 ( .A(u3_u80_z_0), .B(u3_u79_z_0), .Y(r1610_n1) );
  ADDF_X1M_A12TR r1610_u1_1 ( .A(u3_u79_z_1), .B(u3_u80_z_1), .CI(r1610_n1), 
        .CO(r1610_carry_2_), .S(n1319) );
  ADDF_X1M_A12TR r1610_u1_2 ( .A(u3_u79_z_2), .B(u3_u80_z_2), .CI(
        r1610_carry_2_), .CO(r1610_carry_3_), .S(n1320) );
  ADDF_X1M_A12TR r1610_u1_3 ( .A(u3_u79_z_3), .B(u3_u80_z_3), .CI(
        r1610_carry_3_), .CO(r1610_carry_4_), .S(n1321) );
  ADDF_X1M_A12TR r1610_u1_4 ( .A(u3_u79_z_4), .B(u3_u80_z_4), .CI(
        r1610_carry_4_), .CO(r1610_carry_5_), .S(n1322) );
  ADDF_X1M_A12TR r1610_u1_5 ( .A(u3_u79_z_5), .B(u3_u80_z_5), .CI(
        r1610_carry_5_), .CO(r1610_carry_6_), .S(n1323) );
  ADDF_X1M_A12TR r1610_u1_6 ( .A(u3_u79_z_6), .B(u3_u80_z_6), .CI(
        r1610_carry_6_), .CO(r1610_carry_7_), .S(n1324) );
  ADDF_X1M_A12TR r1610_u1_7 ( .A(u3_u79_z_7), .B(u3_u80_z_7), .CI(
        r1610_carry_7_), .CO(r1610_carry_8_), .S(n1325) );
  ADDF_X1M_A12TR r1610_u1_8 ( .A(u3_u79_z_8), .B(u3_u80_z_8), .CI(
        r1610_carry_8_), .CO(r1610_carry_9_), .S(n1326) );
  ADDF_X1M_A12TR r1610_u1_9 ( .A(u3_u79_z_9), .B(u3_u80_z_9), .CI(
        r1610_carry_9_), .CO(r1610_carry_10_), .S(n1327) );
  ADDF_X1M_A12TR r1610_u1_10 ( .A(u3_u79_z_10), .B(u3_u80_z_10), .CI(
        r1610_carry_10_), .CO(r1610_carry_11_), .S(n1328) );
  ADDF_X1M_A12TR r1610_u1_11 ( .A(u3_u79_z_11), .B(u3_u80_z_11), .CI(
        r1610_carry_11_), .CO(r1610_carry_12_), .S(n1329) );
  ADDF_X1M_A12TR r1610_u1_12 ( .A(u3_u79_z_12), .B(u3_u80_z_12), .CI(
        r1610_carry_12_), .CO(r1610_carry_13_), .S(n1330) );
  ADDF_X1M_A12TR r1610_u1_13 ( .A(u3_u79_z_13), .B(u3_u80_z_13), .CI(
        r1610_carry_13_), .CO(r1610_carry_14_), .S(n1331) );
  ADDF_X1M_A12TR r1610_u1_14 ( .A(u3_u79_z_14), .B(u3_u80_z_14), .CI(
        r1610_carry_14_), .CO(r1610_carry_15_), .S(n1332) );
  ADDF_X1M_A12TR r1610_u1_15 ( .A(u3_u79_z_15), .B(u3_u80_z_15), .CI(
        r1610_carry_15_), .CO(n1334), .S(n1333) );
endmodule

