
module router ( clk, reset, currx, curry, flitin_0, flitin_1, flitout_0, 
        flitout_1, creditin_0, creditin_1, creditout_0, creditout_1, seu );
  input [2:0] currx;
  input [2:0] curry;
  input [11:0] flitin_0;
  input [11:0] flitin_1;
  output [11:0] flitout_0;
  output [11:0] flitout_1;
  input clk, reset, creditin_0, creditin_1, seu;
  output creditout_0, creditout_1;
  wire   tailout_1, s0m_no_bufs0, s0m_no_bufs1, s0m_elig_0_, s0m_elig_1_,
         x0m_n6, x0m_n5, x0m_n4, x0m_n3, c0nm_b0m_rdata_1_, c0nm_r0m_n11,
         c0nm_r0m_n10, c0nm_v0m_n64, c0nm_v0m_n62, c0nm_v0m_n61, c0nm_v0m_n58,
         c0nm_v0m_n57, s0m_m0m_n10, s0m_o0nm_n42, s0m_o0nm_n41, s0m_o0nm_n38,
         s0m_o0nm_n37, s0m_o0nm_n36, s0m_o0nm_n35, s0m_o0nm_state_assigned,
         c0sm_b0m_rdata_1_, s0m_m1m_n10, s0m_o0sm_n42, s0m_o0sm_n41,
         s0m_o0sm_n38, s0m_o0sm_n37, s0m_o0sm_n36, s0m_o0sm_n35,
         s0m_o0sm_state_assigned, c0sm_r0m_n11, c0sm_r0m_n10, c0sm_v0m_n64,
         c0sm_v0m_n62, c0sm_v0m_n61, c0sm_v0m_n58, c0sm_v0m_n57,
         c0nm_b0m_v0m_n171, c0nm_b0m_v0m_head_1_, c0sm_b0m_v0m_n171,
         c0sm_b0m_v0m_head_1_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n66, n67, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n134, n135, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n147, n148, n150, n151, n158, n168, n193, n194, n212, n219,
         n220, n221, n239, n240, n241, n242, n243, n244, n245, n313, n314,
         n315, n316, n317, n318, n319, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n970, n971, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487;

  DFFQ_X1M_A12TR s0m_o0sm_state_assigned_reg ( .D(s0m_o0sm_n35), .CK(clk), .Q(
        s0m_o0sm_state_assigned) );
  DFFQ_X1M_A12TR s0m_o0nm_state_assigned_reg ( .D(s0m_o0nm_n35), .CK(clk), .Q(
        s0m_o0nm_state_assigned) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_1_ ( .D(n903), .CK(clk), .Q(
        c0nm_b0m_rdata_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_1_ ( .D(n839), .CK(clk), .Q(
        c0sm_b0m_rdata_1_) );
  DFFQ_X1M_A12TR c0nm_b0m_dqenablereg_reg ( .D(n168), .CK(clk), .Q(n139) );
  DFFQ_X1M_A12TR s0m_o0nm_eligible_reg ( .D(s0m_o0nm_n41), .CK(clk), .Q(
        s0m_elig_0_) );
  DFFQ_X1M_A12TR s0m_o0sm_eligible_reg ( .D(s0m_o0sm_n41), .CK(clk), .Q(
        s0m_elig_1_) );
  DFFQ_X1M_A12TR s0m_o0nm_no_bufs_reg ( .D(s0m_o0nm_n42), .CK(clk), .Q(
        s0m_no_bufs0) );
  DFFQ_X1M_A12TR s0m_o0sm_no_bufs_reg ( .D(s0m_o0sm_n42), .CK(clk), .Q(
        s0m_no_bufs1) );
  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_1_ ( .D(n959), .CK(clk), .Q(
        c0nm_b0m_v0m_head_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_1_ ( .D(n889), .CK(clk), .Q(
        c0sm_b0m_v0m_head_1_) );
  DFFQ_X1M_A12TR c0sm_b0m_dqenablereg_reg ( .D(n158), .CK(clk), .Q(n71) );
  DFFQ_X1M_A12TR c0sm_b0m_v0m_tailout_reg ( .D(c0sm_b0m_v0m_n171), .CK(clk), 
        .Q(tailout_1) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_tailout_reg ( .D(c0nm_b0m_v0m_n171), .CK(clk), 
        .QN(n124) );
  DFFQN_X1M_A12TR s0m_resp0_reg_0_ ( .D(n905), .CK(clk), .QN(n140) );
  DFFQN_X1M_A12TR s0m_resp0_reg_1_ ( .D(n961), .CK(clk), .QN(n6) );
  DFFQN_X1M_A12TR s0m_o0nm_state_invc_reg_1_ ( .D(n891), .CK(clk), .QN(n143)
         );
  DFFQN_X1M_A12TR s0m_o0sm_state_invc_reg_1_ ( .D(n907), .CK(clk), .QN(n2) );
  DFFQN_X1M_A12TR c0nm_r0m_vc_req_reg_0_ ( .D(c0nm_r0m_n10), .CK(clk), .QN(
        n193) );
  DFFQN_X1M_A12TR c0sm_r0m_vc_req_reg_1_ ( .D(c0sm_r0m_n11), .CK(clk), .QN(
        n221) );
  DFFQN_X1M_A12TR c0nm_v0m_state_queuelen_reg_1_ ( .D(c0nm_v0m_n62), .CK(clk), 
        .QN(n137) );
  DFFQN_X1M_A12TR c0nm_r0m_vc_req_reg_1_ ( .D(c0nm_r0m_n11), .CK(clk), .QN(
        n194) );
  DFFQN_X1M_A12TR c0sm_r0m_vc_req_reg_0_ ( .D(c0sm_r0m_n10), .CK(clk), .QN(
        n220) );
  DFFQN_X1M_A12TR c0nm_v0m_full_reg ( .D(c0nm_v0m_n64), .CK(clk), .QN(n138) );
  DFFQN_X1M_A12TR c0sm_v0m_full_reg ( .D(c0sm_v0m_n64), .CK(clk), .QN(n70) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_1_ ( .D(n920), .CK(clk), .QN(n127)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_1_ ( .D(n851), .CK(clk), .QN(n17)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_1_ ( .D(n863), .CK(clk), .QN(n16)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_1_ ( .D(n932), .CK(clk), .QN(n126)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_0_ ( .D(n921), .CK(clk), .QN(n131)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_0_ ( .D(n933), .CK(clk), .QN(n130)
         );
  DFFQN_X1M_A12TR s0m_m1m_state1_reg ( .D(s0m_m1m_n10), .CK(clk), .QN(n73) );
  DFFQN_X1M_A12TR s0m_m0m_state1_reg ( .D(s0m_m0m_n10), .CK(clk), .QN(n7) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_7_ ( .D(n897), .CK(clk), .QN(n245) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_6_ ( .D(n898), .CK(clk), .QN(n244) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_5_ ( .D(n899), .CK(clk), .QN(n243) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_4_ ( .D(n900), .CK(clk), .QN(n242) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_3_ ( .D(n901), .CK(clk), .QN(n241) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_2_ ( .D(n902), .CK(clk), .QN(n240) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_11_ ( .D(n893), .CK(clk), .QN(n119)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_10_ ( .D(n894), .CK(clk), .QN(n114)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_9_ ( .D(n895), .CK(clk), .QN(n109) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_8_ ( .D(n896), .CK(clk), .QN(n104) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_6_ ( .D(n834), .CK(clk), .QN(n318) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_5_ ( .D(n835), .CK(clk), .QN(n317) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_7_ ( .D(n833), .CK(clk), .QN(n319) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_4_ ( .D(n836), .CK(clk), .QN(n316) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_2_ ( .D(n838), .CK(clk), .QN(n314) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_3_ ( .D(n837), .CK(clk), .QN(n315) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_8_ ( .D(n832), .CK(clk), .QN(n24) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_9_ ( .D(n831), .CK(clk), .QN(n23) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_10_ ( .D(n830), .CK(clk), .QN(n22) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_11_ ( .D(n829), .CK(clk), .QN(n21) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_1_ ( .D(n875), .CK(clk), .QN(n15)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_1_ ( .D(n944), .CK(clk), .QN(n125)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_0_ ( .D(n864), .CK(clk), .QN(n20)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_0_ ( .D(n852), .CK(clk), .QN(n145)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_1_ ( .D(n956), .CK(clk), .QN(n128)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_1_ ( .D(n886), .CK(clk), .QN(n18)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_0_ ( .D(n876), .CK(clk), .QN(n19)
         );
  DFFQN_X1M_A12TR c0sm_v0m_state_status_reg_1_ ( .D(c0sm_v0m_n58), .CK(clk), 
        .QN(n13) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_0_ ( .D(n945), .CK(clk), .QN(n129)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_0_ ( .D(n887), .CK(clk), .QN(n144)
         );
  DFFQN_X1M_A12TR c0nm_v0m_state_swreq_reg_1_ ( .D(n908), .CK(clk), .QN(n79)
         );
  DFFQN_X1M_A12TR c0nm_v0m_state_swreq_reg_0_ ( .D(n909), .CK(clk), .QN(n76)
         );
  DFFQN_X1M_A12TR c0sm_v0m_state_queuelen_reg_1_ ( .D(c0sm_v0m_n62), .CK(clk), 
        .QN(n69) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_3_ ( .D(n918), .CK(clk), .QN(n86)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_3_ ( .D(n849), .CK(clk), .QN(n35)
         );
  DFFQN_X1M_A12TR c0nm_v0m_state_queuelen_reg_0_ ( .D(c0nm_v0m_n61), .CK(clk), 
        .QN(n135) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_rdata_reg_0_ ( .D(n904), .CK(clk), .QN(n239) );
  DFFQN_X1M_A12TR c0nm_v0m_state_status_reg_0_ ( .D(c0nm_v0m_n57), .CK(clk), 
        .QN(n77) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_0_ ( .D(n957), .CK(clk), .QN(n132)
         );
  DFFQN_X1M_A12TR s0m_o0sm_state_invc_reg_0_ ( .D(n906), .CK(clk), .QN(n3) );
  DFFQN_X1M_A12TR s0m_o0nm_state_invc_reg_0_ ( .D(n892), .CK(clk), .QN(n1) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_rdata_reg_0_ ( .D(n840), .CK(clk), .QN(n313) );
  DFFQN_X1M_A12TR x0m_colsel0reg_reg_1_ ( .D(x0m_n4), .CK(clk), .QN(n9) );
  DFFQN_X1M_A12TR x0m_colsel1reg_reg_1_ ( .D(x0m_n6), .CK(clk), .QN(n4) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_tail_reg_0_ ( .D(n968), .CK(clk), .QN(n148) );
  DFFQN_X1M_A12TR c0nm_v0m_state_status_reg_1_ ( .D(c0nm_v0m_n58), .CK(clk), 
        .QN(n78) );
  DFFQN_X1M_A12TR s0m_o0nm_state_credits_reg_2_ ( .D(s0m_o0nm_n38), .CK(clk), 
        .QN(n212) );
  DFFQN_X1M_A12TR s0m_o0sm_state_credits_reg_2_ ( .D(s0m_o0sm_n38), .CK(clk), 
        .QN(n219) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_11_ ( .D(n922), .CK(clk), .QN(n121) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_10_ ( .D(n923), .CK(clk), .QN(n116) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_9_ ( .D(n924), .CK(clk), .QN(n111)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_8_ ( .D(n925), .CK(clk), .QN(n106)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_2_ ( .D(n919), .CK(clk), .QN(n82)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_10_ ( .D(n854), .CK(clk), .QN(n62)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_9_ ( .D(n855), .CK(clk), .QN(n58)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_8_ ( .D(n856), .CK(clk), .QN(n54)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_2_ ( .D(n850), .CK(clk), .QN(n31)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_7_ ( .D(n950), .CK(clk), .QN(n103)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_6_ ( .D(n951), .CK(clk), .QN(n99)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_5_ ( .D(n952), .CK(clk), .QN(n95)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_7_ ( .D(n880), .CK(clk), .QN(n52)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_6_ ( .D(n881), .CK(clk), .QN(n48)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_5_ ( .D(n882), .CK(clk), .QN(n44)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_7_ ( .D(n938), .CK(clk), .QN(n100)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_6_ ( .D(n939), .CK(clk), .QN(n96)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_5_ ( .D(n940), .CK(clk), .QN(n92)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_4_ ( .D(n917), .CK(clk), .QN(n90)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_4_ ( .D(n941), .CK(clk), .QN(n88)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_7_ ( .D(n869), .CK(clk), .QN(n49)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_6_ ( .D(n870), .CK(clk), .QN(n45)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_5_ ( .D(n871), .CK(clk), .QN(n41)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_4_ ( .D(n848), .CK(clk), .QN(n39)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_4_ ( .D(n872), .CK(clk), .QN(n37)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_11_ ( .D(n865), .CK(clk), .QN(n25)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_3_ ( .D(n942), .CK(clk), .QN(n84)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_3_ ( .D(n873), .CK(clk), .QN(n33)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_4_ ( .D(n953), .CK(clk), .QN(n91)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_3_ ( .D(n954), .CK(clk), .QN(n87)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_4_ ( .D(n883), .CK(clk), .QN(n40)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_3_ ( .D(n884), .CK(clk), .QN(n36)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_2_ ( .D(n885), .CK(clk), .QN(n32)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_7_ ( .D(n914), .CK(clk), .QN(n102)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_6_ ( .D(n915), .CK(clk), .QN(n98)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_5_ ( .D(n916), .CK(clk), .QN(n94)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_3_ ( .D(n930), .CK(clk), .QN(n85)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_2_ ( .D(n943), .CK(clk), .QN(n80)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_7_ ( .D(n845), .CK(clk), .QN(n51)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_6_ ( .D(n846), .CK(clk), .QN(n47)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_5_ ( .D(n847), .CK(clk), .QN(n43)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_3_ ( .D(n861), .CK(clk), .QN(n34)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_2_ ( .D(n874), .CK(clk), .QN(n29)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_11_ ( .D(n853), .CK(clk), .QN(n26)
         );
  DFFQN_X1M_A12TR c0sm_v0m_state_status_reg_0_ ( .D(c0sm_v0m_n57), .CK(clk), 
        .QN(n12) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_11_ ( .D(n841), .CK(clk), .QN(n27)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_11_ ( .D(n934), .CK(clk), .QN(n120) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_10_ ( .D(n935), .CK(clk), .QN(n115) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_9_ ( .D(n936), .CK(clk), .QN(n110)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_8_ ( .D(n937), .CK(clk), .QN(n105)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_10_ ( .D(n866), .CK(clk), .QN(n61)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_9_ ( .D(n867), .CK(clk), .QN(n57)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_8_ ( .D(n868), .CK(clk), .QN(n53)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_11_ ( .D(n910), .CK(clk), .QN(n122) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_10_ ( .D(n911), .CK(clk), .QN(n117) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_9_ ( .D(n912), .CK(clk), .QN(n112)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_8_ ( .D(n913), .CK(clk), .QN(n107)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_2_ ( .D(n955), .CK(clk), .QN(n83)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_10_ ( .D(n842), .CK(clk), .QN(n63)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_9_ ( .D(n843), .CK(clk), .QN(n59)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_8_ ( .D(n844), .CK(clk), .QN(n55)
         );
  DFFQN_X1M_A12TR s0m_resp1_reg_1_ ( .D(n964), .CK(clk), .QN(n72) );
  DFFQN_X1M_A12TR s0m_resp1_reg_0_ ( .D(n963), .CK(clk), .QN(n10) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_11_ ( .D(n946), .CK(clk), .QN(n123) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_10_ ( .D(n947), .CK(clk), .QN(n118) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_9_ ( .D(n948), .CK(clk), .QN(n113)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_8_ ( .D(n949), .CK(clk), .QN(n108)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_10_ ( .D(n877), .CK(clk), .QN(n64)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_9_ ( .D(n878), .CK(clk), .QN(n60)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_8_ ( .D(n879), .CK(clk), .QN(n56)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_7_ ( .D(n926), .CK(clk), .QN(n101)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_6_ ( .D(n927), .CK(clk), .QN(n97)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_5_ ( .D(n928), .CK(clk), .QN(n93)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_4_ ( .D(n929), .CK(clk), .QN(n89)
         );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_2_ ( .D(n931), .CK(clk), .QN(n81)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_7_ ( .D(n857), .CK(clk), .QN(n50)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_6_ ( .D(n858), .CK(clk), .QN(n46)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_5_ ( .D(n859), .CK(clk), .QN(n42)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_4_ ( .D(n860), .CK(clk), .QN(n38)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_2_ ( .D(n862), .CK(clk), .QN(n30)
         );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_11_ ( .D(n966), .CK(clk), .QN(n28)
         );
  DFFQN_X1M_A12TR c0sm_v0m_state_swreq_reg_1_ ( .D(n965), .CK(clk), .QN(n14)
         );
  DFFQN_X1M_A12TR c0sm_v0m_state_swreq_reg_0_ ( .D(n962), .CK(clk), .QN(n11)
         );
  DFFQN_X1M_A12TR s0m_o0nm_state_credits_reg_1_ ( .D(s0m_o0nm_n37), .CK(clk), 
        .QN(n141) );
  DFFQN_X1M_A12TR s0m_o0sm_state_credits_reg_1_ ( .D(s0m_o0sm_n37), .CK(clk), 
        .QN(n74) );
  DFFQN_X1M_A12TR c0sm_v0m_state_queuelen_reg_0_ ( .D(c0sm_v0m_n61), .CK(clk), 
        .QN(n67) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_head_reg_0_ ( .D(n960), .CK(clk), .QN(n134) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_head_reg_0_ ( .D(n890), .CK(clk), .QN(n66) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_tail_reg_1_ ( .D(n970), .CK(clk), .QN(n150) );
  DFFQN_X1M_A12TR x0m_colsel0reg_reg_0_ ( .D(x0m_n3), .CK(clk), .QN(n8) );
  DFFQN_X1M_A12TR s0m_o0nm_state_credits_reg_0_ ( .D(s0m_o0nm_n36), .CK(clk), 
        .QN(n142) );
  DFFQN_X1M_A12TR s0m_o0sm_state_credits_reg_0_ ( .D(s0m_o0sm_n36), .CK(clk), 
        .QN(n75) );
  DFFQN_X1M_A12TR c0sm_b0m_v0m_tail_reg_1_ ( .D(n967), .CK(clk), .QN(n147) );
  DFFQN_X1M_A12TR x0m_colsel1reg_reg_0_ ( .D(x0m_n5), .CK(clk), .QN(n5) );
  DFFQN_X1M_A12TR c0nm_b0m_v0m_tail_reg_0_ ( .D(n971), .CK(clk), .QN(n151) );
  NAND2B_X0P5M_A12TR u1015 ( .AN(n1261), .B(n1463), .Y(n1163) );
  NAND2_X0P5A_A12TR u1016 ( .A(n1413), .B(curry[0]), .Y(n973) );
  CGENI_X1M_A12TR u1017 ( .A(n1414), .B(n1034), .CI(n973), .CON(n974) );
  CGENI_X1M_A12TR u1018 ( .A(n1416), .B(curry[2]), .CI(n974), .CON(n975) );
  CGEN_X1M_A12TR u1019 ( .A(currx[0]), .B(n1417), .CI(n975), .CO(n976) );
  CGEN_X1M_A12TR u1020 ( .A(n1418), .B(currx[1]), .CI(n976), .CO(n977) );
  CGENI_X1M_A12TR u1021 ( .A(currx[2]), .B(n1419), .CI(n977), .CON(n1040) );
  NAND2_X0P5A_A12TR u1022 ( .A(curry[0]), .B(n1245), .Y(n978) );
  CGENI_X1M_A12TR u1023 ( .A(n1246), .B(n1034), .CI(n978), .CON(n979) );
  CGENI_X1M_A12TR u1024 ( .A(n1248), .B(curry[2]), .CI(n979), .CON(n980) );
  CGEN_X1M_A12TR u1025 ( .A(currx[0]), .B(n1249), .CI(n980), .CO(n981) );
  CGEN_X1M_A12TR u1026 ( .A(n1250), .B(currx[1]), .CI(n981), .CO(n982) );
  CGENI_X1M_A12TR u1027 ( .A(currx[2]), .B(n1251), .CI(n982), .CON(n1009) );
  NOR2_X0P5A_A12TR u1028 ( .A(n1472), .B(n1473), .Y(n983) );
  AOI22_X0P5M_A12TR u1029 ( .A0(n75), .A1(n1474), .B0(n1476), .B1(n1471), .Y(
        n984) );
  NAND2_X0P5A_A12TR u1030 ( .A(n74), .B(n984), .Y(n985) );
  OAI211_X0P5M_A12TR u1031 ( .A0(n983), .A1(n74), .B0(n1485), .C0(n985), .Y(
        s0m_o0sm_n37) );
  NOR2_X0P5A_A12TR u1032 ( .A(n1450), .B(n1451), .Y(n986) );
  AOI22_X0P5M_A12TR u1033 ( .A0(n142), .A1(n1452), .B0(n1454), .B1(n1449), .Y(
        n987) );
  NAND2_X0P5A_A12TR u1034 ( .A(n141), .B(n987), .Y(n988) );
  OAI211_X0P5M_A12TR u1035 ( .A0(n986), .A1(n141), .B0(n1485), .C0(n988), .Y(
        s0m_o0nm_n37) );
  OAI21_X0P5M_A12TR u1036 ( .A0(n1463), .A1(n1167), .B0(n1485), .Y(n989) );
  NAND3B_X0P5M_A12TR u1037 ( .AN(n1090), .B(n1018), .C(n1017), .Y(n990) );
  OAI22_X0P5M_A12TR u1038 ( .A0(n138), .A1(n989), .B0(n1268), .B1(n990), .Y(
        c0nm_v0m_n64) );
  INV_X1M_A12TR u1039 ( .A(reset), .Y(n1485) );
  OAI221_X1M_A12TR u1040 ( .A0(n1244), .A1(n1243), .B0(n1463), .B1(n1242), 
        .C0(n1485), .Y(n903) );
  OAI221_X1M_A12TR u1041 ( .A0(n1466), .A1(n1412), .B0(n1411), .B1(n1410), 
        .C0(n1485), .Y(n839) );
  NOR2_X1M_A12TR u1042 ( .A(s0m_o0nm_n42), .B(s0m_o0nm_n35), .Y(s0m_o0nm_n41)
         );
  NOR2_X1M_A12TR u1043 ( .A(n1442), .B(n1441), .Y(s0m_o0nm_n35) );
  NOR2_X1M_A12TR u1044 ( .A(n1443), .B(s0m_o0nm_state_assigned), .Y(n1442) );
  NOR2_X1M_A12TR u1045 ( .A(s0m_o0sm_n42), .B(s0m_o0sm_n35), .Y(s0m_o0sm_n41)
         );
  NOR2_X1M_A12TR u1046 ( .A(n1462), .B(n1461), .Y(s0m_o0sm_n35) );
  NOR2_X1M_A12TR u1047 ( .A(n1464), .B(s0m_o0sm_state_assigned), .Y(n1462) );
  OA21A1OI2_X1M_A12TR u1048 ( .A0(n1460), .A1(n1459), .B0(n1458), .C0(reset), 
        .Y(s0m_o0nm_n42) );
  NAND2_X1M_A12TR u1049 ( .A(s0m_no_bufs0), .B(n1457), .Y(n1458) );
  OA21A1OI2_X1M_A12TR u1050 ( .A0(n1482), .A1(n1481), .B0(n1480), .C0(reset), 
        .Y(s0m_o0sm_n42) );
  NAND2_X1M_A12TR u1051 ( .A(s0m_no_bufs1), .B(n1479), .Y(n1480) );
  AOI221_X1M_A12TR u1052 ( .A0(n1183), .A1(n1244), .B0(n1089), .B1(n1463), 
        .C0(n1088), .Y(n959) );
  NAND2_X1M_A12TR u1053 ( .A(n1485), .B(n1261), .Y(n1088) );
  AOI221_X1M_A12TR u1054 ( .A0(n1362), .A1(n1466), .B0(n1276), .B1(n1411), 
        .C0(n1275), .Y(n889) );
  NAND2_X1M_A12TR u1055 ( .A(n1485), .B(n1429), .Y(n1275) );
  OA21A1OI2_X1M_A12TR u1056 ( .A0(n1486), .A1(n1437), .B0(n140), .C0(n1240), 
        .Y(n905) );
  OA21A1OI2_X1M_A12TR u1057 ( .A0(n1483), .A1(n1439), .B0(n6), .C0(n1240), .Y(
        n961) );
  OA21A1OI2_X1M_A12TR u1058 ( .A0(n143), .A1(n1443), .B0(n1273), .C0(n1441), 
        .Y(n891) );
  OA21A1OI2_X1M_A12TR u1059 ( .A0(n2), .A1(n1464), .B0(n1238), .C0(n1461), .Y(
        n907) );
  NOR2_X1M_A12TR u1060 ( .A(n1009), .B(n1008), .Y(c0nm_r0m_n10) );
  OA21A1OI2_X1M_A12TR u1061 ( .A0(n137), .A1(n1244), .B0(n1016), .C0(reset), 
        .Y(c0nm_v0m_n62) );
  OAI22_X1M_A12TR u1062 ( .A0(n1015), .A1(n1018), .B0(n1014), .B1(n1017), .Y(
        n1016) );
  NAND3_X1M_A12TR u1063 ( .A(n1241), .B(n1485), .C(n1099), .Y(n1008) );
  NOR2_X1M_A12TR u1064 ( .A(n1040), .B(n1039), .Y(c0sm_r0m_n10) );
  NAND3_X1M_A12TR u1065 ( .A(n1409), .B(n1485), .C(n1284), .Y(n1039) );
  INV_X1M_A12TR u1066 ( .A(curry[1]), .Y(n1034) );
  OAI31_X1M_A12TR u1067 ( .A0(n1051), .A1(n1436), .A2(n1077), .B0(n1050), .Y(
        c0sm_v0m_n64) );
  OAI211_X1M_A12TR u1068 ( .A0(n1411), .A1(n1346), .B0(n1485), .C0(n1049), .Y(
        n1050) );
  INV_X1M_A12TR u1069 ( .A(n70), .Y(n1049) );
  AOI32_X1M_A12TR u1070 ( .A0(n1203), .A1(n1229), .A2(n1485), .B0(n1202), .B1(
        n127), .Y(n920) );
  AOI22_X1M_A12TR u1071 ( .A0(n1206), .A1(n1201), .B0(n1200), .B1(n1204), .Y(
        n1203) );
  AOI32_X1M_A12TR u1072 ( .A0(n1382), .A1(n1408), .A2(n1485), .B0(n1381), .B1(
        n17), .Y(n851) );
  AOI22_X1M_A12TR u1073 ( .A0(n1385), .A1(n1380), .B0(n1379), .B1(n1383), .Y(
        n1382) );
  AOI32_X1M_A12TR u1074 ( .A0(n1369), .A1(n1375), .A2(n1485), .B0(n1368), .B1(
        n16), .Y(n863) );
  AOI22_X1M_A12TR u1075 ( .A0(n1372), .A1(n1380), .B0(n1379), .B1(n1370), .Y(
        n1369) );
  AOI32_X1M_A12TR u1076 ( .A0(n1190), .A1(n1196), .A2(n1485), .B0(n1189), .B1(
        n126), .Y(n932) );
  AOI22_X1M_A12TR u1077 ( .A0(n1193), .A1(n1201), .B0(n1200), .B1(n1191), .Y(
        n1190) );
  AOI32_X1M_A12TR u1078 ( .A0(n1199), .A1(n1229), .A2(n1485), .B0(n1202), .B1(
        n131), .Y(n921) );
  INV_X1M_A12TR u1079 ( .A(n1229), .Y(n1202) );
  AOI22_X1M_A12TR u1080 ( .A0(n1206), .A1(n1198), .B0(n1197), .B1(n1204), .Y(
        n1199) );
  AOI32_X1M_A12TR u1081 ( .A0(n1188), .A1(n1196), .A2(n1485), .B0(n1189), .B1(
        n130), .Y(n933) );
  INV_X1M_A12TR u1082 ( .A(n1196), .Y(n1189) );
  AOI22_X1M_A12TR u1083 ( .A0(n1193), .A1(n1198), .B0(n1197), .B1(n1191), .Y(
        n1188) );
  OA21A1OI2_X1M_A12TR u1084 ( .A0(n1440), .A1(n73), .B0(n1439), .C0(reset), 
        .Y(s0m_m1m_n10) );
  OA21A1OI2_X1M_A12TR u1085 ( .A0(n1438), .A1(n7), .B0(n1437), .C0(reset), .Y(
        s0m_m0m_n10) );
  OAI22_X1M_A12TR u1086 ( .A0(n1251), .A1(n168), .B0(n245), .B1(n1268), .Y(
        n897) );
  NOR2_X1M_A12TR u1087 ( .A(n997), .B(n996), .Y(n1251) );
  OAI22_X1M_A12TR u1088 ( .A0(n101), .A1(n1263), .B0(n100), .B1(n1264), .Y(
        n996) );
  OAI22_X1M_A12TR u1089 ( .A0(n102), .A1(n1262), .B0(n103), .B1(n1261), .Y(
        n997) );
  OAI22_X1M_A12TR u1090 ( .A0(n1250), .A1(n168), .B0(n244), .B1(n1268), .Y(
        n898) );
  NOR2_X1M_A12TR u1091 ( .A(n1007), .B(n1006), .Y(n1250) );
  OAI22_X1M_A12TR u1092 ( .A0(n97), .A1(n1263), .B0(n96), .B1(n1264), .Y(n1006) );
  OAI22_X1M_A12TR u1093 ( .A0(n98), .A1(n1262), .B0(n99), .B1(n1261), .Y(n1007) );
  OAI22_X1M_A12TR u1094 ( .A0(n1249), .A1(n168), .B0(n243), .B1(n1268), .Y(
        n899) );
  NOR2_X1M_A12TR u1095 ( .A(n1005), .B(n1004), .Y(n1249) );
  OAI22_X1M_A12TR u1096 ( .A0(n93), .A1(n1263), .B0(n92), .B1(n1264), .Y(n1004) );
  OAI22_X1M_A12TR u1097 ( .A0(n94), .A1(n1262), .B0(n95), .B1(n1261), .Y(n1005) );
  OAI22_X1M_A12TR u1098 ( .A0(n1248), .A1(n168), .B0(n242), .B1(n1268), .Y(
        n900) );
  NOR2_X1M_A12TR u1099 ( .A(n999), .B(n998), .Y(n1248) );
  OAI22_X1M_A12TR u1100 ( .A0(n88), .A1(n1264), .B0(n90), .B1(n1262), .Y(n998)
         );
  OAI22_X1M_A12TR u1101 ( .A0(n91), .A1(n1261), .B0(n89), .B1(n1263), .Y(n999)
         );
  OAI22_X1M_A12TR u1102 ( .A0(n1247), .A1(n168), .B0(n241), .B1(n1268), .Y(
        n901) );
  INV_X1M_A12TR u1103 ( .A(n1246), .Y(n1247) );
  OAI21_X1M_A12TR u1104 ( .A0(n84), .A1(n1264), .B0(n1001), .Y(n1246) );
  AOI21_X1M_A12TR u1105 ( .A0(n1205), .A1(n1115), .B0(n1000), .Y(n1001) );
  OAI22_X1M_A12TR u1106 ( .A0(n87), .A1(n1261), .B0(n85), .B1(n1263), .Y(n1000) );
  OAI22_X1M_A12TR u1107 ( .A0(n1245), .A1(n168), .B0(n240), .B1(n1268), .Y(
        n902) );
  NOR2_X1M_A12TR u1108 ( .A(n1003), .B(n1002), .Y(n1245) );
  OAI22_X1M_A12TR u1109 ( .A0(n81), .A1(n1263), .B0(n82), .B1(n1262), .Y(n1002) );
  OAI22_X1M_A12TR u1110 ( .A0(n83), .A1(n1261), .B0(n80), .B1(n1264), .Y(n1003) );
  OAI21_X1M_A12TR u1111 ( .A0(n119), .A1(n1268), .B0(n1267), .Y(n893) );
  OAI21_X1M_A12TR u1112 ( .A0(n1266), .A1(n1265), .B0(creditout_0), .Y(n1267)
         );
  OAI22_X1M_A12TR u1113 ( .A0(n120), .A1(n1264), .B0(n121), .B1(n1263), .Y(
        n1265) );
  OAI22_X1M_A12TR u1114 ( .A0(n122), .A1(n1262), .B0(n123), .B1(n1261), .Y(
        n1266) );
  OAI21_X1M_A12TR u1115 ( .A0(n114), .A1(n1268), .B0(n1260), .Y(n894) );
  OAI21_X1M_A12TR u1116 ( .A0(n1259), .A1(n1258), .B0(creditout_0), .Y(n1260)
         );
  OAI22_X1M_A12TR u1117 ( .A0(n115), .A1(n1264), .B0(n116), .B1(n1263), .Y(
        n1258) );
  OAI22_X1M_A12TR u1118 ( .A0(n117), .A1(n1262), .B0(n118), .B1(n1261), .Y(
        n1259) );
  OAI21_X1M_A12TR u1119 ( .A0(n109), .A1(n1268), .B0(n1257), .Y(n895) );
  OAI21_X1M_A12TR u1120 ( .A0(n1256), .A1(n1255), .B0(creditout_0), .Y(n1257)
         );
  OAI22_X1M_A12TR u1121 ( .A0(n110), .A1(n1264), .B0(n111), .B1(n1263), .Y(
        n1255) );
  OAI22_X1M_A12TR u1122 ( .A0(n112), .A1(n1262), .B0(n113), .B1(n1261), .Y(
        n1256) );
  OAI21_X1M_A12TR u1123 ( .A0(n104), .A1(n1268), .B0(n1254), .Y(n896) );
  OAI21_X1M_A12TR u1124 ( .A0(n1253), .A1(n1252), .B0(creditout_0), .Y(n1254)
         );
  OAI22_X1M_A12TR u1125 ( .A0(n105), .A1(n1264), .B0(n106), .B1(n1263), .Y(
        n1252) );
  OAI22_X1M_A12TR u1126 ( .A0(n107), .A1(n1262), .B0(n108), .B1(n1261), .Y(
        n1253) );
  OAI22_X1M_A12TR u1127 ( .A0(n1418), .A1(n158), .B0(n318), .B1(n1436), .Y(
        n834) );
  NOR2_X1M_A12TR u1128 ( .A(n1038), .B(n1037), .Y(n1418) );
  OAI22_X1M_A12TR u1129 ( .A0(n46), .A1(n1431), .B0(n45), .B1(n1432), .Y(n1037) );
  OAI22_X1M_A12TR u1130 ( .A0(n47), .A1(n1430), .B0(n48), .B1(n1429), .Y(n1038) );
  OAI22_X1M_A12TR u1131 ( .A0(n1417), .A1(n158), .B0(n317), .B1(n1436), .Y(
        n835) );
  NOR2_X1M_A12TR u1132 ( .A(n1036), .B(n1035), .Y(n1417) );
  OAI22_X1M_A12TR u1133 ( .A0(n42), .A1(n1431), .B0(n41), .B1(n1432), .Y(n1035) );
  OAI22_X1M_A12TR u1134 ( .A0(n43), .A1(n1430), .B0(n44), .B1(n1429), .Y(n1036) );
  OAI22_X1M_A12TR u1135 ( .A0(n1419), .A1(n158), .B0(n319), .B1(n1436), .Y(
        n833) );
  NOR2_X1M_A12TR u1136 ( .A(n1027), .B(n1026), .Y(n1419) );
  OAI22_X1M_A12TR u1137 ( .A0(n50), .A1(n1431), .B0(n49), .B1(n1432), .Y(n1026) );
  OAI22_X1M_A12TR u1138 ( .A0(n51), .A1(n1430), .B0(n52), .B1(n1429), .Y(n1027) );
  OAI22_X1M_A12TR u1139 ( .A0(n1416), .A1(n158), .B0(n316), .B1(n1436), .Y(
        n836) );
  NOR2_X1M_A12TR u1140 ( .A(n1029), .B(n1028), .Y(n1416) );
  OAI22_X1M_A12TR u1141 ( .A0(n37), .A1(n1432), .B0(n39), .B1(n1430), .Y(n1028) );
  OAI22_X1M_A12TR u1142 ( .A0(n40), .A1(n1429), .B0(n38), .B1(n1431), .Y(n1029) );
  OAI22_X1M_A12TR u1143 ( .A0(n1413), .A1(n158), .B0(n314), .B1(n1436), .Y(
        n838) );
  NOR2_X1M_A12TR u1144 ( .A(n1033), .B(n1032), .Y(n1413) );
  OAI22_X1M_A12TR u1145 ( .A0(n30), .A1(n1431), .B0(n31), .B1(n1430), .Y(n1032) );
  OAI22_X1M_A12TR u1146 ( .A0(n32), .A1(n1429), .B0(n29), .B1(n1432), .Y(n1033) );
  OAI22_X1M_A12TR u1147 ( .A0(n1415), .A1(n158), .B0(n315), .B1(n1436), .Y(
        n837) );
  INV_X1M_A12TR u1148 ( .A(n1414), .Y(n1415) );
  OAI21_X1M_A12TR u1149 ( .A0(n33), .A1(n1432), .B0(n1031), .Y(n1414) );
  AOI21_X1M_A12TR u1150 ( .A0(n1384), .A1(n1300), .B0(n1030), .Y(n1031) );
  OAI22_X1M_A12TR u1151 ( .A0(n36), .A1(n1429), .B0(n34), .B1(n1431), .Y(n1030) );
  OAI21_X1M_A12TR u1152 ( .A0(n24), .A1(n1436), .B0(n1422), .Y(n832) );
  OAI21_X1M_A12TR u1153 ( .A0(n1421), .A1(n1420), .B0(creditout_1), .Y(n1422)
         );
  OAI22_X1M_A12TR u1154 ( .A0(n53), .A1(n1432), .B0(n54), .B1(n1431), .Y(n1420) );
  OAI22_X1M_A12TR u1155 ( .A0(n55), .A1(n1430), .B0(n56), .B1(n1429), .Y(n1421) );
  OAI21_X1M_A12TR u1156 ( .A0(n23), .A1(n1436), .B0(n1425), .Y(n831) );
  OAI21_X1M_A12TR u1157 ( .A0(n1424), .A1(n1423), .B0(creditout_1), .Y(n1425)
         );
  OAI22_X1M_A12TR u1158 ( .A0(n57), .A1(n1432), .B0(n58), .B1(n1431), .Y(n1423) );
  OAI22_X1M_A12TR u1159 ( .A0(n59), .A1(n1430), .B0(n60), .B1(n1429), .Y(n1424) );
  OAI21_X1M_A12TR u1160 ( .A0(n22), .A1(n1436), .B0(n1428), .Y(n830) );
  OAI21_X1M_A12TR u1161 ( .A0(n1427), .A1(n1426), .B0(creditout_1), .Y(n1428)
         );
  OAI22_X1M_A12TR u1162 ( .A0(n61), .A1(n1432), .B0(n62), .B1(n1431), .Y(n1426) );
  OAI22_X1M_A12TR u1163 ( .A0(n63), .A1(n1430), .B0(n64), .B1(n1429), .Y(n1427) );
  OAI21_X1M_A12TR u1164 ( .A0(n21), .A1(n1436), .B0(n1435), .Y(n829) );
  OAI21_X1M_A12TR u1165 ( .A0(n1434), .A1(n1433), .B0(creditout_1), .Y(n1435)
         );
  OAI22_X1M_A12TR u1166 ( .A0(n25), .A1(n1432), .B0(n26), .B1(n1431), .Y(n1433) );
  OAI22_X1M_A12TR u1167 ( .A0(n27), .A1(n1430), .B0(n28), .B1(n1429), .Y(n1434) );
  AOI32_X1M_A12TR u1168 ( .A0(n1360), .A1(n1366), .A2(n1485), .B0(n1359), .B1(
        n15), .Y(n875) );
  AOI22_X1M_A12TR u1169 ( .A0(n1363), .A1(n1380), .B0(n1379), .B1(n1361), .Y(
        n1360) );
  AOI32_X1M_A12TR u1170 ( .A0(n1181), .A1(n1187), .A2(n1485), .B0(n1180), .B1(
        n125), .Y(n944) );
  AOI22_X1M_A12TR u1171 ( .A0(n1184), .A1(n1201), .B0(n1200), .B1(n1182), .Y(
        n1181) );
  AOI32_X1M_A12TR u1172 ( .A0(n1367), .A1(n1375), .A2(n1485), .B0(n1368), .B1(
        n20), .Y(n864) );
  INV_X1M_A12TR u1173 ( .A(n1375), .Y(n1368) );
  AOI22_X1M_A12TR u1174 ( .A0(n1372), .A1(n1377), .B0(n1376), .B1(n1370), .Y(
        n1367) );
  AOI32_X1M_A12TR u1175 ( .A0(n1378), .A1(n1408), .A2(n1485), .B0(n1381), .B1(
        n145), .Y(n852) );
  INV_X1M_A12TR u1176 ( .A(n1408), .Y(n1381) );
  AOI22_X1M_A12TR u1177 ( .A0(n1385), .A1(n1377), .B0(n1376), .B1(n1383), .Y(
        n1378) );
  AOI32_X1M_A12TR u1178 ( .A0(n1101), .A1(n1176), .A2(n1485), .B0(n1100), .B1(
        n128), .Y(n956) );
  AOI22_X1M_A12TR u1179 ( .A0(n1105), .A1(n1201), .B0(n1200), .B1(n1102), .Y(
        n1101) );
  NAND2_X1M_A12TR u1180 ( .A(n1242), .B(n1463), .Y(n1200) );
  INV_X1M_A12TR u1181 ( .A(n1099), .Y(n1242) );
  OAI21_X1M_A12TR u1182 ( .A0(n125), .A1(n1264), .B0(n995), .Y(n1099) );
  OAI22_X1M_A12TR u1183 ( .A0(n126), .A1(n1263), .B0(n128), .B1(n1261), .Y(
        n994) );
  OAI211_X1M_A12TR u1184 ( .A0(n125), .A1(n1173), .B0(n1098), .C0(n1097), .Y(
        n1201) );
  AOI22_X1M_A12TR u1185 ( .A0(flitin_0[1]), .A1(n1167), .B0(n1169), .B1(n1096), 
        .Y(n1098) );
  INV_X1M_A12TR u1186 ( .A(n128), .Y(n1096) );
  AOI32_X1M_A12TR u1187 ( .A0(n1288), .A1(n1355), .A2(n1485), .B0(n1287), .B1(
        n18), .Y(n886) );
  AOI22_X1M_A12TR u1188 ( .A0(n1286), .A1(n1380), .B0(n1379), .B1(n1285), .Y(
        n1288) );
  NAND2_X1M_A12TR u1189 ( .A(n1410), .B(n1411), .Y(n1379) );
  INV_X1M_A12TR u1190 ( .A(n1284), .Y(n1410) );
  OAI21_X1M_A12TR u1191 ( .A0(n16), .A1(n1431), .B0(n1025), .Y(n1284) );
  OAI22_X1M_A12TR u1192 ( .A0(n15), .A1(n1432), .B0(n18), .B1(n1429), .Y(n1024) );
  OAI211_X1M_A12TR u1193 ( .A0(n15), .A1(n1352), .B0(n1283), .C0(n1282), .Y(
        n1380) );
  AOI22_X1M_A12TR u1194 ( .A0(flitin_1[1]), .A1(n1346), .B0(n1348), .B1(n1281), 
        .Y(n1283) );
  INV_X1M_A12TR u1195 ( .A(n18), .Y(n1281) );
  AOI32_X1M_A12TR u1196 ( .A0(n1358), .A1(n1366), .A2(n1485), .B0(n1359), .B1(
        n19), .Y(n876) );
  INV_X1M_A12TR u1197 ( .A(n1366), .Y(n1359) );
  AOI22_X1M_A12TR u1198 ( .A0(n1363), .A1(n1377), .B0(n1376), .B1(n1361), .Y(
        n1358) );
  OAI21_X1M_A12TR u1199 ( .A0(n13), .A1(n1082), .B0(n1081), .Y(c0sm_v0m_n58)
         );
  AOI32_X1M_A12TR u1200 ( .A0(n1179), .A1(n1187), .A2(n1485), .B0(n1180), .B1(
        n129), .Y(n945) );
  INV_X1M_A12TR u1201 ( .A(n1187), .Y(n1180) );
  AOI22_X1M_A12TR u1202 ( .A0(n1184), .A1(n1198), .B0(n1197), .B1(n1182), .Y(
        n1179) );
  AOI32_X1M_A12TR u1203 ( .A0(n1280), .A1(n1355), .A2(n1485), .B0(n1287), .B1(
        n144), .Y(n887) );
  INV_X1M_A12TR u1204 ( .A(n1355), .Y(n1287) );
  AOI22_X1M_A12TR u1205 ( .A0(n1286), .A1(n1377), .B0(n1376), .B1(n1285), .Y(
        n1280) );
  NAND2_X1M_A12TR u1206 ( .A(n1409), .B(n1411), .Y(n1376) );
  OAI21_X1M_A12TR u1207 ( .A0(n19), .A1(n1352), .B0(n1279), .Y(n1377) );
  AOI211_X1M_A12TR u1208 ( .A0(flitin_1[0]), .A1(n1346), .B0(n1278), .C0(n1277), .Y(n1279) );
  OAI22_X1M_A12TR u1209 ( .A0(n145), .A1(n1350), .B0(n20), .B1(n1351), .Y(
        n1277) );
  NOR2_X1M_A12TR u1210 ( .A(n144), .B(n1323), .Y(n1278) );
  OAI22_X1M_A12TR u1211 ( .A0(n194), .A1(n1234), .B0(n79), .B1(n1233), .Y(n908) );
  OAI22_X1M_A12TR u1212 ( .A0(n193), .A1(n1234), .B0(n76), .B1(n1233), .Y(n909) );
  NAND2_X1M_A12TR u1213 ( .A(n1230), .B(n1232), .Y(n1234) );
  OA21A1OI2_X1M_A12TR u1214 ( .A0(n69), .A1(n1466), .B0(n1048), .C0(reset), 
        .Y(c0sm_v0m_n62) );
  OAI22_X1M_A12TR u1215 ( .A0(n1047), .A1(n1046), .B0(n1045), .B1(n1044), .Y(
        n1048) );
  OAI222_X1M_A12TR u1216 ( .A0(n1229), .A1(n86), .B0(n1228), .B1(n1210), .C0(
        n1226), .C1(n1209), .Y(n918) );
  OAI222_X1M_A12TR u1217 ( .A0(n1408), .A1(n35), .B0(n1407), .B1(n1389), .C0(
        n1405), .C1(n1388), .Y(n849) );
  AOI21_X1M_A12TR u1218 ( .A0(n135), .A1(n1014), .B0(n1013), .Y(c0nm_v0m_n61)
         );
  OAI21_X1M_A12TR u1219 ( .A0(n135), .A1(n1014), .B0(n1485), .Y(n1013) );
  AOI31_X1M_A12TR u1220 ( .A0(n1090), .A1(n1244), .A2(n138), .B0(n1015), .Y(
        n1014) );
  AOI211_X1M_A12TR u1221 ( .A0(n1018), .A1(n1017), .B0(n1090), .C0(n1244), .Y(
        n1015) );
  OAI221_X1M_A12TR u1222 ( .A0(n1244), .A1(n239), .B0(n1463), .B1(n1241), .C0(
        n1485), .Y(n904) );
  INV_X1M_A12TR u1223 ( .A(n1463), .Y(n1244) );
  AOI32_X1M_A12TR u1224 ( .A0(n1095), .A1(n1176), .A2(n1485), .B0(n1100), .B1(
        n132), .Y(n957) );
  INV_X1M_A12TR u1225 ( .A(n1176), .Y(n1100) );
  AOI22_X1M_A12TR u1226 ( .A0(n1105), .A1(n1198), .B0(n1197), .B1(n1102), .Y(
        n1095) );
  NAND2_X1M_A12TR u1227 ( .A(n1241), .B(n1463), .Y(n1197) );
  NOR2_X1M_A12TR u1228 ( .A(n993), .B(n992), .Y(n1241) );
  OAI222_X1M_A12TR u1229 ( .A0(n1261), .A1(n132), .B0(n1263), .B1(n130), .C0(
        n1262), .C1(n131), .Y(n992) );
  NOR2_X1M_A12TR u1230 ( .A(n129), .B(n1264), .Y(n993) );
  OAI211_X1M_A12TR u1231 ( .A0(n129), .A1(n1173), .B0(n1094), .C0(n1093), .Y(
        n1198) );
  AOI22_X1M_A12TR u1232 ( .A0(flitin_0[0]), .A1(n1167), .B0(n1169), .B1(n1091), 
        .Y(n1094) );
  INV_X1M_A12TR u1233 ( .A(n132), .Y(n1091) );
  OA21A1OI2_X1M_A12TR u1234 ( .A0(n3), .A1(n1464), .B0(n1439), .C0(n1461), .Y(
        n906) );
  NAND2_X1M_A12TR u1235 ( .A(n1237), .B(n1485), .Y(n1461) );
  AOI22_X1M_A12TR u1236 ( .A0(tailout_1), .A1(n1467), .B0(n1270), .B1(n1236), 
        .Y(n1237) );
  OAI211_X1M_A12TR u1237 ( .A0(n14), .A1(n73), .B0(s0m_elig_1_), .C0(n1086), 
        .Y(n1439) );
  OA21A1OI2_X1M_A12TR u1238 ( .A0(n1), .A1(n1443), .B0(n1437), .C0(n1441), .Y(
        n892) );
  NAND2_X1M_A12TR u1239 ( .A(n1272), .B(n1485), .Y(n1441) );
  AOI22_X1M_A12TR u1240 ( .A0(tailout_1), .A1(n1445), .B0(n1271), .B1(n1270), 
        .Y(n1272) );
  OAI211_X1M_A12TR u1241 ( .A0(n11), .A1(n7), .B0(s0m_elig_0_), .C0(n1239), 
        .Y(n1437) );
  OAI221_X1M_A12TR u1242 ( .A0(n1466), .A1(n313), .B0(n1411), .B1(n1409), .C0(
        n1485), .Y(n840) );
  NOR2_X1M_A12TR u1243 ( .A(n1023), .B(n1022), .Y(n1409) );
  OAI222_X1M_A12TR u1244 ( .A0(n1430), .A1(n145), .B0(n1429), .B1(n144), .C0(
        n1432), .C1(n19), .Y(n1022) );
  NOR2_X1M_A12TR u1245 ( .A(n20), .B(n1431), .Y(n1023) );
  OAI21_X1M_A12TR u1246 ( .A0(n1484), .A1(n1483), .B0(n1485), .Y(x0m_n4) );
  OAI21_X1M_A12TR u1247 ( .A0(n1487), .A1(n1486), .B0(n1485), .Y(x0m_n6) );
  OAI21_X1M_A12TR u1248 ( .A0(n78), .A1(n1232), .B0(n1231), .Y(c0nm_v0m_n58)
         );
  NOR2_X1M_A12TR u1249 ( .A(n1012), .B(n1240), .Y(n1231) );
  INV_X1M_A12TR u1250 ( .A(n1230), .Y(n1240) );
  NOR2_X1M_A12TR u1251 ( .A(reset), .B(n1270), .Y(n1230) );
  AOI211_X1M_A12TR u1252 ( .A0(n193), .A1(n194), .B0(n77), .C0(n78), .Y(n1232)
         );
  OA21A1OI2_X1M_A12TR u1253 ( .A0(n212), .A1(n1456), .B0(n1455), .C0(reset), 
        .Y(s0m_o0nm_n38) );
  OAI21_X1M_A12TR u1254 ( .A0(n212), .A1(n1454), .B0(n1453), .Y(n1455) );
  OA21A1OI2_X1M_A12TR u1255 ( .A0(n142), .A1(n1454), .B0(n212), .C0(n141), .Y(
        n1453) );
  AOI21_X1M_A12TR u1256 ( .A0(n141), .A1(n1452), .B0(n1451), .Y(n1456) );
  OA21A1OI2_X1M_A12TR u1257 ( .A0(n219), .A1(n1478), .B0(n1477), .C0(reset), 
        .Y(s0m_o0sm_n38) );
  OAI21_X1M_A12TR u1258 ( .A0(n219), .A1(n1476), .B0(n1475), .Y(n1477) );
  OA21A1OI2_X1M_A12TR u1259 ( .A0(n75), .A1(n1476), .B0(n219), .C0(n74), .Y(
        n1475) );
  AOI21_X1M_A12TR u1260 ( .A0(n74), .A1(n1474), .B0(n1473), .Y(n1478) );
  OAI222_X1M_A12TR u1261 ( .A0(n1196), .A1(n121), .B0(n1195), .B1(n1227), .C0(
        n1194), .C1(n1225), .Y(n922) );
  OAI222_X1M_A12TR u1262 ( .A0(n1196), .A1(n116), .B0(n1195), .B1(n1224), .C0(
        n1194), .C1(n1223), .Y(n923) );
  OAI222_X1M_A12TR u1263 ( .A0(n1196), .A1(n111), .B0(n1195), .B1(n1222), .C0(
        n1194), .C1(n1221), .Y(n924) );
  OAI222_X1M_A12TR u1264 ( .A0(n1196), .A1(n106), .B0(n1195), .B1(n1220), .C0(
        n1194), .C1(n1219), .Y(n925) );
  OAI222_X1M_A12TR u1265 ( .A0(n1229), .A1(n82), .B0(n1228), .B1(n1208), .C0(
        n1226), .C1(n1207), .Y(n919) );
  OAI222_X1M_A12TR u1266 ( .A0(n1375), .A1(n62), .B0(n1374), .B1(n1403), .C0(
        n1373), .C1(n1402), .Y(n854) );
  OAI222_X1M_A12TR u1267 ( .A0(n1375), .A1(n58), .B0(n1374), .B1(n1401), .C0(
        n1373), .C1(n1400), .Y(n855) );
  NAND3_X1M_A12TR u1268 ( .A(n72), .B(n1485), .C(n1486), .Y(x0m_n5) );
  AOI21_X1M_A12TR u1269 ( .A0(n147), .A1(n1070), .B0(n1069), .Y(n967) );
  OAI21_X1M_A12TR u1270 ( .A0(n147), .A1(n1070), .B0(n1485), .Y(n1069) );
  NAND2_X1M_A12TR u1271 ( .A(n1076), .B(n1346), .Y(n1070) );
  OAI221_X1M_A12TR u1272 ( .A0(n75), .A1(n1469), .B0(n1471), .B1(n1472), .C0(
        n1485), .Y(s0m_o0sm_n36) );
  OAI221_X1M_A12TR u1273 ( .A0(n142), .A1(n1447), .B0(n1449), .B1(n1450), .C0(
        n1485), .Y(s0m_o0nm_n36) );
  NAND3_X1M_A12TR u1274 ( .A(n10), .B(n1485), .C(n1483), .Y(x0m_n3) );
  AOI21_X1M_A12TR u1275 ( .A0(n150), .A1(n1068), .B0(n1067), .Y(n970) );
  OAI21_X1M_A12TR u1276 ( .A0(n150), .A1(n1068), .B0(n1485), .Y(n1067) );
  INV_X1M_A12TR u1277 ( .A(n1066), .Y(n1068) );
  AOI22_X1M_A12TR u1278 ( .A0(n66), .A1(n158), .B0(n1436), .B1(n1274), .Y(n890) );
  NAND2_X1M_A12TR u1279 ( .A(n1485), .B(n1411), .Y(n1436) );
  INV_X1M_A12TR u1280 ( .A(creditout_1), .Y(n158) );
  AOI22_X1M_A12TR u1281 ( .A0(n134), .A1(n168), .B0(n1268), .B1(n1087), .Y(
        n960) );
  NAND2_X1M_A12TR u1282 ( .A(n1485), .B(n1463), .Y(n1268) );
  INV_X1M_A12TR u1283 ( .A(creditout_0), .Y(n168) );
  AOI21_X1M_A12TR u1284 ( .A0(n67), .A1(n1045), .B0(n1043), .Y(c0sm_v0m_n61)
         );
  OAI21_X1M_A12TR u1285 ( .A0(n67), .A1(n1045), .B0(n1485), .Y(n1043) );
  AOI31_X1M_A12TR u1286 ( .A0(n1077), .A1(n1466), .A2(n70), .B0(n1047), .Y(
        n1045) );
  NAND2_X1M_A12TR u1287 ( .A(n1046), .B(n1044), .Y(n1051) );
  INV_X1M_A12TR u1288 ( .A(n67), .Y(n1044) );
  INV_X1M_A12TR u1289 ( .A(n69), .Y(n1046) );
  AOI22_X1M_A12TR u1290 ( .A0(n75), .A1(n1476), .B0(n1482), .B1(n1471), .Y(
        n1473) );
  INV_X1M_A12TR u1291 ( .A(n75), .Y(n1471) );
  INV_X1M_A12TR u1292 ( .A(n1470), .Y(n1482) );
  INV_X1M_A12TR u1293 ( .A(n1469), .Y(n1472) );
  NAND2_X1M_A12TR u1294 ( .A(n1474), .B(n1476), .Y(n1469) );
  NAND2_X1M_A12TR u1295 ( .A(creditin_1), .B(n1468), .Y(n1479) );
  NAND2_X1M_A12TR u1296 ( .A(n1470), .B(n1481), .Y(n1474) );
  NAND3_X1M_A12TR u1297 ( .A(n219), .B(n74), .C(n75), .Y(n1481) );
  NOR2_X1M_A12TR u1298 ( .A(creditin_1), .B(n1468), .Y(n1470) );
  AOI211_X1M_A12TR u1299 ( .A0(n1467), .A1(n1466), .B0(n1465), .C0(n1464), .Y(
        n1468) );
  AOI21_X1M_A12TR u1300 ( .A0(n79), .A1(n14), .B0(n1235), .Y(n1464) );
  NOR2_X1M_A12TR u1301 ( .A(n3), .B(n1463), .Y(n1465) );
  NOR2_X1M_A12TR u1302 ( .A(n2), .B(n1236), .Y(n1467) );
  INV_X1M_A12TR u1303 ( .A(n3), .Y(n1236) );
  AOI22_X1M_A12TR u1304 ( .A0(n142), .A1(n1454), .B0(n1460), .B1(n1449), .Y(
        n1451) );
  INV_X1M_A12TR u1305 ( .A(n142), .Y(n1449) );
  INV_X1M_A12TR u1306 ( .A(n1448), .Y(n1460) );
  INV_X1M_A12TR u1307 ( .A(n1447), .Y(n1450) );
  NAND2_X1M_A12TR u1308 ( .A(n1452), .B(n1454), .Y(n1447) );
  NAND2_X1M_A12TR u1309 ( .A(creditin_0), .B(n1446), .Y(n1457) );
  NAND2_X1M_A12TR u1310 ( .A(n1448), .B(n1459), .Y(n1452) );
  NAND3_X1M_A12TR u1311 ( .A(n212), .B(n141), .C(n142), .Y(n1459) );
  NOR2_X1M_A12TR u1312 ( .A(creditin_0), .B(n1446), .Y(n1448) );
  AOI211_X1M_A12TR u1313 ( .A0(n1445), .A1(n1466), .B0(n1444), .C0(n1443), .Y(
        n1446) );
  AOI21_X1M_A12TR u1314 ( .A0(n76), .A1(n11), .B0(n1269), .Y(n1443) );
  NOR2_X1M_A12TR u1315 ( .A(n1), .B(n1463), .Y(n1444) );
  NOR2_X1M_A12TR u1316 ( .A(n143), .B(n1271), .Y(n1445) );
  INV_X1M_A12TR u1317 ( .A(n1), .Y(n1271) );
  OAI22_X1M_A12TR u1318 ( .A0(n220), .A1(n1085), .B0(n11), .B1(n1084), .Y(n962) );
  OAI22_X1M_A12TR u1319 ( .A0(n221), .A1(n1085), .B0(n14), .B1(n1084), .Y(n965) );
  NOR2_X1M_A12TR u1320 ( .A(n1042), .B(n1083), .Y(n1081) );
  NAND2_X1M_A12TR u1321 ( .A(n1080), .B(n1082), .Y(n1085) );
  AOI211_X1M_A12TR u1322 ( .A0(n221), .A1(n220), .B0(n12), .C0(n13), .Y(n1082)
         );
  OAI222_X1M_A12TR u1323 ( .A0(n1355), .A1(n28), .B0(n1357), .B1(n1406), .C0(
        n1356), .C1(n1404), .Y(n966) );
  OAI222_X1M_A12TR u1324 ( .A0(n1375), .A1(n30), .B0(n1374), .B1(n1387), .C0(
        n1373), .C1(n1386), .Y(n862) );
  OAI222_X1M_A12TR u1325 ( .A0(n1375), .A1(n38), .B0(n1374), .B1(n1391), .C0(
        n1373), .C1(n1390), .Y(n860) );
  OAI222_X1M_A12TR u1326 ( .A0(n1375), .A1(n42), .B0(n1374), .B1(n1393), .C0(
        n1373), .C1(n1392), .Y(n859) );
  OAI222_X1M_A12TR u1327 ( .A0(n1375), .A1(n46), .B0(n1374), .B1(n1395), .C0(
        n1373), .C1(n1394), .Y(n858) );
  OAI222_X1M_A12TR u1328 ( .A0(n1375), .A1(n50), .B0(n1374), .B1(n1397), .C0(
        n1373), .C1(n1396), .Y(n857) );
  OAI222_X1M_A12TR u1329 ( .A0(n1196), .A1(n81), .B0(n1195), .B1(n1208), .C0(
        n1194), .C1(n1207), .Y(n931) );
  OAI222_X1M_A12TR u1330 ( .A0(n1196), .A1(n89), .B0(n1195), .B1(n1212), .C0(
        n1194), .C1(n1211), .Y(n929) );
  OAI222_X1M_A12TR u1331 ( .A0(n1196), .A1(n93), .B0(n1195), .B1(n1214), .C0(
        n1194), .C1(n1213), .Y(n928) );
  OAI222_X1M_A12TR u1332 ( .A0(n1196), .A1(n97), .B0(n1195), .B1(n1216), .C0(
        n1194), .C1(n1215), .Y(n927) );
  OAI222_X1M_A12TR u1333 ( .A0(n1196), .A1(n101), .B0(n1195), .B1(n1218), .C0(
        n1194), .C1(n1217), .Y(n926) );
  OAI222_X1M_A12TR u1334 ( .A0(n1357), .A1(n1399), .B0(n1356), .B1(n1398), 
        .C0(n1355), .C1(n56), .Y(n879) );
  OAI222_X1M_A12TR u1335 ( .A0(n1357), .A1(n1401), .B0(n1356), .B1(n1400), 
        .C0(n1355), .C1(n60), .Y(n878) );
  OAI222_X1M_A12TR u1336 ( .A0(n1357), .A1(n1403), .B0(n1356), .B1(n1402), 
        .C0(n1355), .C1(n64), .Y(n877) );
  OAI222_X1M_A12TR u1337 ( .A0(n1178), .A1(n1220), .B0(n1177), .B1(n1219), 
        .C0(n1176), .C1(n108), .Y(n949) );
  OAI222_X1M_A12TR u1338 ( .A0(n1178), .A1(n1222), .B0(n1177), .B1(n1221), 
        .C0(n1176), .C1(n113), .Y(n948) );
  OAI222_X1M_A12TR u1339 ( .A0(n1178), .A1(n1224), .B0(n1177), .B1(n1223), 
        .C0(n1176), .C1(n118), .Y(n947) );
  OAI222_X1M_A12TR u1340 ( .A0(n1178), .A1(n1227), .B0(n1177), .B1(n1225), 
        .C0(n1176), .C1(n123), .Y(n946) );
  OA21A1OI2_X1M_A12TR u1341 ( .A0(n1487), .A1(n1273), .B0(n10), .C0(n1083), 
        .Y(n963) );
  NOR2_X1M_A12TR u1342 ( .A(n11), .B(n1269), .Y(n1438) );
  INV_X1M_A12TR u1343 ( .A(s0m_elig_0_), .Y(n1269) );
  INV_X1M_A12TR u1344 ( .A(n76), .Y(n1239) );
  INV_X1M_A12TR u1345 ( .A(n72), .Y(n1487) );
  OA21A1OI2_X1M_A12TR u1346 ( .A0(n1484), .A1(n1238), .B0(n72), .C0(n1083), 
        .Y(n964) );
  INV_X1M_A12TR u1347 ( .A(n1080), .Y(n1083) );
  NOR2_X1M_A12TR u1348 ( .A(n14), .B(n1235), .Y(n1440) );
  INV_X1M_A12TR u1349 ( .A(s0m_elig_1_), .Y(n1235) );
  INV_X1M_A12TR u1350 ( .A(n79), .Y(n1086) );
  INV_X1M_A12TR u1351 ( .A(n10), .Y(n1484) );
  OAI222_X1M_A12TR u1352 ( .A0(n1408), .A1(n55), .B0(n1407), .B1(n1399), .C0(
        n1405), .C1(n1398), .Y(n844) );
  OAI222_X1M_A12TR u1353 ( .A0(n1408), .A1(n59), .B0(n1407), .B1(n1401), .C0(
        n1405), .C1(n1400), .Y(n843) );
  OAI222_X1M_A12TR u1354 ( .A0(n1408), .A1(n63), .B0(n1407), .B1(n1403), .C0(
        n1405), .C1(n1402), .Y(n842) );
  OAI222_X1M_A12TR u1355 ( .A0(n1176), .A1(n83), .B0(n1178), .B1(n1208), .C0(
        n1177), .C1(n1207), .Y(n955) );
  OAI222_X1M_A12TR u1356 ( .A0(n1229), .A1(n107), .B0(n1228), .B1(n1220), .C0(
        n1226), .C1(n1219), .Y(n913) );
  OAI222_X1M_A12TR u1357 ( .A0(n1229), .A1(n112), .B0(n1228), .B1(n1222), .C0(
        n1226), .C1(n1221), .Y(n912) );
  OAI222_X1M_A12TR u1358 ( .A0(n1229), .A1(n117), .B0(n1228), .B1(n1224), .C0(
        n1226), .C1(n1223), .Y(n911) );
  OAI222_X1M_A12TR u1359 ( .A0(n1229), .A1(n122), .B0(n1228), .B1(n1227), .C0(
        n1226), .C1(n1225), .Y(n910) );
  OAI222_X1M_A12TR u1360 ( .A0(n1366), .A1(n53), .B0(n1365), .B1(n1399), .C0(
        n1364), .C1(n1398), .Y(n868) );
  OAI222_X1M_A12TR u1361 ( .A0(n1366), .A1(n57), .B0(n1365), .B1(n1401), .C0(
        n1364), .C1(n1400), .Y(n867) );
  NOR2_X1M_A12TR u1362 ( .A(n1339), .B(n1338), .Y(n1400) );
  OAI22_X1M_A12TR u1363 ( .A0(n57), .A1(n1352), .B0(n58), .B1(n1351), .Y(n1338) );
  OAI21_X1M_A12TR u1364 ( .A0(n59), .A1(n1350), .B0(n1337), .Y(n1339) );
  AOI22_X1M_A12TR u1365 ( .A0(n1348), .A1(n1336), .B0(flitin_1[9]), .B1(n1346), 
        .Y(n1337) );
  INV_X1M_A12TR u1366 ( .A(n60), .Y(n1336) );
  NOR2_X1M_A12TR u1367 ( .A(n1335), .B(n1334), .Y(n1401) );
  OAI22_X1M_A12TR u1368 ( .A0(n59), .A1(n1343), .B0(n60), .B1(n1342), .Y(n1334) );
  OAI22_X1M_A12TR u1369 ( .A0(n57), .A1(n1341), .B0(n58), .B1(n1340), .Y(n1335) );
  OAI222_X1M_A12TR u1370 ( .A0(n1366), .A1(n61), .B0(n1365), .B1(n1403), .C0(
        n1364), .C1(n1402), .Y(n866) );
  NOR2_X1M_A12TR u1371 ( .A(n1354), .B(n1353), .Y(n1402) );
  OAI22_X1M_A12TR u1372 ( .A0(n61), .A1(n1352), .B0(n62), .B1(n1351), .Y(n1353) );
  OAI21_X1M_A12TR u1373 ( .A0(n63), .A1(n1350), .B0(n1349), .Y(n1354) );
  AOI22_X1M_A12TR u1374 ( .A0(n1348), .A1(n1347), .B0(flitin_1[10]), .B1(n1346), .Y(n1349) );
  INV_X1M_A12TR u1375 ( .A(n64), .Y(n1347) );
  NOR2_X1M_A12TR u1376 ( .A(n1345), .B(n1344), .Y(n1403) );
  OAI22_X1M_A12TR u1377 ( .A0(n63), .A1(n1343), .B0(n64), .B1(n1342), .Y(n1344) );
  OAI22_X1M_A12TR u1378 ( .A0(n61), .A1(n1341), .B0(n62), .B1(n1340), .Y(n1345) );
  AOI211_X1M_A12TR u1379 ( .A0(n151), .A1(n1090), .B0(reset), .C0(n1066), .Y(
        n971) );
  NOR2_X1M_A12TR u1380 ( .A(n151), .B(n1090), .Y(n1066) );
  OAI222_X1M_A12TR u1381 ( .A0(n1187), .A1(n105), .B0(n1186), .B1(n1220), .C0(
        n1185), .C1(n1219), .Y(n937) );
  NOR2_X1M_A12TR u1382 ( .A(n1148), .B(n1147), .Y(n1219) );
  OAI22_X1M_A12TR u1383 ( .A0(n105), .A1(n1173), .B0(n106), .B1(n1172), .Y(
        n1147) );
  OAI21_X1M_A12TR u1384 ( .A0(n107), .A1(n1171), .B0(n1146), .Y(n1148) );
  AOI22_X1M_A12TR u1385 ( .A0(n1169), .A1(n1145), .B0(flitin_0[8]), .B1(n1167), 
        .Y(n1146) );
  INV_X1M_A12TR u1386 ( .A(n108), .Y(n1145) );
  NOR2_X1M_A12TR u1387 ( .A(n1144), .B(n1143), .Y(n1220) );
  OAI22_X1M_A12TR u1388 ( .A0(n107), .A1(n1164), .B0(n108), .B1(n1163), .Y(
        n1143) );
  OAI22_X1M_A12TR u1389 ( .A0(n105), .A1(n1162), .B0(n106), .B1(n1161), .Y(
        n1144) );
  OAI222_X1M_A12TR u1390 ( .A0(n1187), .A1(n110), .B0(n1186), .B1(n1222), .C0(
        n1185), .C1(n1221), .Y(n936) );
  NOR2_X1M_A12TR u1391 ( .A(n1154), .B(n1153), .Y(n1221) );
  OAI22_X1M_A12TR u1392 ( .A0(n110), .A1(n1173), .B0(n111), .B1(n1172), .Y(
        n1153) );
  OAI21_X1M_A12TR u1393 ( .A0(n112), .A1(n1171), .B0(n1152), .Y(n1154) );
  AOI22_X1M_A12TR u1394 ( .A0(n1169), .A1(n1151), .B0(flitin_0[9]), .B1(n1167), 
        .Y(n1152) );
  INV_X1M_A12TR u1395 ( .A(n113), .Y(n1151) );
  NOR2_X1M_A12TR u1396 ( .A(n1150), .B(n1149), .Y(n1222) );
  OAI22_X1M_A12TR u1397 ( .A0(n112), .A1(n1164), .B0(n113), .B1(n1163), .Y(
        n1149) );
  OAI22_X1M_A12TR u1398 ( .A0(n110), .A1(n1162), .B0(n111), .B1(n1161), .Y(
        n1150) );
  OAI222_X1M_A12TR u1399 ( .A0(n1187), .A1(n115), .B0(n1186), .B1(n1224), .C0(
        n1185), .C1(n1223), .Y(n935) );
  NOR2_X1M_A12TR u1400 ( .A(n1160), .B(n1159), .Y(n1223) );
  OAI22_X1M_A12TR u1401 ( .A0(n115), .A1(n1173), .B0(n116), .B1(n1172), .Y(
        n1159) );
  OAI21_X1M_A12TR u1402 ( .A0(n117), .A1(n1171), .B0(n1158), .Y(n1160) );
  AOI22_X1M_A12TR u1403 ( .A0(n1169), .A1(n1157), .B0(flitin_0[10]), .B1(n1167), .Y(n1158) );
  INV_X1M_A12TR u1404 ( .A(n118), .Y(n1157) );
  NOR2_X1M_A12TR u1405 ( .A(n1156), .B(n1155), .Y(n1224) );
  OAI22_X1M_A12TR u1406 ( .A0(n117), .A1(n1164), .B0(n118), .B1(n1163), .Y(
        n1155) );
  OAI22_X1M_A12TR u1407 ( .A0(n115), .A1(n1162), .B0(n116), .B1(n1161), .Y(
        n1156) );
  OAI222_X1M_A12TR u1408 ( .A0(n1187), .A1(n120), .B0(n1186), .B1(n1227), .C0(
        n1185), .C1(n1225), .Y(n934) );
  NOR2_X1M_A12TR u1409 ( .A(n1175), .B(n1174), .Y(n1225) );
  OAI22_X1M_A12TR u1410 ( .A0(n120), .A1(n1173), .B0(n121), .B1(n1172), .Y(
        n1174) );
  OAI21_X1M_A12TR u1411 ( .A0(n122), .A1(n1171), .B0(n1170), .Y(n1175) );
  AOI22_X1M_A12TR u1412 ( .A0(n1169), .A1(n1168), .B0(flitin_0[11]), .B1(n1167), .Y(n1170) );
  INV_X1M_A12TR u1413 ( .A(n123), .Y(n1168) );
  NOR2_X1M_A12TR u1414 ( .A(n1166), .B(n1165), .Y(n1227) );
  OAI22_X1M_A12TR u1415 ( .A0(n122), .A1(n1164), .B0(n123), .B1(n1163), .Y(
        n1165) );
  OAI22_X1M_A12TR u1416 ( .A0(n120), .A1(n1162), .B0(n121), .B1(n1161), .Y(
        n1166) );
  OAI222_X1M_A12TR u1417 ( .A0(n1408), .A1(n27), .B0(n1407), .B1(n1406), .C0(
        n1405), .C1(n1404), .Y(n841) );
  OAI21_X1M_A12TR u1418 ( .A0(n12), .A1(n1041), .B0(n1080), .Y(c0sm_v0m_n57)
         );
  NOR2_X1M_A12TR u1419 ( .A(reset), .B(tailout_1), .Y(n1080) );
  OAI222_X1M_A12TR u1420 ( .A0(n1375), .A1(n26), .B0(n1374), .B1(n1406), .C0(
        n1373), .C1(n1404), .Y(n853) );
  OAI222_X1M_A12TR u1421 ( .A0(n1366), .A1(n29), .B0(n1365), .B1(n1387), .C0(
        n1364), .C1(n1386), .Y(n874) );
  OAI222_X1M_A12TR u1422 ( .A0(n1375), .A1(n34), .B0(n1374), .B1(n1389), .C0(
        n1373), .C1(n1388), .Y(n861) );
  OAI222_X1M_A12TR u1423 ( .A0(n1408), .A1(n43), .B0(n1407), .B1(n1393), .C0(
        n1405), .C1(n1392), .Y(n847) );
  OAI222_X1M_A12TR u1424 ( .A0(n1408), .A1(n47), .B0(n1407), .B1(n1395), .C0(
        n1405), .C1(n1394), .Y(n846) );
  OAI222_X1M_A12TR u1425 ( .A0(n1408), .A1(n51), .B0(n1407), .B1(n1397), .C0(
        n1405), .C1(n1396), .Y(n845) );
  OAI222_X1M_A12TR u1426 ( .A0(n1187), .A1(n80), .B0(n1186), .B1(n1208), .C0(
        n1185), .C1(n1207), .Y(n943) );
  AOI211_X1M_A12TR u1427 ( .A0(n1142), .A1(n1109), .B0(n1108), .C0(n1107), .Y(
        n1207) );
  OAI22_X1M_A12TR u1428 ( .A0(n80), .A1(n1173), .B0(n82), .B1(n1171), .Y(n1107) );
  OAI21_X1M_A12TR u1429 ( .A0(n83), .A1(n1138), .B0(n1106), .Y(n1108) );
  NAND2_X1M_A12TR u1430 ( .A(flitin_0[2]), .B(n1167), .Y(n1106) );
  INV_X1M_A12TR u1431 ( .A(n81), .Y(n1109) );
  NOR2_X1M_A12TR u1432 ( .A(n1104), .B(n1103), .Y(n1208) );
  OAI22_X1M_A12TR u1433 ( .A0(n83), .A1(n1163), .B0(n82), .B1(n1164), .Y(n1103) );
  OAI22_X1M_A12TR u1434 ( .A0(n80), .A1(n1162), .B0(n81), .B1(n1161), .Y(n1104) );
  OAI222_X1M_A12TR u1435 ( .A0(n1196), .A1(n85), .B0(n1195), .B1(n1210), .C0(
        n1194), .C1(n1209), .Y(n930) );
  NAND2_X1M_A12TR u1436 ( .A(n1193), .B(n1485), .Y(n1194) );
  INV_X1M_A12TR u1437 ( .A(n1191), .Y(n1193) );
  NAND3_X1M_A12TR u1438 ( .A(n1192), .B(n1485), .C(n1191), .Y(n1195) );
  NAND3_X1M_A12TR u1439 ( .A(n1485), .B(n1263), .C(n1191), .Y(n1196) );
  OAI222_X1M_A12TR u1440 ( .A0(n1229), .A1(n94), .B0(n1228), .B1(n1214), .C0(
        n1226), .C1(n1213), .Y(n916) );
  OAI222_X1M_A12TR u1441 ( .A0(n1229), .A1(n98), .B0(n1228), .B1(n1216), .C0(
        n1226), .C1(n1215), .Y(n915) );
  OAI222_X1M_A12TR u1442 ( .A0(n1229), .A1(n102), .B0(n1228), .B1(n1218), .C0(
        n1226), .C1(n1217), .Y(n914) );
  OAI222_X1M_A12TR u1443 ( .A0(n1357), .A1(n1387), .B0(n1355), .B1(n32), .C0(
        n1356), .C1(n1386), .Y(n885) );
  OAI222_X1M_A12TR u1444 ( .A0(n1357), .A1(n1389), .B0(n1355), .B1(n36), .C0(
        n1356), .C1(n1388), .Y(n884) );
  OAI222_X1M_A12TR u1445 ( .A0(n1357), .A1(n1391), .B0(n1355), .B1(n40), .C0(
        n1356), .C1(n1390), .Y(n883) );
  OAI222_X1M_A12TR u1446 ( .A0(n1178), .A1(n1210), .B0(n1176), .B1(n87), .C0(
        n1177), .C1(n1209), .Y(n954) );
  OAI222_X1M_A12TR u1447 ( .A0(n1178), .A1(n1212), .B0(n1176), .B1(n91), .C0(
        n1177), .C1(n1211), .Y(n953) );
  OAI222_X1M_A12TR u1448 ( .A0(n1366), .A1(n33), .B0(n1365), .B1(n1389), .C0(
        n1364), .C1(n1388), .Y(n873) );
  AOI211_X1M_A12TR u1449 ( .A0(n1301), .A1(n1300), .B0(n1299), .C0(n1298), .Y(
        n1388) );
  OAI22_X1M_A12TR u1450 ( .A0(n34), .A1(n1351), .B0(n33), .B1(n1352), .Y(n1298) );
  OAI21_X1M_A12TR u1451 ( .A0(n36), .A1(n1323), .B0(n1297), .Y(n1299) );
  NAND2_X1M_A12TR u1452 ( .A(flitin_1[3]), .B(n1346), .Y(n1297) );
  INV_X1M_A12TR u1453 ( .A(n35), .Y(n1300) );
  INV_X1M_A12TR u1454 ( .A(n1350), .Y(n1301) );
  NOR2_X1M_A12TR u1455 ( .A(n1296), .B(n1295), .Y(n1389) );
  OAI22_X1M_A12TR u1456 ( .A0(n36), .A1(n1342), .B0(n35), .B1(n1343), .Y(n1295) );
  OAI22_X1M_A12TR u1457 ( .A0(n34), .A1(n1340), .B0(n33), .B1(n1341), .Y(n1296) );
  OAI222_X1M_A12TR u1458 ( .A0(n1187), .A1(n84), .B0(n1186), .B1(n1210), .C0(
        n1185), .C1(n1209), .Y(n942) );
  AOI211_X1M_A12TR u1459 ( .A0(n1116), .A1(n1115), .B0(n1114), .C0(n1113), .Y(
        n1209) );
  OAI22_X1M_A12TR u1460 ( .A0(n85), .A1(n1172), .B0(n84), .B1(n1173), .Y(n1113) );
  INV_X1M_A12TR u1461 ( .A(n1142), .Y(n1172) );
  OAI21_X1M_A12TR u1462 ( .A0(n87), .A1(n1138), .B0(n1112), .Y(n1114) );
  NAND2_X1M_A12TR u1463 ( .A(flitin_0[3]), .B(n1167), .Y(n1112) );
  INV_X1M_A12TR u1464 ( .A(n86), .Y(n1115) );
  NOR2_X1M_A12TR u1465 ( .A(n1111), .B(n1110), .Y(n1210) );
  OAI22_X1M_A12TR u1466 ( .A0(n87), .A1(n1163), .B0(n86), .B1(n1164), .Y(n1110) );
  OAI22_X1M_A12TR u1467 ( .A0(n85), .A1(n1161), .B0(n84), .B1(n1162), .Y(n1111) );
  OAI222_X1M_A12TR u1468 ( .A0(n1366), .A1(n25), .B0(n1365), .B1(n1406), .C0(
        n1364), .C1(n1404), .Y(n865) );
  NOR2_X1M_A12TR u1469 ( .A(n1079), .B(n1078), .Y(n1404) );
  OAI22_X1M_A12TR u1470 ( .A0(n26), .A1(n1351), .B0(n25), .B1(n1352), .Y(n1078) );
  OAI21_X1M_A12TR u1471 ( .A0(n27), .A1(n1350), .B0(n1075), .Y(n1079) );
  AOI22_X1M_A12TR u1472 ( .A0(flitin_1[11]), .A1(n1346), .B0(n1348), .B1(n1074), .Y(n1075) );
  INV_X1M_A12TR u1473 ( .A(n28), .Y(n1074) );
  NOR2_X1M_A12TR u1474 ( .A(n1073), .B(n1072), .Y(n1406) );
  OAI22_X1M_A12TR u1475 ( .A0(n28), .A1(n1342), .B0(n27), .B1(n1343), .Y(n1072) );
  OAI22_X1M_A12TR u1476 ( .A0(n26), .A1(n1340), .B0(n25), .B1(n1341), .Y(n1073) );
  OAI222_X1M_A12TR u1477 ( .A0(n1366), .A1(n37), .B0(n1365), .B1(n1391), .C0(
        n1364), .C1(n1390), .Y(n872) );
  OAI222_X1M_A12TR u1478 ( .A0(n1408), .A1(n39), .B0(n1407), .B1(n1391), .C0(
        n1405), .C1(n1390), .Y(n848) );
  AOI211_X1M_A12TR u1479 ( .A0(n1327), .A1(n1307), .B0(n1306), .C0(n1305), .Y(
        n1390) );
  OAI22_X1M_A12TR u1480 ( .A0(n39), .A1(n1350), .B0(n37), .B1(n1352), .Y(n1305) );
  OAI21_X1M_A12TR u1481 ( .A0(n40), .A1(n1323), .B0(n1304), .Y(n1306) );
  NAND2_X1M_A12TR u1482 ( .A(flitin_1[4]), .B(n1346), .Y(n1304) );
  INV_X1M_A12TR u1483 ( .A(n38), .Y(n1307) );
  NOR2_X1M_A12TR u1484 ( .A(n1303), .B(n1302), .Y(n1391) );
  OAI22_X1M_A12TR u1485 ( .A0(n40), .A1(n1342), .B0(n39), .B1(n1343), .Y(n1302) );
  OAI22_X1M_A12TR u1486 ( .A0(n38), .A1(n1340), .B0(n37), .B1(n1341), .Y(n1303) );
  OAI222_X1M_A12TR u1487 ( .A0(n1366), .A1(n41), .B0(n1365), .B1(n1393), .C0(
        n1364), .C1(n1392), .Y(n871) );
  OAI222_X1M_A12TR u1488 ( .A0(n1366), .A1(n45), .B0(n1365), .B1(n1395), .C0(
        n1364), .C1(n1394), .Y(n870) );
  OAI222_X1M_A12TR u1489 ( .A0(n1366), .A1(n49), .B0(n1365), .B1(n1397), .C0(
        n1364), .C1(n1396), .Y(n869) );
  NAND2_X1M_A12TR u1490 ( .A(n1363), .B(n1485), .Y(n1364) );
  NAND3_X1M_A12TR u1491 ( .A(n1362), .B(n1485), .C(n1361), .Y(n1365) );
  NAND3_X1M_A12TR u1492 ( .A(n1485), .B(n1432), .C(n1361), .Y(n1366) );
  INV_X1M_A12TR u1493 ( .A(n1363), .Y(n1361) );
  OAI222_X1M_A12TR u1494 ( .A0(n1187), .A1(n88), .B0(n1186), .B1(n1212), .C0(
        n1185), .C1(n1211), .Y(n941) );
  OAI222_X1M_A12TR u1495 ( .A0(n1229), .A1(n90), .B0(n1228), .B1(n1212), .C0(
        n1226), .C1(n1211), .Y(n917) );
  AOI211_X1M_A12TR u1496 ( .A0(n1142), .A1(n1122), .B0(n1121), .C0(n1120), .Y(
        n1211) );
  OAI22_X1M_A12TR u1497 ( .A0(n90), .A1(n1171), .B0(n88), .B1(n1173), .Y(n1120) );
  OAI21_X1M_A12TR u1498 ( .A0(n91), .A1(n1138), .B0(n1119), .Y(n1121) );
  NAND2_X1M_A12TR u1499 ( .A(flitin_0[4]), .B(n1167), .Y(n1119) );
  INV_X1M_A12TR u1500 ( .A(n89), .Y(n1122) );
  NAND2_X1M_A12TR u1501 ( .A(n1206), .B(n1485), .Y(n1226) );
  NOR2_X1M_A12TR u1502 ( .A(n1118), .B(n1117), .Y(n1212) );
  OAI22_X1M_A12TR u1503 ( .A0(n91), .A1(n1163), .B0(n90), .B1(n1164), .Y(n1117) );
  OAI22_X1M_A12TR u1504 ( .A0(n89), .A1(n1161), .B0(n88), .B1(n1162), .Y(n1118) );
  NAND3_X1M_A12TR u1505 ( .A(n1205), .B(n1485), .C(n1204), .Y(n1228) );
  NAND3_X1M_A12TR u1506 ( .A(n1485), .B(n1262), .C(n1204), .Y(n1229) );
  OAI222_X1M_A12TR u1507 ( .A0(n1187), .A1(n92), .B0(n1186), .B1(n1214), .C0(
        n1185), .C1(n1213), .Y(n940) );
  OAI222_X1M_A12TR u1508 ( .A0(n1187), .A1(n96), .B0(n1186), .B1(n1216), .C0(
        n1185), .C1(n1215), .Y(n939) );
  OAI222_X1M_A12TR u1509 ( .A0(n1187), .A1(n100), .B0(n1186), .B1(n1218), .C0(
        n1185), .C1(n1217), .Y(n938) );
  NAND2_X1M_A12TR u1510 ( .A(n1184), .B(n1485), .Y(n1185) );
  NAND3_X1M_A12TR u1511 ( .A(n1183), .B(n1485), .C(n1182), .Y(n1186) );
  NAND3_X1M_A12TR u1512 ( .A(n1485), .B(n1264), .C(n1182), .Y(n1187) );
  INV_X1M_A12TR u1513 ( .A(n1184), .Y(n1182) );
  OAI222_X1M_A12TR u1514 ( .A0(n1357), .A1(n1393), .B0(n1355), .B1(n44), .C0(
        n1356), .C1(n1392), .Y(n882) );
  AOI211_X1M_A12TR u1515 ( .A0(n1327), .A1(n1313), .B0(n1312), .C0(n1311), .Y(
        n1392) );
  OAI22_X1M_A12TR u1516 ( .A0(n43), .A1(n1350), .B0(n41), .B1(n1352), .Y(n1311) );
  OAI21_X1M_A12TR u1517 ( .A0(n44), .A1(n1323), .B0(n1310), .Y(n1312) );
  NAND2_X1M_A12TR u1518 ( .A(flitin_1[5]), .B(n1346), .Y(n1310) );
  INV_X1M_A12TR u1519 ( .A(n42), .Y(n1313) );
  NOR2_X1M_A12TR u1520 ( .A(n1309), .B(n1308), .Y(n1393) );
  OAI22_X1M_A12TR u1521 ( .A0(n44), .A1(n1342), .B0(n43), .B1(n1343), .Y(n1308) );
  OAI22_X1M_A12TR u1522 ( .A0(n41), .A1(n1341), .B0(n42), .B1(n1340), .Y(n1309) );
  OAI222_X1M_A12TR u1523 ( .A0(n1357), .A1(n1395), .B0(n1355), .B1(n48), .C0(
        n1356), .C1(n1394), .Y(n881) );
  AOI211_X1M_A12TR u1524 ( .A0(n1327), .A1(n1319), .B0(n1318), .C0(n1317), .Y(
        n1394) );
  OAI22_X1M_A12TR u1525 ( .A0(n47), .A1(n1350), .B0(n45), .B1(n1352), .Y(n1317) );
  OAI21_X1M_A12TR u1526 ( .A0(n48), .A1(n1323), .B0(n1316), .Y(n1318) );
  NAND2_X1M_A12TR u1527 ( .A(flitin_1[6]), .B(n1346), .Y(n1316) );
  INV_X1M_A12TR u1528 ( .A(n46), .Y(n1319) );
  NOR2_X1M_A12TR u1529 ( .A(n1315), .B(n1314), .Y(n1395) );
  OAI22_X1M_A12TR u1530 ( .A0(n48), .A1(n1342), .B0(n47), .B1(n1343), .Y(n1314) );
  OAI22_X1M_A12TR u1531 ( .A0(n45), .A1(n1341), .B0(n46), .B1(n1340), .Y(n1315) );
  OAI222_X1M_A12TR u1532 ( .A0(n1357), .A1(n1397), .B0(n1355), .B1(n52), .C0(
        n1356), .C1(n1396), .Y(n880) );
  AOI211_X1M_A12TR u1533 ( .A0(n1327), .A1(n1326), .B0(n1325), .C0(n1324), .Y(
        n1396) );
  OAI22_X1M_A12TR u1534 ( .A0(n51), .A1(n1350), .B0(n49), .B1(n1352), .Y(n1324) );
  OAI21_X1M_A12TR u1535 ( .A0(n52), .A1(n1323), .B0(n1322), .Y(n1325) );
  NAND2_X1M_A12TR u1536 ( .A(flitin_1[7]), .B(n1346), .Y(n1322) );
  INV_X1M_A12TR u1537 ( .A(n50), .Y(n1326) );
  NAND2_X1M_A12TR u1538 ( .A(n1286), .B(n1485), .Y(n1356) );
  INV_X1M_A12TR u1539 ( .A(n1285), .Y(n1286) );
  NAND3_X1M_A12TR u1540 ( .A(n1485), .B(n1429), .C(n1285), .Y(n1355) );
  NOR2_X1M_A12TR u1541 ( .A(n1321), .B(n1320), .Y(n1397) );
  OAI22_X1M_A12TR u1542 ( .A0(n52), .A1(n1342), .B0(n51), .B1(n1343), .Y(n1320) );
  OAI22_X1M_A12TR u1543 ( .A0(n49), .A1(n1341), .B0(n50), .B1(n1340), .Y(n1321) );
  NAND3_X1M_A12TR u1544 ( .A(n1071), .B(n1485), .C(n1285), .Y(n1357) );
  OAI222_X1M_A12TR u1545 ( .A0(n1178), .A1(n1214), .B0(n1176), .B1(n95), .C0(
        n1177), .C1(n1213), .Y(n952) );
  AOI211_X1M_A12TR u1546 ( .A0(n1142), .A1(n1128), .B0(n1127), .C0(n1126), .Y(
        n1213) );
  OAI22_X1M_A12TR u1547 ( .A0(n94), .A1(n1171), .B0(n92), .B1(n1173), .Y(n1126) );
  OAI21_X1M_A12TR u1548 ( .A0(n95), .A1(n1138), .B0(n1125), .Y(n1127) );
  NAND2_X1M_A12TR u1549 ( .A(flitin_0[5]), .B(n1167), .Y(n1125) );
  INV_X1M_A12TR u1550 ( .A(n93), .Y(n1128) );
  NOR2_X1M_A12TR u1551 ( .A(n1124), .B(n1123), .Y(n1214) );
  OAI22_X1M_A12TR u1552 ( .A0(n95), .A1(n1163), .B0(n94), .B1(n1164), .Y(n1123) );
  OAI22_X1M_A12TR u1553 ( .A0(n92), .A1(n1162), .B0(n93), .B1(n1161), .Y(n1124) );
  OAI222_X1M_A12TR u1554 ( .A0(n1178), .A1(n1216), .B0(n1176), .B1(n99), .C0(
        n1177), .C1(n1215), .Y(n951) );
  AOI211_X1M_A12TR u1555 ( .A0(n1142), .A1(n1134), .B0(n1133), .C0(n1132), .Y(
        n1215) );
  OAI22_X1M_A12TR u1556 ( .A0(n98), .A1(n1171), .B0(n96), .B1(n1173), .Y(n1132) );
  OAI21_X1M_A12TR u1557 ( .A0(n99), .A1(n1138), .B0(n1131), .Y(n1133) );
  NAND2_X1M_A12TR u1558 ( .A(flitin_0[6]), .B(n1167), .Y(n1131) );
  INV_X1M_A12TR u1559 ( .A(n97), .Y(n1134) );
  NOR2_X1M_A12TR u1560 ( .A(n1130), .B(n1129), .Y(n1216) );
  OAI22_X1M_A12TR u1561 ( .A0(n99), .A1(n1163), .B0(n98), .B1(n1164), .Y(n1129) );
  OAI22_X1M_A12TR u1562 ( .A0(n96), .A1(n1162), .B0(n97), .B1(n1161), .Y(n1130) );
  OAI222_X1M_A12TR u1563 ( .A0(n1178), .A1(n1218), .B0(n1176), .B1(n103), .C0(
        n1177), .C1(n1217), .Y(n950) );
  AOI211_X1M_A12TR u1564 ( .A0(n1142), .A1(n1141), .B0(n1140), .C0(n1139), .Y(
        n1217) );
  OAI22_X1M_A12TR u1565 ( .A0(n102), .A1(n1171), .B0(n100), .B1(n1173), .Y(
        n1139) );
  NAND2_X1M_A12TR u1566 ( .A(n1090), .B(n1184), .Y(n1173) );
  NOR2_X1M_A12TR u1567 ( .A(n151), .B(n150), .Y(n1184) );
  INV_X1M_A12TR u1568 ( .A(n1167), .Y(n1090) );
  INV_X1M_A12TR u1569 ( .A(n1116), .Y(n1171) );
  NOR2_X1M_A12TR u1570 ( .A(n1167), .B(n1204), .Y(n1116) );
  INV_X1M_A12TR u1571 ( .A(n1206), .Y(n1204) );
  NOR2_X1M_A12TR u1572 ( .A(n1092), .B(n151), .Y(n1206) );
  OAI21_X1M_A12TR u1573 ( .A0(n103), .A1(n1138), .B0(n1137), .Y(n1140) );
  NAND2_X1M_A12TR u1574 ( .A(flitin_0[7]), .B(n1167), .Y(n1137) );
  INV_X1M_A12TR u1575 ( .A(n1169), .Y(n1138) );
  NOR2_X1M_A12TR u1576 ( .A(n1102), .B(n1167), .Y(n1169) );
  INV_X1M_A12TR u1577 ( .A(n101), .Y(n1141) );
  NOR2_X1M_A12TR u1578 ( .A(n1167), .B(n1191), .Y(n1142) );
  NAND2_X1M_A12TR u1579 ( .A(n151), .B(n1092), .Y(n1191) );
  INV_X1M_A12TR u1580 ( .A(n150), .Y(n1092) );
  NAND2_X1M_A12TR u1581 ( .A(flitin_0[0]), .B(flitin_0[1]), .Y(n1167) );
  NAND2_X1M_A12TR u1582 ( .A(n1105), .B(n1485), .Y(n1177) );
  INV_X1M_A12TR u1583 ( .A(n1102), .Y(n1105) );
  NOR2_X1M_A12TR u1584 ( .A(n1136), .B(n1135), .Y(n1218) );
  OAI22_X1M_A12TR u1585 ( .A0(n103), .A1(n1163), .B0(n102), .B1(n1164), .Y(
        n1135) );
  NAND2_X1M_A12TR u1586 ( .A(n1205), .B(n1463), .Y(n1164) );
  INV_X1M_A12TR u1587 ( .A(n1262), .Y(n1205) );
  NAND2_X1M_A12TR u1588 ( .A(n1089), .B(n1087), .Y(n1262) );
  OAI22_X1M_A12TR u1589 ( .A0(n100), .A1(n1162), .B0(n101), .B1(n1161), .Y(
        n1136) );
  NAND2_X1M_A12TR u1590 ( .A(n1192), .B(n1463), .Y(n1161) );
  INV_X1M_A12TR u1591 ( .A(n1263), .Y(n1192) );
  NAND2_X1M_A12TR u1592 ( .A(c0nm_b0m_v0m_head_1_), .B(n134), .Y(n1263) );
  NAND2_X1M_A12TR u1593 ( .A(n1183), .B(n1463), .Y(n1162) );
  INV_X1M_A12TR u1594 ( .A(n1264), .Y(n1183) );
  NAND2_X1M_A12TR u1595 ( .A(c0nm_b0m_v0m_head_1_), .B(n1087), .Y(n1264) );
  INV_X1M_A12TR u1596 ( .A(n134), .Y(n1087) );
  NAND3_X1M_A12TR u1597 ( .A(n1485), .B(n1102), .C(n1176), .Y(n1178) );
  NAND3_X1M_A12TR u1598 ( .A(n1485), .B(n1261), .C(n1102), .Y(n1176) );
  NAND2_X1M_A12TR u1599 ( .A(n134), .B(n1089), .Y(n1261) );
  INV_X1M_A12TR u1600 ( .A(c0nm_b0m_v0m_head_1_), .Y(n1089) );
  NAND2_X1M_A12TR u1601 ( .A(n151), .B(n150), .Y(n1102) );
  OAI222_X1M_A12TR u1602 ( .A0(n1408), .A1(n31), .B0(n1407), .B1(n1387), .C0(
        n1405), .C1(n1386), .Y(n850) );
  AOI211_X1M_A12TR u1603 ( .A0(n1327), .A1(n1294), .B0(n1293), .C0(n1292), .Y(
        n1386) );
  OAI22_X1M_A12TR u1604 ( .A0(n29), .A1(n1352), .B0(n31), .B1(n1350), .Y(n1292) );
  OAI21_X1M_A12TR u1605 ( .A0(n32), .A1(n1323), .B0(n1291), .Y(n1293) );
  NAND2_X1M_A12TR u1606 ( .A(flitin_1[2]), .B(n1346), .Y(n1291) );
  INV_X1M_A12TR u1607 ( .A(n1348), .Y(n1323) );
  INV_X1M_A12TR u1608 ( .A(n30), .Y(n1294) );
  INV_X1M_A12TR u1609 ( .A(n1351), .Y(n1327) );
  NAND2_X1M_A12TR u1610 ( .A(n1385), .B(n1485), .Y(n1405) );
  NOR2_X1M_A12TR u1611 ( .A(n1290), .B(n1289), .Y(n1387) );
  OAI22_X1M_A12TR u1612 ( .A0(n32), .A1(n1342), .B0(n31), .B1(n1343), .Y(n1289) );
  OAI22_X1M_A12TR u1613 ( .A0(n29), .A1(n1341), .B0(n30), .B1(n1340), .Y(n1290) );
  NAND3_X1M_A12TR u1614 ( .A(n1384), .B(n1485), .C(n1383), .Y(n1407) );
  NAND3_X1M_A12TR u1615 ( .A(n1485), .B(n1430), .C(n1383), .Y(n1408) );
  OAI222_X1M_A12TR u1616 ( .A0(n1375), .A1(n54), .B0(n1374), .B1(n1399), .C0(
        n1373), .C1(n1398), .Y(n856) );
  NOR2_X1M_A12TR u1617 ( .A(n1333), .B(n1332), .Y(n1398) );
  OAI22_X1M_A12TR u1618 ( .A0(n53), .A1(n1352), .B0(n54), .B1(n1351), .Y(n1332) );
  NAND2_X1M_A12TR u1619 ( .A(n1077), .B(n1372), .Y(n1351) );
  NAND2_X1M_A12TR u1620 ( .A(n1077), .B(n1363), .Y(n1352) );
  NOR2_X1M_A12TR u1621 ( .A(n148), .B(n147), .Y(n1363) );
  OAI21_X1M_A12TR u1622 ( .A0(n55), .A1(n1350), .B0(n1331), .Y(n1333) );
  AOI22_X1M_A12TR u1623 ( .A0(n1348), .A1(n1330), .B0(flitin_1[8]), .B1(n1346), 
        .Y(n1331) );
  INV_X1M_A12TR u1624 ( .A(n56), .Y(n1330) );
  NOR2_X1M_A12TR u1625 ( .A(n1285), .B(n1346), .Y(n1348) );
  NAND2_X1M_A12TR u1626 ( .A(n148), .B(n147), .Y(n1285) );
  NAND2_X1M_A12TR u1627 ( .A(n1077), .B(n1385), .Y(n1350) );
  INV_X1M_A12TR u1628 ( .A(n1383), .Y(n1385) );
  NAND2_X1M_A12TR u1629 ( .A(n1076), .B(n147), .Y(n1383) );
  NAND2_X1M_A12TR u1630 ( .A(flitin_1[0]), .B(flitin_1[1]), .Y(n1346) );
  NAND2_X1M_A12TR u1631 ( .A(n1372), .B(n1485), .Y(n1373) );
  NOR2_X1M_A12TR u1632 ( .A(n1329), .B(n1328), .Y(n1399) );
  OAI22_X1M_A12TR u1633 ( .A0(n55), .A1(n1343), .B0(n56), .B1(n1342), .Y(n1328) );
  NAND2_X1M_A12TR u1634 ( .A(n1071), .B(n1411), .Y(n1342) );
  INV_X1M_A12TR u1635 ( .A(n1429), .Y(n1071) );
  NAND2_X1M_A12TR u1636 ( .A(n66), .B(n1276), .Y(n1429) );
  NAND2_X1M_A12TR u1637 ( .A(n1384), .B(n1411), .Y(n1343) );
  INV_X1M_A12TR u1638 ( .A(n1430), .Y(n1384) );
  NAND2_X1M_A12TR u1639 ( .A(n1276), .B(n1274), .Y(n1430) );
  INV_X1M_A12TR u1640 ( .A(c0sm_b0m_v0m_head_1_), .Y(n1276) );
  OAI22_X1M_A12TR u1641 ( .A0(n53), .A1(n1341), .B0(n54), .B1(n1340), .Y(n1329) );
  NAND2_X1M_A12TR u1642 ( .A(n1371), .B(n1411), .Y(n1340) );
  NAND2_X1M_A12TR u1643 ( .A(n1362), .B(n1411), .Y(n1341) );
  INV_X1M_A12TR u1644 ( .A(n1432), .Y(n1362) );
  NAND2_X1M_A12TR u1645 ( .A(c0sm_b0m_v0m_head_1_), .B(n1274), .Y(n1432) );
  INV_X1M_A12TR u1646 ( .A(n66), .Y(n1274) );
  NAND3_X1M_A12TR u1647 ( .A(n1371), .B(n1485), .C(n1370), .Y(n1374) );
  INV_X1M_A12TR u1648 ( .A(n1431), .Y(n1371) );
  NAND3_X1M_A12TR u1649 ( .A(n1485), .B(n1431), .C(n1370), .Y(n1375) );
  INV_X1M_A12TR u1650 ( .A(n1372), .Y(n1370) );
  NOR2_X1M_A12TR u1651 ( .A(n147), .B(n1076), .Y(n1372) );
  NAND2_X1M_A12TR u1652 ( .A(c0sm_b0m_v0m_head_1_), .B(n66), .Y(n1431) );
  NOR2_X1M_A12TR u1653 ( .A(reset), .B(n1411), .Y(creditout_1) );
  AOI21_X1M_A12TR u1654 ( .A0(n69), .A1(n67), .B0(n1021), .Y(n1466) );
  AOI31_X1M_A12TR u1655 ( .A0(n12), .A1(n1020), .A2(n1019), .B0(n1042), .Y(
        n1021) );
  AOI21_X1M_A12TR u1656 ( .A0(n72), .A1(n10), .B0(n1020), .Y(n1041) );
  INV_X1M_A12TR u1657 ( .A(tailout_1), .Y(n1019) );
  INV_X1M_A12TR u1658 ( .A(n13), .Y(n1020) );
  NOR2_X1M_A12TR u1659 ( .A(reset), .B(n1463), .Y(creditout_0) );
  OAI22_X1M_A12TR u1660 ( .A0(n1012), .A1(n991), .B0(n1017), .B1(n1018), .Y(
        n1463) );
  INV_X1M_A12TR u1661 ( .A(n137), .Y(n1018) );
  INV_X1M_A12TR u1662 ( .A(n135), .Y(n1017) );
  NOR3_X1M_A12TR u1663 ( .A(n78), .B(n1011), .C(n1270), .Y(n991) );
  INV_X1M_A12TR u1664 ( .A(n124), .Y(n1270) );
  INV_X1M_A12TR u1665 ( .A(n77), .Y(n1011) );
  NOR2_X1M_A12TR u1666 ( .A(n77), .B(n1010), .Y(n1012) );
  OAI21_X1M_A12TR u1667 ( .A0(n1486), .A1(n1483), .B0(n78), .Y(n1010) );
  INV_X1M_A12TR u1668 ( .A(n140), .Y(n1483) );
  INV_X1M_A12TR u1669 ( .A(n6), .Y(n1486) );
  OAI221_X1M_A12TR u1670 ( .A0(n5), .A1(n313), .B0(n1063), .B1(n239), .C0(
        n1062), .Y(flitout_1[0]) );
  OAI221_X1M_A12TR u1671 ( .A0(n5), .A1(n1412), .B0(n1063), .B1(n1243), .C0(
        n1062), .Y(flitout_1[1]) );
  OA21A1OI2_X1M_A12TR u1672 ( .A0(n71), .A1(n5), .B0(n1061), .C0(n1059), .Y(
        n1062) );
  INV_X1M_A12TR u1673 ( .A(n4), .Y(n1059) );
  INV_X1M_A12TR u1674 ( .A(n5), .Y(n1063) );
  OAI22_X1M_A12TR u1675 ( .A0(n314), .A1(n1065), .B0(n240), .B1(n1064), .Y(
        flitout_1[2]) );
  OAI22_X1M_A12TR u1676 ( .A0(n315), .A1(n1065), .B0(n241), .B1(n1064), .Y(
        flitout_1[3]) );
  OAI22_X1M_A12TR u1677 ( .A0(n316), .A1(n1065), .B0(n242), .B1(n1064), .Y(
        flitout_1[4]) );
  OAI22_X1M_A12TR u1678 ( .A0(n317), .A1(n1065), .B0(n243), .B1(n1064), .Y(
        flitout_1[5]) );
  OAI22_X1M_A12TR u1679 ( .A0(n318), .A1(n1065), .B0(n244), .B1(n1064), .Y(
        flitout_1[6]) );
  OAI22_X1M_A12TR u1680 ( .A0(n319), .A1(n1065), .B0(n245), .B1(n1064), .Y(
        flitout_1[7]) );
  OAI22_X1M_A12TR u1681 ( .A0(n24), .A1(n1065), .B0(n104), .B1(n1064), .Y(
        flitout_1[8]) );
  OAI22_X1M_A12TR u1682 ( .A0(n23), .A1(n1065), .B0(n109), .B1(n1064), .Y(
        flitout_1[9]) );
  OAI22_X1M_A12TR u1683 ( .A0(n22), .A1(n1065), .B0(n114), .B1(n1064), .Y(
        flitout_1[10]) );
  OAI22_X1M_A12TR u1684 ( .A0(n21), .A1(n1065), .B0(n119), .B1(n1064), .Y(
        flitout_1[11]) );
  NAND2_X1M_A12TR u1685 ( .A(n4), .B(n1060), .Y(n1065) );
  NOR2_X1M_A12TR u1686 ( .A(n71), .B(n5), .Y(n1060) );
  OAI221_X1M_A12TR u1687 ( .A0(n8), .A1(n313), .B0(n1056), .B1(n239), .C0(
        n1055), .Y(flitout_0[0]) );
  OAI221_X1M_A12TR u1688 ( .A0(n8), .A1(n1412), .B0(n1056), .B1(n1243), .C0(
        n1055), .Y(flitout_0[1]) );
  OA21A1OI2_X1M_A12TR u1689 ( .A0(n8), .A1(n71), .B0(n1054), .C0(n1052), .Y(
        n1055) );
  INV_X1M_A12TR u1690 ( .A(n9), .Y(n1052) );
  INV_X1M_A12TR u1691 ( .A(c0nm_b0m_rdata_1_), .Y(n1243) );
  INV_X1M_A12TR u1692 ( .A(n8), .Y(n1056) );
  INV_X1M_A12TR u1693 ( .A(c0sm_b0m_rdata_1_), .Y(n1412) );
  OAI22_X1M_A12TR u1694 ( .A0(n314), .A1(n1058), .B0(n240), .B1(n1057), .Y(
        flitout_0[2]) );
  OAI22_X1M_A12TR u1695 ( .A0(n315), .A1(n1058), .B0(n241), .B1(n1057), .Y(
        flitout_0[3]) );
  OAI22_X1M_A12TR u1696 ( .A0(n316), .A1(n1058), .B0(n242), .B1(n1057), .Y(
        flitout_0[4]) );
  OAI22_X1M_A12TR u1697 ( .A0(n317), .A1(n1058), .B0(n243), .B1(n1057), .Y(
        flitout_0[5]) );
  OAI22_X1M_A12TR u1698 ( .A0(n318), .A1(n1058), .B0(n244), .B1(n1057), .Y(
        flitout_0[6]) );
  OAI22_X1M_A12TR u1699 ( .A0(n319), .A1(n1058), .B0(n245), .B1(n1057), .Y(
        flitout_0[7]) );
  OAI22_X1M_A12TR u1700 ( .A0(n24), .A1(n1058), .B0(n104), .B1(n1057), .Y(
        flitout_0[8]) );
  OAI22_X1M_A12TR u1701 ( .A0(n23), .A1(n1058), .B0(n109), .B1(n1057), .Y(
        flitout_0[9]) );
  OAI22_X1M_A12TR u1702 ( .A0(n22), .A1(n1058), .B0(n114), .B1(n1057), .Y(
        flitout_0[10]) );
  OAI22_X1M_A12TR u1703 ( .A0(n21), .A1(n1058), .B0(n119), .B1(n1057), .Y(
        flitout_0[11]) );
  NAND2_X1M_A12TR u1704 ( .A(n9), .B(n1053), .Y(n1058) );
  NOR2_X1M_A12TR u1705 ( .A(n71), .B(n8), .Y(n1053) );
  NOR2XB_X1M_A12TR u1706 ( .BN(n1040), .A(n1039), .Y(c0sm_r0m_n11) );
  NOR2XB_X1M_A12TR u1707 ( .BN(n1009), .A(n1008), .Y(c0nm_r0m_n11) );
  AOI2XB1_X1M_A12TR u1708 ( .A1N(n127), .A0(n1205), .B0(n994), .Y(n995) );
  OA22_X1M_A12TR u1709 ( .A0(n1171), .A1(n127), .B0(n1172), .B1(n126), .Y(
        n1097) );
  AOI2XB1_X1M_A12TR u1710 ( .A1N(n17), .A0(n1384), .B0(n1024), .Y(n1025) );
  OA22_X1M_A12TR u1711 ( .A0(n1350), .A1(n17), .B0(n16), .B1(n1351), .Y(n1282)
         );
  NAND2XB_X1M_A12TR u1712 ( .BN(n1232), .A(n1231), .Y(n1233) );
  AO21B_X1M_A12TR u1713 ( .A0(n1011), .A1(n1010), .B0N(n1230), .Y(c0nm_v0m_n57) );
  OA22_X1M_A12TR u1714 ( .A0(n1171), .A1(n131), .B0(n1172), .B1(n130), .Y(
        n1093) );
  OA211_X1M_A12TR u1715 ( .A0(n1076), .A1(n1346), .B0(n1485), .C0(n1070), .Y(
        n968) );
  AND3_X1M_A12TR u1716 ( .A(n1411), .B(n1346), .C(n1051), .Y(n1047) );
  OR2_X1M_A12TR u1717 ( .A(s0m_no_bufs1), .B(n1479), .Y(n1476) );
  OR2_X1M_A12TR u1718 ( .A(s0m_no_bufs0), .B(n1457), .Y(n1454) );
  NAND2XB_X1M_A12TR u1719 ( .BN(n1082), .A(n1081), .Y(n1084) );
  AO21B_X1M_A12TR u1720 ( .A0(n1239), .A1(n7), .B0N(n1438), .Y(n1273) );
  AO21B_X1M_A12TR u1721 ( .A0(n1086), .A1(n73), .B0N(n1440), .Y(n1238) );
  INV_X1M_A12TR u1722 ( .A(n1346), .Y(n1077) );
  INV_X1M_A12TR u1723 ( .A(n148), .Y(n1076) );
  INV_X1M_A12TR u1724 ( .A(n1466), .Y(n1411) );
  NOR2XB_X1M_A12TR u1725 ( .BN(n1041), .A(n12), .Y(n1042) );
  NAND2XB_X1M_A12TR u1726 ( .BN(n1061), .A(n4), .Y(n1064) );
  NAND2XB_X1M_A12TR u1727 ( .BN(n139), .A(n5), .Y(n1061) );
  NAND2XB_X1M_A12TR u1728 ( .BN(n1054), .A(n9), .Y(n1057) );
  NAND2XB_X1M_A12TR u1729 ( .BN(n139), .A(n8), .Y(n1054) );
  NOR3_X0P5A_A12TR u1730 ( .A(n1241), .B(n1099), .C(n168), .Y(
        c0nm_b0m_v0m_n171) );
  NOR3_X0P5A_A12TR u1731 ( .A(n1409), .B(n1284), .C(n158), .Y(
        c0sm_b0m_v0m_n171) );
endmodule

