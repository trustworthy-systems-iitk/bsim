
module oc8051_top ( wb_rst_i, wb_clk_i, wbi_adr_o, wbi_dat_i, wbi_stb_o, 
        wbi_ack_i, wbi_cyc_o, wbi_err_i, wbd_dat_i, wbd_dat_o, wbd_adr_o, 
        wbd_we_o, wbd_ack_i, wbd_stb_o, wbd_cyc_o, wbd_err_i, int0_i, int1_i, 
        p0_i, p0_o, p1_i, p1_o, p2_i, p2_o, p3_i, p3_o, rxd_i, txd_o, t0_i, 
        t1_i, t2_i, t2ex_i, ea_in );
  output [15:0] wbi_adr_o;
  input [31:0] wbi_dat_i;
  input [7:0] wbd_dat_i;
  output [7:0] wbd_dat_o;
  output [15:0] wbd_adr_o;
  input [7:0] p0_i;
  output [7:0] p0_o;
  input [7:0] p1_i;
  output [7:0] p1_o;
  input [7:0] p2_i;
  output [7:0] p2_o;
  input [7:0] p3_i;
  output [7:0] p3_o;
  input wb_rst_i, wb_clk_i, wbi_ack_i, wbi_err_i, wbd_ack_i, wbd_err_i, int0_i,
         int1_i, rxd_i, t0_i, t1_i, t2_i, t2ex_i, ea_in;
  output wbi_stb_o, wbi_cyc_o, wbd_we_o, wbd_stb_o, wbd_cyc_o, txd_o;
  wire   wbd_cyc_o, src_sel3, pc_wr, eq, rd, rmw, istb, mem_wait, wait_data,
         alu_cy, srcac, descy, desac, desov, bit_out, bit_addr_o, n_0_net_,
         bit_data, wr_o, wr_ind, cy, wbi_cyc_o, sfr_bit, intr, int_ack, reti,
         n_3_net_, comp_wait, n_5_net_, n2, n3, oc8051_decoder1_n444,
         oc8051_decoder1_n441, oc8051_decoder1_n440, oc8051_decoder1_n439,
         oc8051_decoder1_n438, oc8051_decoder1_n437, oc8051_decoder1_n436,
         oc8051_decoder1_n435, oc8051_decoder1_n434, oc8051_decoder1_n433,
         oc8051_decoder1_n432, oc8051_decoder1_n431, oc8051_decoder1_n430,
         oc8051_decoder1_n429, oc8051_decoder1_n428, oc8051_decoder1_n427,
         oc8051_decoder1_n426, oc8051_decoder1_n425, oc8051_decoder1_n411,
         oc8051_decoder1_n410, oc8051_decoder1_n409, oc8051_decoder1_n404,
         oc8051_decoder1_n387, oc8051_decoder1_n386, oc8051_decoder1_n385,
         oc8051_decoder1_n384, oc8051_decoder1_n383, oc8051_decoder1_n382,
         oc8051_decoder1_n381, oc8051_decoder1_n380, oc8051_decoder1_n379,
         oc8051_decoder1_n378, oc8051_decoder1_n377, oc8051_decoder1_n376,
         oc8051_decoder1_n375, oc8051_decoder1_n374, oc8051_decoder1_n373,
         oc8051_decoder1_n372, oc8051_decoder1_n371, oc8051_decoder1_n370,
         oc8051_decoder1_n369, oc8051_decoder1_n368, oc8051_decoder1_n367,
         oc8051_decoder1_n366, oc8051_decoder1_n365, oc8051_decoder1_n364,
         oc8051_decoder1_n363, oc8051_decoder1_n362, oc8051_decoder1_n361,
         oc8051_decoder1_n360, oc8051_decoder1_n359, oc8051_decoder1_n358,
         oc8051_decoder1_n357, oc8051_decoder1_n356, oc8051_decoder1_n355,
         oc8051_decoder1_n354, oc8051_decoder1_n353, oc8051_decoder1_n352,
         oc8051_decoder1_n351, oc8051_decoder1_n350, oc8051_decoder1_n349,
         oc8051_decoder1_n348, oc8051_decoder1_n347, oc8051_decoder1_n346,
         oc8051_decoder1_n345, oc8051_decoder1_n344, oc8051_decoder1_n343,
         oc8051_decoder1_n342, oc8051_decoder1_n341, oc8051_decoder1_n340,
         oc8051_decoder1_n339, oc8051_decoder1_n338, oc8051_decoder1_n337,
         oc8051_decoder1_n336, oc8051_decoder1_n335, oc8051_decoder1_n334,
         oc8051_decoder1_n333, oc8051_decoder1_n332, oc8051_decoder1_n331,
         oc8051_decoder1_n330, oc8051_decoder1_n329, oc8051_decoder1_n328,
         oc8051_decoder1_n327, oc8051_decoder1_n326, oc8051_decoder1_n325,
         oc8051_decoder1_n324, oc8051_decoder1_n323, oc8051_decoder1_n322,
         oc8051_decoder1_n321, oc8051_decoder1_n320, oc8051_decoder1_n319,
         oc8051_decoder1_n318, oc8051_decoder1_n317, oc8051_decoder1_n316,
         oc8051_decoder1_n315, oc8051_decoder1_n314, oc8051_decoder1_n313,
         oc8051_decoder1_n312, oc8051_decoder1_n311, oc8051_decoder1_n310,
         oc8051_decoder1_n309, oc8051_decoder1_n308, oc8051_decoder1_n307,
         oc8051_decoder1_n306, oc8051_decoder1_n305, oc8051_decoder1_n304,
         oc8051_decoder1_n303, oc8051_decoder1_n302, oc8051_decoder1_n301,
         oc8051_decoder1_n300, oc8051_decoder1_n299, oc8051_decoder1_n298,
         oc8051_decoder1_n297, oc8051_decoder1_n296, oc8051_decoder1_n295,
         oc8051_decoder1_n294, oc8051_decoder1_n293, oc8051_decoder1_n292,
         oc8051_decoder1_n291, oc8051_decoder1_n290, oc8051_decoder1_n289,
         oc8051_decoder1_n288, oc8051_decoder1_n287, oc8051_decoder1_n286,
         oc8051_decoder1_n285, oc8051_decoder1_n284, oc8051_decoder1_n283,
         oc8051_decoder1_n282, oc8051_decoder1_n281, oc8051_decoder1_n280,
         oc8051_decoder1_n279, oc8051_decoder1_n278, oc8051_decoder1_n277,
         oc8051_decoder1_n276, oc8051_decoder1_n275, oc8051_decoder1_n274,
         oc8051_decoder1_n273, oc8051_decoder1_n272, oc8051_decoder1_n271,
         oc8051_decoder1_n270, oc8051_decoder1_n269, oc8051_decoder1_n268,
         oc8051_decoder1_n267, oc8051_decoder1_n266, oc8051_decoder1_n265,
         oc8051_decoder1_n264, oc8051_decoder1_n263, oc8051_decoder1_n262,
         oc8051_decoder1_n261, oc8051_decoder1_n260, oc8051_decoder1_n259,
         oc8051_decoder1_n258, oc8051_decoder1_n257, oc8051_decoder1_n256,
         oc8051_decoder1_n255, oc8051_decoder1_n254, oc8051_decoder1_n253,
         oc8051_decoder1_n252, oc8051_decoder1_n251, oc8051_decoder1_n250,
         oc8051_decoder1_n249, oc8051_decoder1_n248, oc8051_decoder1_n247,
         oc8051_decoder1_n246, oc8051_decoder1_n245, oc8051_decoder1_n244,
         oc8051_decoder1_n243, oc8051_decoder1_n242, oc8051_decoder1_n241,
         oc8051_decoder1_n240, oc8051_decoder1_n239, oc8051_decoder1_n238,
         oc8051_decoder1_n237, oc8051_decoder1_n236, oc8051_decoder1_n235,
         oc8051_decoder1_n234, oc8051_decoder1_n233, oc8051_decoder1_n232,
         oc8051_decoder1_n231, oc8051_decoder1_n230, oc8051_decoder1_n229,
         oc8051_decoder1_n228, oc8051_decoder1_n227, oc8051_decoder1_n226,
         oc8051_decoder1_n225, oc8051_decoder1_n224, oc8051_decoder1_n223,
         oc8051_decoder1_n222, oc8051_decoder1_n221, oc8051_decoder1_n220,
         oc8051_decoder1_n219, oc8051_decoder1_n218, oc8051_decoder1_n217,
         oc8051_decoder1_n216, oc8051_decoder1_n215, oc8051_decoder1_n214,
         oc8051_decoder1_n213, oc8051_decoder1_n212, oc8051_decoder1_n211,
         oc8051_decoder1_n210, oc8051_decoder1_n209, oc8051_decoder1_n208,
         oc8051_decoder1_n207, oc8051_decoder1_n206, oc8051_decoder1_n205,
         oc8051_decoder1_n204, oc8051_decoder1_n203, oc8051_decoder1_n202,
         oc8051_decoder1_n201, oc8051_decoder1_n200, oc8051_decoder1_n199,
         oc8051_decoder1_n198, oc8051_decoder1_n197, oc8051_decoder1_n196,
         oc8051_decoder1_n195, oc8051_decoder1_n194, oc8051_decoder1_n193,
         oc8051_decoder1_n192, oc8051_decoder1_n191, oc8051_decoder1_n190,
         oc8051_decoder1_n189, oc8051_decoder1_n188, oc8051_decoder1_n187,
         oc8051_decoder1_n186, oc8051_decoder1_n185, oc8051_decoder1_n184,
         oc8051_decoder1_n183, oc8051_decoder1_n182, oc8051_decoder1_n181,
         oc8051_decoder1_n180, oc8051_decoder1_n179, oc8051_decoder1_n178,
         oc8051_decoder1_n177, oc8051_decoder1_n176, oc8051_decoder1_n175,
         oc8051_decoder1_n174, oc8051_decoder1_n173, oc8051_decoder1_n172,
         oc8051_decoder1_n171, oc8051_decoder1_n170, oc8051_decoder1_n169,
         oc8051_decoder1_n168, oc8051_decoder1_n167, oc8051_decoder1_n166,
         oc8051_decoder1_n165, oc8051_decoder1_n164, oc8051_decoder1_n163,
         oc8051_decoder1_n162, oc8051_decoder1_n161, oc8051_decoder1_n160,
         oc8051_decoder1_n159, oc8051_decoder1_n158, oc8051_decoder1_n157,
         oc8051_decoder1_n156, oc8051_decoder1_n155, oc8051_decoder1_n154,
         oc8051_decoder1_n153, oc8051_decoder1_n152, oc8051_decoder1_n151,
         oc8051_decoder1_n150, oc8051_decoder1_n149, oc8051_decoder1_n148,
         oc8051_decoder1_n147, oc8051_decoder1_n146, oc8051_decoder1_n145,
         oc8051_decoder1_n144, oc8051_decoder1_n143, oc8051_decoder1_n142,
         oc8051_decoder1_n141, oc8051_decoder1_n140, oc8051_decoder1_n139,
         oc8051_decoder1_n138, oc8051_decoder1_n137, oc8051_decoder1_n136,
         oc8051_decoder1_n135, oc8051_decoder1_n134, oc8051_decoder1_n133,
         oc8051_decoder1_n132, oc8051_decoder1_n131, oc8051_decoder1_n130,
         oc8051_decoder1_n129, oc8051_decoder1_n128, oc8051_decoder1_n127,
         oc8051_decoder1_n126, oc8051_decoder1_n125, oc8051_decoder1_n124,
         oc8051_decoder1_n123, oc8051_decoder1_n122, oc8051_decoder1_n121,
         oc8051_decoder1_n120, oc8051_decoder1_n119, oc8051_decoder1_n118,
         oc8051_decoder1_n117, oc8051_decoder1_n116, oc8051_decoder1_n115,
         oc8051_decoder1_n114, oc8051_decoder1_n113, oc8051_decoder1_n112,
         oc8051_decoder1_n111, oc8051_decoder1_n110, oc8051_decoder1_n109,
         oc8051_decoder1_n108, oc8051_decoder1_n107, oc8051_decoder1_n106,
         oc8051_decoder1_n105, oc8051_decoder1_n104, oc8051_decoder1_n103,
         oc8051_decoder1_n102, oc8051_decoder1_n101, oc8051_decoder1_n100,
         oc8051_decoder1_n99, oc8051_decoder1_n98, oc8051_decoder1_n97,
         oc8051_decoder1_n96, oc8051_decoder1_n95, oc8051_decoder1_n94,
         oc8051_decoder1_n93, oc8051_decoder1_n92, oc8051_decoder1_n91,
         oc8051_decoder1_n90, oc8051_decoder1_n89, oc8051_decoder1_n88,
         oc8051_decoder1_n87, oc8051_decoder1_n86, oc8051_decoder1_n85,
         oc8051_decoder1_n84, oc8051_decoder1_n83, oc8051_decoder1_n82,
         oc8051_decoder1_n81, oc8051_decoder1_n80, oc8051_decoder1_n79,
         oc8051_decoder1_n78, oc8051_decoder1_n77, oc8051_decoder1_n76,
         oc8051_decoder1_n75, oc8051_decoder1_n74, oc8051_decoder1_n73,
         oc8051_decoder1_n72, oc8051_decoder1_n71, oc8051_decoder1_n70,
         oc8051_decoder1_n69, oc8051_decoder1_n68, oc8051_decoder1_n67,
         oc8051_decoder1_n66, oc8051_decoder1_n65, oc8051_decoder1_n64,
         oc8051_decoder1_n63, oc8051_decoder1_n62, oc8051_decoder1_n61,
         oc8051_decoder1_n60, oc8051_decoder1_n59, oc8051_decoder1_n58,
         oc8051_decoder1_n57, oc8051_decoder1_n56, oc8051_decoder1_n55,
         oc8051_decoder1_n54, oc8051_decoder1_n53, oc8051_decoder1_n52,
         oc8051_decoder1_n51, oc8051_decoder1_n50, oc8051_decoder1_n49,
         oc8051_decoder1_n48, oc8051_decoder1_n47, oc8051_decoder1_n46,
         oc8051_decoder1_n45, oc8051_decoder1_n44, oc8051_decoder1_n43,
         oc8051_decoder1_n42, oc8051_decoder1_n41, oc8051_decoder1_n40,
         oc8051_decoder1_n39, oc8051_decoder1_n38, oc8051_decoder1_n37,
         oc8051_decoder1_n36, oc8051_decoder1_n35, oc8051_decoder1_n34,
         oc8051_decoder1_n33, oc8051_decoder1_n32, oc8051_decoder1_n31,
         oc8051_decoder1_n30, oc8051_decoder1_n29, oc8051_decoder1_n28,
         oc8051_decoder1_n27, oc8051_decoder1_n26, oc8051_decoder1_n25,
         oc8051_decoder1_n24, oc8051_decoder1_n23, oc8051_decoder1_n22,
         oc8051_decoder1_n21, oc8051_decoder1_n20, oc8051_decoder1_n19,
         oc8051_decoder1_n18, oc8051_decoder1_n17, oc8051_decoder1_n16,
         oc8051_decoder1_n15, oc8051_decoder1_n14, oc8051_decoder1_n13,
         oc8051_decoder1_n12, oc8051_decoder1_n11, oc8051_decoder1_n10,
         oc8051_decoder1_n9, oc8051_decoder1_n8, oc8051_decoder1_n7,
         oc8051_decoder1_n6, oc8051_decoder1_n5, oc8051_decoder1_n4,
         oc8051_decoder1_n3, oc8051_decoder1_n2, oc8051_decoder1_n1,
         oc8051_decoder1_n424, oc8051_decoder1_n423, oc8051_decoder1_n422,
         oc8051_decoder1_n421, oc8051_decoder1_n420, oc8051_decoder1_n419,
         oc8051_decoder1_n418, oc8051_decoder1_n417, oc8051_decoder1_n416,
         oc8051_decoder1_n415, oc8051_decoder1_n414, oc8051_decoder1_n413,
         oc8051_decoder1_n412, oc8051_decoder1_n408, oc8051_decoder1_n407,
         oc8051_decoder1_n406, oc8051_decoder1_n405, oc8051_decoder1_n403,
         oc8051_decoder1_n402, oc8051_decoder1_n401, oc8051_decoder1_n400,
         oc8051_decoder1_n399, oc8051_decoder1_n398, oc8051_decoder1_n397,
         oc8051_decoder1_n396, oc8051_decoder1_n395, oc8051_decoder1_n394,
         oc8051_decoder1_n393, oc8051_decoder1_n392, oc8051_decoder1_n391,
         oc8051_decoder1_n390, oc8051_decoder1_n389, oc8051_decoder1_n388,
         oc8051_decoder1_n1806, oc8051_decoder1_n1805, oc8051_decoder1_n1804,
         oc8051_decoder1_wr, oc8051_decoder1_ram_wr_sel_0_,
         oc8051_decoder1_ram_wr_sel_1_, oc8051_decoder1_ram_rd_sel_0_,
         oc8051_decoder1_ram_rd_sel_1_, oc8051_decoder1_alu_op_0_,
         oc8051_decoder1_alu_op_1_, oc8051_decoder1_alu_op_2_,
         oc8051_decoder1_alu_op_3_, oc8051_decoder1_state_0_,
         oc8051_decoder1_state_1_, oc8051_alu1_n290, oc8051_alu1_n289,
         oc8051_alu1_n288, oc8051_alu1_n283, oc8051_alu1_n282,
         oc8051_alu1_n281, oc8051_alu1_n280, oc8051_alu1_n279,
         oc8051_alu1_n278, oc8051_alu1_n277, oc8051_alu1_n276,
         oc8051_alu1_n275, oc8051_alu1_n274, oc8051_alu1_n273,
         oc8051_alu1_n272, oc8051_alu1_n271, oc8051_alu1_n270,
         oc8051_alu1_n269, oc8051_alu1_n268, oc8051_alu1_n267,
         oc8051_alu1_n266, oc8051_alu1_n265, oc8051_alu1_n264,
         oc8051_alu1_n263, oc8051_alu1_n262, oc8051_alu1_n261,
         oc8051_alu1_n260, oc8051_alu1_n259, oc8051_alu1_n258,
         oc8051_alu1_n257, oc8051_alu1_n256, oc8051_alu1_n255,
         oc8051_alu1_n254, oc8051_alu1_n253, oc8051_alu1_n252,
         oc8051_alu1_n251, oc8051_alu1_n250, oc8051_alu1_n249,
         oc8051_alu1_n248, oc8051_alu1_n247, oc8051_alu1_n246,
         oc8051_alu1_n245, oc8051_alu1_n244, oc8051_alu1_n243,
         oc8051_alu1_n242, oc8051_alu1_n241, oc8051_alu1_n240,
         oc8051_alu1_n239, oc8051_alu1_n238, oc8051_alu1_n237,
         oc8051_alu1_n236, oc8051_alu1_n235, oc8051_alu1_n234,
         oc8051_alu1_n233, oc8051_alu1_n232, oc8051_alu1_n231,
         oc8051_alu1_n230, oc8051_alu1_n229, oc8051_alu1_n228,
         oc8051_alu1_n227, oc8051_alu1_n226, oc8051_alu1_n225,
         oc8051_alu1_n224, oc8051_alu1_n223, oc8051_alu1_n222,
         oc8051_alu1_n221, oc8051_alu1_n220, oc8051_alu1_n219,
         oc8051_alu1_n218, oc8051_alu1_n217, oc8051_alu1_n216,
         oc8051_alu1_n215, oc8051_alu1_n214, oc8051_alu1_n213,
         oc8051_alu1_n212, oc8051_alu1_n211, oc8051_alu1_n210,
         oc8051_alu1_n209, oc8051_alu1_n208, oc8051_alu1_n207,
         oc8051_alu1_n206, oc8051_alu1_n205, oc8051_alu1_n204,
         oc8051_alu1_n203, oc8051_alu1_n202, oc8051_alu1_n201,
         oc8051_alu1_n200, oc8051_alu1_n199, oc8051_alu1_n198,
         oc8051_alu1_n197, oc8051_alu1_n196, oc8051_alu1_n195,
         oc8051_alu1_n194, oc8051_alu1_n193, oc8051_alu1_n192,
         oc8051_alu1_n191, oc8051_alu1_n190, oc8051_alu1_n189,
         oc8051_alu1_n188, oc8051_alu1_n187, oc8051_alu1_n186,
         oc8051_alu1_n185, oc8051_alu1_n184, oc8051_alu1_n183,
         oc8051_alu1_n182, oc8051_alu1_n181, oc8051_alu1_n180,
         oc8051_alu1_n179, oc8051_alu1_n178, oc8051_alu1_n177,
         oc8051_alu1_n176, oc8051_alu1_n175, oc8051_alu1_n174,
         oc8051_alu1_n173, oc8051_alu1_n172, oc8051_alu1_n171,
         oc8051_alu1_n170, oc8051_alu1_n169, oc8051_alu1_n168,
         oc8051_alu1_n167, oc8051_alu1_n166, oc8051_alu1_n165,
         oc8051_alu1_n164, oc8051_alu1_n163, oc8051_alu1_n162,
         oc8051_alu1_n161, oc8051_alu1_n160, oc8051_alu1_n159,
         oc8051_alu1_n158, oc8051_alu1_n157, oc8051_alu1_n156,
         oc8051_alu1_n155, oc8051_alu1_n154, oc8051_alu1_n153,
         oc8051_alu1_n152, oc8051_alu1_n151, oc8051_alu1_n150,
         oc8051_alu1_n149, oc8051_alu1_n148, oc8051_alu1_n147,
         oc8051_alu1_n146, oc8051_alu1_n145, oc8051_alu1_n144,
         oc8051_alu1_n143, oc8051_alu1_n142, oc8051_alu1_n141,
         oc8051_alu1_n140, oc8051_alu1_n139, oc8051_alu1_n138,
         oc8051_alu1_n137, oc8051_alu1_n136, oc8051_alu1_n135,
         oc8051_alu1_n134, oc8051_alu1_n133, oc8051_alu1_n132,
         oc8051_alu1_n131, oc8051_alu1_n130, oc8051_alu1_n129,
         oc8051_alu1_n128, oc8051_alu1_n127, oc8051_alu1_n126,
         oc8051_alu1_n125, oc8051_alu1_n124, oc8051_alu1_n123,
         oc8051_alu1_n122, oc8051_alu1_n121, oc8051_alu1_n120,
         oc8051_alu1_n119, oc8051_alu1_n118, oc8051_alu1_n117,
         oc8051_alu1_n116, oc8051_alu1_n115, oc8051_alu1_n114,
         oc8051_alu1_n113, oc8051_alu1_n112, oc8051_alu1_n111,
         oc8051_alu1_n110, oc8051_alu1_n109, oc8051_alu1_n108,
         oc8051_alu1_n107, oc8051_alu1_n106, oc8051_alu1_n105,
         oc8051_alu1_n104, oc8051_alu1_n103, oc8051_alu1_n102,
         oc8051_alu1_n101, oc8051_alu1_n100, oc8051_alu1_n99, oc8051_alu1_n98,
         oc8051_alu1_n97, oc8051_alu1_n96, oc8051_alu1_n95, oc8051_alu1_n94,
         oc8051_alu1_n93, oc8051_alu1_n92, oc8051_alu1_n91, oc8051_alu1_n90,
         oc8051_alu1_n89, oc8051_alu1_n88, oc8051_alu1_n87, oc8051_alu1_n86,
         oc8051_alu1_n85, oc8051_alu1_n84, oc8051_alu1_n83, oc8051_alu1_n82,
         oc8051_alu1_n81, oc8051_alu1_n80, oc8051_alu1_n79, oc8051_alu1_n78,
         oc8051_alu1_n77, oc8051_alu1_n76, oc8051_alu1_n75, oc8051_alu1_n74,
         oc8051_alu1_n73, oc8051_alu1_n72, oc8051_alu1_n71, oc8051_alu1_n70,
         oc8051_alu1_n69, oc8051_alu1_n68, oc8051_alu1_n67, oc8051_alu1_n66,
         oc8051_alu1_n65, oc8051_alu1_n64, oc8051_alu1_n63, oc8051_alu1_n62,
         oc8051_alu1_n61, oc8051_alu1_n60, oc8051_alu1_n59, oc8051_alu1_n58,
         oc8051_alu1_n57, oc8051_alu1_n56, oc8051_alu1_n55, oc8051_alu1_n54,
         oc8051_alu1_n53, oc8051_alu1_n52, oc8051_alu1_n51, oc8051_alu1_n50,
         oc8051_alu1_n49, oc8051_alu1_n48, oc8051_alu1_n47, oc8051_alu1_n46,
         oc8051_alu1_n45, oc8051_alu1_n44, oc8051_alu1_n43, oc8051_alu1_n42,
         oc8051_alu1_n41, oc8051_alu1_n40, oc8051_alu1_n39, oc8051_alu1_n38,
         oc8051_alu1_n37, oc8051_alu1_n36, oc8051_alu1_n35, oc8051_alu1_n34,
         oc8051_alu1_n33, oc8051_alu1_n32, oc8051_alu1_n31, oc8051_alu1_n30,
         oc8051_alu1_n29, oc8051_alu1_n28, oc8051_alu1_n27, oc8051_alu1_n26,
         oc8051_alu1_n25, oc8051_alu1_n24, oc8051_alu1_n23, oc8051_alu1_n22,
         oc8051_alu1_n21, oc8051_alu1_n20, oc8051_alu1_n19, oc8051_alu1_n18,
         oc8051_alu1_n17, oc8051_alu1_n16, oc8051_alu1_n15, oc8051_alu1_n13,
         oc8051_alu1_n12, oc8051_alu1_n11, oc8051_alu1_n10, oc8051_alu1_n9,
         oc8051_alu1_n8, oc8051_alu1_n7, oc8051_alu1_n6, oc8051_alu1_n5,
         oc8051_alu1_n4, oc8051_alu1_n3, oc8051_alu1_n2, oc8051_alu1_n1,
         oc8051_alu1_n14, oc8051_alu1_n2400, oc8051_alu1_n2200,
         oc8051_alu1_n2190, oc8051_alu1_n2180, oc8051_alu1_n2170,
         oc8051_alu1_n2160, oc8051_alu1_n2150, oc8051_alu1_n2140,
         oc8051_alu1_n2130, oc8051_alu1_divov, oc8051_alu1_mulov,
         oc8051_alu1_malicious1, oc8051_alu1_alu_malicious_n7,
         oc8051_alu1_alu_malicious_n6, oc8051_alu1_alu_malicious_n5,
         oc8051_alu1_alu_malicious_n4, oc8051_alu1_alu_malicious_n3,
         oc8051_alu1_alu_malicious_n2, oc8051_alu1_alu_malicious_n1,
         oc8051_alu1_alu_malicious_n9, oc8051_alu1_alu_malicious_n8,
         oc8051_alu1_alu_malicious_n70, oc8051_alu1_alu_malicious_state_0_,
         oc8051_alu1_alu_malicious_state_1_, oc8051_alu1_oc8051_mul1_n55,
         oc8051_alu1_oc8051_mul1_n54, oc8051_alu1_oc8051_mul1_n53,
         oc8051_alu1_oc8051_mul1_n52, oc8051_alu1_oc8051_mul1_n51,
         oc8051_alu1_oc8051_mul1_n50, oc8051_alu1_oc8051_mul1_n49,
         oc8051_alu1_oc8051_mul1_n48, oc8051_alu1_oc8051_mul1_n47,
         oc8051_alu1_oc8051_mul1_n46, oc8051_alu1_oc8051_mul1_n45,
         oc8051_alu1_oc8051_mul1_n44, oc8051_alu1_oc8051_mul1_n43,
         oc8051_alu1_oc8051_mul1_n42, oc8051_alu1_oc8051_mul1_n41,
         oc8051_alu1_oc8051_mul1_n40, oc8051_alu1_oc8051_mul1_n39,
         oc8051_alu1_oc8051_mul1_n38, oc8051_alu1_oc8051_mul1_n37,
         oc8051_alu1_oc8051_mul1_n36, oc8051_alu1_oc8051_mul1_n35,
         oc8051_alu1_oc8051_mul1_n34, oc8051_alu1_oc8051_mul1_n33,
         oc8051_alu1_oc8051_mul1_n32, oc8051_alu1_oc8051_mul1_n31,
         oc8051_alu1_oc8051_mul1_n30, oc8051_alu1_oc8051_mul1_n29,
         oc8051_alu1_oc8051_mul1_n28, oc8051_alu1_oc8051_mul1_n27,
         oc8051_alu1_oc8051_mul1_n26, oc8051_alu1_oc8051_mul1_n25,
         oc8051_alu1_oc8051_mul1_n24, oc8051_alu1_oc8051_mul1_n23,
         oc8051_alu1_oc8051_mul1_n22, oc8051_alu1_oc8051_mul1_n21,
         oc8051_alu1_oc8051_mul1_n20, oc8051_alu1_oc8051_mul1_n19,
         oc8051_alu1_oc8051_mul1_n18, oc8051_alu1_oc8051_mul1_n16,
         oc8051_alu1_oc8051_mul1_n15, oc8051_alu1_oc8051_mul1_n14,
         oc8051_alu1_oc8051_mul1_n13, oc8051_alu1_oc8051_mul1_n12,
         oc8051_alu1_oc8051_mul1_n11, oc8051_alu1_oc8051_mul1_n10,
         oc8051_alu1_oc8051_mul1_n9, oc8051_alu1_oc8051_mul1_n8,
         oc8051_alu1_oc8051_mul1_n7, oc8051_alu1_oc8051_mul1_n6,
         oc8051_alu1_oc8051_mul1_n5, oc8051_alu1_oc8051_mul1_n4,
         oc8051_alu1_oc8051_mul1_n3, oc8051_alu1_oc8051_mul1_n2,
         oc8051_alu1_oc8051_mul1_n1, oc8051_alu1_oc8051_mul1_n17,
         oc8051_alu1_oc8051_mul1_tmp_mul_0_,
         oc8051_alu1_oc8051_mul1_tmp_mul_1_,
         oc8051_alu1_oc8051_mul1_tmp_mul_2_,
         oc8051_alu1_oc8051_mul1_tmp_mul_3_,
         oc8051_alu1_oc8051_mul1_tmp_mul_4_,
         oc8051_alu1_oc8051_mul1_tmp_mul_5_,
         oc8051_alu1_oc8051_mul1_tmp_mul_6_,
         oc8051_alu1_oc8051_mul1_tmp_mul_7_,
         oc8051_alu1_oc8051_mul1_tmp_mul_8_,
         oc8051_alu1_oc8051_mul1_tmp_mul_9_,
         oc8051_alu1_oc8051_mul1_tmp_mul_10_,
         oc8051_alu1_oc8051_mul1_tmp_mul_11_,
         oc8051_alu1_oc8051_mul1_tmp_mul_12_,
         oc8051_alu1_oc8051_mul1_tmp_mul_13_,
         oc8051_alu1_oc8051_mul1_mul_result1_2_,
         oc8051_alu1_oc8051_mul1_mul_result1_3_,
         oc8051_alu1_oc8051_mul1_mul_result1_4_,
         oc8051_alu1_oc8051_mul1_mul_result1_5_,
         oc8051_alu1_oc8051_mul1_mul_result1_6_,
         oc8051_alu1_oc8051_mul1_mul_result1_7_,
         oc8051_alu1_oc8051_mul1_mul_result1_8_,
         oc8051_alu1_oc8051_mul1_mul_result1_9_, oc8051_alu1_oc8051_mul1_n80,
         oc8051_alu1_oc8051_mul1_n70, oc8051_alu1_oc8051_mul1_cycle_0_,
         oc8051_alu1_oc8051_mul1_cycle_1_, oc8051_alu1_oc8051_mul1_mult_90_n33,
         oc8051_alu1_oc8051_mul1_mult_90_n32,
         oc8051_alu1_oc8051_mul1_mult_90_n31,
         oc8051_alu1_oc8051_mul1_mult_90_n30,
         oc8051_alu1_oc8051_mul1_mult_90_n29,
         oc8051_alu1_oc8051_mul1_mult_90_n28,
         oc8051_alu1_oc8051_mul1_mult_90_n27,
         oc8051_alu1_oc8051_mul1_mult_90_n26,
         oc8051_alu1_oc8051_mul1_mult_90_n25,
         oc8051_alu1_oc8051_mul1_mult_90_n24,
         oc8051_alu1_oc8051_mul1_mult_90_n23,
         oc8051_alu1_oc8051_mul1_mult_90_n22,
         oc8051_alu1_oc8051_mul1_mult_90_n21,
         oc8051_alu1_oc8051_mul1_mult_90_n20,
         oc8051_alu1_oc8051_mul1_mult_90_n19,
         oc8051_alu1_oc8051_mul1_mult_90_n18,
         oc8051_alu1_oc8051_mul1_mult_90_n17,
         oc8051_alu1_oc8051_mul1_mult_90_n16,
         oc8051_alu1_oc8051_mul1_mult_90_n15,
         oc8051_alu1_oc8051_mul1_mult_90_n14,
         oc8051_alu1_oc8051_mul1_mult_90_n13,
         oc8051_alu1_oc8051_mul1_mult_90_n12,
         oc8051_alu1_oc8051_mul1_mult_90_n11,
         oc8051_alu1_oc8051_mul1_mult_90_n10,
         oc8051_alu1_oc8051_mul1_mult_90_n9,
         oc8051_alu1_oc8051_mul1_mult_90_n8,
         oc8051_alu1_oc8051_mul1_mult_90_n7,
         oc8051_alu1_oc8051_mul1_mult_90_n6,
         oc8051_alu1_oc8051_mul1_mult_90_n5,
         oc8051_alu1_oc8051_mul1_mult_90_n4,
         oc8051_alu1_oc8051_mul1_mult_90_n3,
         oc8051_alu1_oc8051_mul1_mult_90_n2, oc8051_alu1_oc8051_div1_n30,
         oc8051_alu1_oc8051_div1_n29, oc8051_alu1_oc8051_div1_n28,
         oc8051_alu1_oc8051_div1_n27, oc8051_alu1_oc8051_div1_n24,
         oc8051_alu1_oc8051_div1_n23, oc8051_alu1_oc8051_div1_n22,
         oc8051_alu1_oc8051_div1_n21, oc8051_alu1_oc8051_div1_n20,
         oc8051_alu1_oc8051_div1_n19, oc8051_alu1_oc8051_div1_n18,
         oc8051_alu1_oc8051_div1_n17, oc8051_alu1_oc8051_div1_n16,
         oc8051_alu1_oc8051_div1_n15, oc8051_alu1_oc8051_div1_n14,
         oc8051_alu1_oc8051_div1_n13, oc8051_alu1_oc8051_div1_n12,
         oc8051_alu1_oc8051_div1_n11, oc8051_alu1_oc8051_div1_n10,
         oc8051_alu1_oc8051_div1_n9, oc8051_alu1_oc8051_div1_n8,
         oc8051_alu1_oc8051_div1_n7, oc8051_alu1_oc8051_div1_n6,
         oc8051_alu1_oc8051_div1_n5, oc8051_alu1_oc8051_div1_n4,
         oc8051_alu1_oc8051_div1_n3, oc8051_alu1_oc8051_div1_n2,
         oc8051_alu1_oc8051_div1_n26, oc8051_alu1_oc8051_div1_n25,
         oc8051_alu1_oc8051_div1_cmp1_0_, oc8051_alu1_oc8051_div1_rem1_0_,
         oc8051_alu1_oc8051_div1_rem1_1_, oc8051_alu1_oc8051_div1_rem1_2_,
         oc8051_alu1_oc8051_div1_rem1_3_, oc8051_alu1_oc8051_div1_rem1_4_,
         oc8051_alu1_oc8051_div1_rem1_5_, oc8051_alu1_oc8051_div1_rem1_6_,
         oc8051_alu1_oc8051_div1_rem1_7_, oc8051_alu1_oc8051_div1_rem2_1_,
         oc8051_alu1_oc8051_div1_rem2_2_, oc8051_alu1_oc8051_div1_rem2_3_,
         oc8051_alu1_oc8051_div1_rem2_4_, oc8051_alu1_oc8051_div1_rem2_5_,
         oc8051_alu1_oc8051_div1_rem2_6_, oc8051_alu1_oc8051_div1_rem2_7_,
         oc8051_alu1_oc8051_div1_cmp0_7_, oc8051_alu1_oc8051_div1_cmp1_1_,
         oc8051_alu1_oc8051_div1_cmp1_2_, oc8051_alu1_oc8051_div1_cmp1_3_,
         oc8051_alu1_oc8051_div1_cmp1_4_, oc8051_alu1_oc8051_div1_cmp1_5_,
         oc8051_alu1_oc8051_div1_cmp1_6_, oc8051_alu1_oc8051_div1_cmp1_7_,
         oc8051_alu1_oc8051_div1_cycle_0_, oc8051_alu1_oc8051_div1_cycle_1_,
         oc8051_alu1_oc8051_div1_sub_98_n10, oc8051_alu1_oc8051_div1_sub_98_n9,
         oc8051_alu1_oc8051_div1_sub_98_n8, oc8051_alu1_oc8051_div1_sub_98_n7,
         oc8051_alu1_oc8051_div1_sub_98_n6, oc8051_alu1_oc8051_div1_sub_98_n5,
         oc8051_alu1_oc8051_div1_sub_98_n4, oc8051_alu1_oc8051_div1_sub_98_n3,
         oc8051_alu1_oc8051_div1_sub_98_n1, oc8051_alu1_oc8051_div1_sub_94_n9,
         oc8051_alu1_oc8051_div1_sub_94_n8, oc8051_alu1_oc8051_div1_sub_94_n7,
         oc8051_alu1_oc8051_div1_sub_94_n6, oc8051_alu1_oc8051_div1_sub_94_n5,
         oc8051_alu1_oc8051_div1_sub_94_n4, oc8051_alu1_oc8051_div1_sub_94_n3,
         oc8051_alu1_oc8051_div1_sub_94_n1, oc8051_alu1_sub_205_n14,
         oc8051_alu1_sub_205_n13, oc8051_alu1_sub_205_n12,
         oc8051_alu1_sub_205_n11, oc8051_alu1_sub_205_n10,
         oc8051_alu1_sub_205_n9, oc8051_alu1_sub_205_n8,
         oc8051_alu1_sub_205_n7, oc8051_alu1_sub_205_n6,
         oc8051_alu1_sub_205_n5, oc8051_alu1_sub_205_n4,
         oc8051_alu1_sub_205_n3, oc8051_alu1_sub_205_n2,
         oc8051_alu1_sub_205_n1, oc8051_ram_top1_n76, oc8051_ram_top1_n75,
         oc8051_ram_top1_n74, oc8051_ram_top1_n73, oc8051_ram_top1_n72,
         oc8051_ram_top1_n71, oc8051_ram_top1_n70, oc8051_ram_top1_n69,
         oc8051_ram_top1_n68, oc8051_ram_top1_n67, oc8051_ram_top1_n66,
         oc8051_ram_top1_n65, oc8051_ram_top1_n64, oc8051_ram_top1_n63,
         oc8051_ram_top1_n62, oc8051_ram_top1_n61, oc8051_ram_top1_n60,
         oc8051_ram_top1_n59, oc8051_ram_top1_n58, oc8051_ram_top1_n57,
         oc8051_ram_top1_n56, oc8051_ram_top1_n55, oc8051_ram_top1_n54,
         oc8051_ram_top1_n52, oc8051_ram_top1_n51, oc8051_ram_top1_n50,
         oc8051_ram_top1_n49, oc8051_ram_top1_n48, oc8051_ram_top1_n47,
         oc8051_ram_top1_n46, oc8051_ram_top1_n45, oc8051_ram_top1_n44,
         oc8051_ram_top1_n43, oc8051_ram_top1_n42, oc8051_ram_top1_n41,
         oc8051_ram_top1_n40, oc8051_ram_top1_n39, oc8051_ram_top1_n38,
         oc8051_ram_top1_n37, oc8051_ram_top1_n36, oc8051_ram_top1_n35,
         oc8051_ram_top1_n34, oc8051_ram_top1_n33, oc8051_ram_top1_n32,
         oc8051_ram_top1_n31, oc8051_ram_top1_n30, oc8051_ram_top1_n29,
         oc8051_ram_top1_n28, oc8051_ram_top1_n27, oc8051_ram_top1_n26,
         oc8051_ram_top1_n25, oc8051_ram_top1_n24, oc8051_ram_top1_n23,
         oc8051_ram_top1_n22, oc8051_ram_top1_n21, oc8051_ram_top1_n20,
         oc8051_ram_top1_n19, oc8051_ram_top1_n18, oc8051_ram_top1_n17,
         oc8051_ram_top1_n16, oc8051_ram_top1_n15, oc8051_ram_top1_n14,
         oc8051_ram_top1_n13, oc8051_ram_top1_n12, oc8051_ram_top1_n11,
         oc8051_ram_top1_n10, oc8051_ram_top1_n9, oc8051_ram_top1_n8,
         oc8051_ram_top1_n7, oc8051_ram_top1_n6, oc8051_ram_top1_n5,
         oc8051_ram_top1_n4, oc8051_ram_top1_n3, oc8051_ram_top1_n2,
         oc8051_ram_top1_n1, oc8051_ram_top1_n53, oc8051_ram_top1_bit_addr_r,
         oc8051_ram_top1_wr_addr_m_0_, oc8051_ram_top1_wr_addr_m_1_,
         oc8051_ram_top1_wr_addr_m_2_, oc8051_ram_top1_wr_addr_m_3_,
         oc8051_ram_top1_wr_addr_m_4_, oc8051_ram_top1_wr_addr_m_5_,
         oc8051_ram_top1_wr_addr_m_6_, oc8051_ram_top1_rd_addr_m_0_,
         oc8051_ram_top1_rd_addr_m_1_, oc8051_ram_top1_rd_addr_m_2_,
         oc8051_ram_top1_rd_addr_m_3_, oc8051_ram_top1_rd_addr_m_4_,
         oc8051_ram_top1_rd_addr_m_5_, oc8051_ram_top1_rd_addr_m_6_,
         oc8051_ram_top1_rd_en_r, oc8051_ram_top1__logic1_,
         oc8051_ram_top1_n280, oc8051_ram_top1_n270, oc8051_ram_top1_n260,
         oc8051_ram_top1_oc8051_idata_n4654,
         oc8051_ram_top1_oc8051_idata_n4653,
         oc8051_ram_top1_oc8051_idata_n4652,
         oc8051_ram_top1_oc8051_idata_n4651,
         oc8051_ram_top1_oc8051_idata_n4650,
         oc8051_ram_top1_oc8051_idata_n4649,
         oc8051_ram_top1_oc8051_idata_n4648,
         oc8051_ram_top1_oc8051_idata_n4647,
         oc8051_ram_top1_oc8051_idata_n4646,
         oc8051_ram_top1_oc8051_idata_n4645,
         oc8051_ram_top1_oc8051_idata_n4644,
         oc8051_ram_top1_oc8051_idata_n4643,
         oc8051_ram_top1_oc8051_idata_n4642,
         oc8051_ram_top1_oc8051_idata_n4641,
         oc8051_ram_top1_oc8051_idata_n4640,
         oc8051_ram_top1_oc8051_idata_n4639,
         oc8051_ram_top1_oc8051_idata_n4638,
         oc8051_ram_top1_oc8051_idata_n4637,
         oc8051_ram_top1_oc8051_idata_n4636,
         oc8051_ram_top1_oc8051_idata_n4635,
         oc8051_ram_top1_oc8051_idata_n4634,
         oc8051_ram_top1_oc8051_idata_n4633,
         oc8051_ram_top1_oc8051_idata_n4632,
         oc8051_ram_top1_oc8051_idata_n4631,
         oc8051_ram_top1_oc8051_idata_n4630,
         oc8051_ram_top1_oc8051_idata_n4629,
         oc8051_ram_top1_oc8051_idata_n4628,
         oc8051_ram_top1_oc8051_idata_n4627,
         oc8051_ram_top1_oc8051_idata_n4626,
         oc8051_ram_top1_oc8051_idata_n4625,
         oc8051_ram_top1_oc8051_idata_n4624,
         oc8051_ram_top1_oc8051_idata_n4623,
         oc8051_ram_top1_oc8051_idata_n4622,
         oc8051_ram_top1_oc8051_idata_n4621,
         oc8051_ram_top1_oc8051_idata_n4620,
         oc8051_ram_top1_oc8051_idata_n4619,
         oc8051_ram_top1_oc8051_idata_n4618,
         oc8051_ram_top1_oc8051_idata_n4617,
         oc8051_ram_top1_oc8051_idata_n4616,
         oc8051_ram_top1_oc8051_idata_n4615,
         oc8051_ram_top1_oc8051_idata_n4614,
         oc8051_ram_top1_oc8051_idata_n4613,
         oc8051_ram_top1_oc8051_idata_n4612,
         oc8051_ram_top1_oc8051_idata_n4611,
         oc8051_ram_top1_oc8051_idata_n4610,
         oc8051_ram_top1_oc8051_idata_n4609,
         oc8051_ram_top1_oc8051_idata_n4608,
         oc8051_ram_top1_oc8051_idata_n4607,
         oc8051_ram_top1_oc8051_idata_n4606,
         oc8051_ram_top1_oc8051_idata_n4605,
         oc8051_ram_top1_oc8051_idata_n4604,
         oc8051_ram_top1_oc8051_idata_n4603,
         oc8051_ram_top1_oc8051_idata_n4602,
         oc8051_ram_top1_oc8051_idata_n4601,
         oc8051_ram_top1_oc8051_idata_n4600,
         oc8051_ram_top1_oc8051_idata_n4599,
         oc8051_ram_top1_oc8051_idata_n4598,
         oc8051_ram_top1_oc8051_idata_n4597,
         oc8051_ram_top1_oc8051_idata_n4596,
         oc8051_ram_top1_oc8051_idata_n4595,
         oc8051_ram_top1_oc8051_idata_n4594,
         oc8051_ram_top1_oc8051_idata_n4593,
         oc8051_ram_top1_oc8051_idata_n4592,
         oc8051_ram_top1_oc8051_idata_n4591,
         oc8051_ram_top1_oc8051_idata_n4590,
         oc8051_ram_top1_oc8051_idata_n4589,
         oc8051_ram_top1_oc8051_idata_n4588,
         oc8051_ram_top1_oc8051_idata_n4587,
         oc8051_ram_top1_oc8051_idata_n4586,
         oc8051_ram_top1_oc8051_idata_n4585,
         oc8051_ram_top1_oc8051_idata_n4584,
         oc8051_ram_top1_oc8051_idata_n4583,
         oc8051_ram_top1_oc8051_idata_n4582,
         oc8051_ram_top1_oc8051_idata_n4581,
         oc8051_ram_top1_oc8051_idata_n4580,
         oc8051_ram_top1_oc8051_idata_n4579,
         oc8051_ram_top1_oc8051_idata_n4578,
         oc8051_ram_top1_oc8051_idata_n4577,
         oc8051_ram_top1_oc8051_idata_n4576,
         oc8051_ram_top1_oc8051_idata_n4575,
         oc8051_ram_top1_oc8051_idata_n4574,
         oc8051_ram_top1_oc8051_idata_n4573,
         oc8051_ram_top1_oc8051_idata_n4572,
         oc8051_ram_top1_oc8051_idata_n4571,
         oc8051_ram_top1_oc8051_idata_n4570,
         oc8051_ram_top1_oc8051_idata_n4569,
         oc8051_ram_top1_oc8051_idata_n4568,
         oc8051_ram_top1_oc8051_idata_n4567,
         oc8051_ram_top1_oc8051_idata_n4566,
         oc8051_ram_top1_oc8051_idata_n4565,
         oc8051_ram_top1_oc8051_idata_n4564,
         oc8051_ram_top1_oc8051_idata_n4563,
         oc8051_ram_top1_oc8051_idata_n4562,
         oc8051_ram_top1_oc8051_idata_n4561,
         oc8051_ram_top1_oc8051_idata_n4560,
         oc8051_ram_top1_oc8051_idata_n4559,
         oc8051_ram_top1_oc8051_idata_n4558,
         oc8051_ram_top1_oc8051_idata_n4557,
         oc8051_ram_top1_oc8051_idata_n4556,
         oc8051_ram_top1_oc8051_idata_n4555,
         oc8051_ram_top1_oc8051_idata_n4554,
         oc8051_ram_top1_oc8051_idata_n4553,
         oc8051_ram_top1_oc8051_idata_n4552,
         oc8051_ram_top1_oc8051_idata_n4551,
         oc8051_ram_top1_oc8051_idata_n4550,
         oc8051_ram_top1_oc8051_idata_n4549,
         oc8051_ram_top1_oc8051_idata_n4548,
         oc8051_ram_top1_oc8051_idata_n4547,
         oc8051_ram_top1_oc8051_idata_n4546,
         oc8051_ram_top1_oc8051_idata_n4545,
         oc8051_ram_top1_oc8051_idata_n4544,
         oc8051_ram_top1_oc8051_idata_n4543,
         oc8051_ram_top1_oc8051_idata_n4542,
         oc8051_ram_top1_oc8051_idata_n4541,
         oc8051_ram_top1_oc8051_idata_n4540,
         oc8051_ram_top1_oc8051_idata_n4539,
         oc8051_ram_top1_oc8051_idata_n4538,
         oc8051_ram_top1_oc8051_idata_n4537,
         oc8051_ram_top1_oc8051_idata_n4536,
         oc8051_ram_top1_oc8051_idata_n4535,
         oc8051_ram_top1_oc8051_idata_n4534,
         oc8051_ram_top1_oc8051_idata_n4533,
         oc8051_ram_top1_oc8051_idata_n4532,
         oc8051_ram_top1_oc8051_idata_n4531,
         oc8051_ram_top1_oc8051_idata_n2474,
         oc8051_ram_top1_oc8051_idata_n2473,
         oc8051_ram_top1_oc8051_idata_n2472,
         oc8051_ram_top1_oc8051_idata_n2471,
         oc8051_ram_top1_oc8051_idata_n2470,
         oc8051_ram_top1_oc8051_idata_n2469,
         oc8051_ram_top1_oc8051_idata_n2468,
         oc8051_ram_top1_oc8051_idata_n2467,
         oc8051_ram_top1_oc8051_idata_n2466,
         oc8051_ram_top1_oc8051_idata_n2465,
         oc8051_ram_top1_oc8051_idata_n2464,
         oc8051_ram_top1_oc8051_idata_n2463,
         oc8051_ram_top1_oc8051_idata_n2462,
         oc8051_ram_top1_oc8051_idata_n2461,
         oc8051_ram_top1_oc8051_idata_n2460,
         oc8051_ram_top1_oc8051_idata_n2459,
         oc8051_ram_top1_oc8051_idata_n2458,
         oc8051_ram_top1_oc8051_idata_n2457,
         oc8051_ram_top1_oc8051_idata_n2456,
         oc8051_ram_top1_oc8051_idata_n2455,
         oc8051_ram_top1_oc8051_idata_n2454,
         oc8051_ram_top1_oc8051_idata_n2453,
         oc8051_ram_top1_oc8051_idata_n2452,
         oc8051_ram_top1_oc8051_idata_n2451,
         oc8051_ram_top1_oc8051_idata_n2450,
         oc8051_ram_top1_oc8051_idata_n2449,
         oc8051_ram_top1_oc8051_idata_n2448,
         oc8051_ram_top1_oc8051_idata_n2447,
         oc8051_ram_top1_oc8051_idata_n2446,
         oc8051_ram_top1_oc8051_idata_n2445,
         oc8051_ram_top1_oc8051_idata_n2444,
         oc8051_ram_top1_oc8051_idata_n2443,
         oc8051_ram_top1_oc8051_idata_n2442,
         oc8051_ram_top1_oc8051_idata_n2441,
         oc8051_ram_top1_oc8051_idata_n2440,
         oc8051_ram_top1_oc8051_idata_n2439,
         oc8051_ram_top1_oc8051_idata_n2438,
         oc8051_ram_top1_oc8051_idata_n2437,
         oc8051_ram_top1_oc8051_idata_n2436,
         oc8051_ram_top1_oc8051_idata_n2435,
         oc8051_ram_top1_oc8051_idata_n2434,
         oc8051_ram_top1_oc8051_idata_n2433,
         oc8051_ram_top1_oc8051_idata_n2432,
         oc8051_ram_top1_oc8051_idata_n2431,
         oc8051_ram_top1_oc8051_idata_n2430,
         oc8051_ram_top1_oc8051_idata_n2429,
         oc8051_ram_top1_oc8051_idata_n2428,
         oc8051_ram_top1_oc8051_idata_n2427,
         oc8051_ram_top1_oc8051_idata_n2426,
         oc8051_ram_top1_oc8051_idata_n2425,
         oc8051_ram_top1_oc8051_idata_n2424,
         oc8051_ram_top1_oc8051_idata_n2423,
         oc8051_ram_top1_oc8051_idata_n2422,
         oc8051_ram_top1_oc8051_idata_n2421,
         oc8051_ram_top1_oc8051_idata_n2420,
         oc8051_ram_top1_oc8051_idata_n2419,
         oc8051_ram_top1_oc8051_idata_n2418,
         oc8051_ram_top1_oc8051_idata_n2417,
         oc8051_ram_top1_oc8051_idata_n2416,
         oc8051_ram_top1_oc8051_idata_n2415,
         oc8051_ram_top1_oc8051_idata_n2414,
         oc8051_ram_top1_oc8051_idata_n2413,
         oc8051_ram_top1_oc8051_idata_n2412,
         oc8051_ram_top1_oc8051_idata_n2411,
         oc8051_ram_top1_oc8051_idata_n2410,
         oc8051_ram_top1_oc8051_idata_n2409,
         oc8051_ram_top1_oc8051_idata_n2408,
         oc8051_ram_top1_oc8051_idata_n2407,
         oc8051_ram_top1_oc8051_idata_n2406,
         oc8051_ram_top1_oc8051_idata_n2405,
         oc8051_ram_top1_oc8051_idata_n2404,
         oc8051_ram_top1_oc8051_idata_n2403,
         oc8051_ram_top1_oc8051_idata_n2402,
         oc8051_ram_top1_oc8051_idata_n2401,
         oc8051_ram_top1_oc8051_idata_n2400,
         oc8051_ram_top1_oc8051_idata_n2399,
         oc8051_ram_top1_oc8051_idata_n2398,
         oc8051_ram_top1_oc8051_idata_n2397,
         oc8051_ram_top1_oc8051_idata_n2396,
         oc8051_ram_top1_oc8051_idata_n2395,
         oc8051_ram_top1_oc8051_idata_n2394,
         oc8051_ram_top1_oc8051_idata_n2393,
         oc8051_ram_top1_oc8051_idata_n2392,
         oc8051_ram_top1_oc8051_idata_n2391,
         oc8051_ram_top1_oc8051_idata_n2390,
         oc8051_ram_top1_oc8051_idata_n2389,
         oc8051_ram_top1_oc8051_idata_n2388,
         oc8051_ram_top1_oc8051_idata_n2387,
         oc8051_ram_top1_oc8051_idata_n2386,
         oc8051_ram_top1_oc8051_idata_n2385,
         oc8051_ram_top1_oc8051_idata_n2384,
         oc8051_ram_top1_oc8051_idata_n2383,
         oc8051_ram_top1_oc8051_idata_n2382,
         oc8051_ram_top1_oc8051_idata_n2381,
         oc8051_ram_top1_oc8051_idata_n2380,
         oc8051_ram_top1_oc8051_idata_n2379,
         oc8051_ram_top1_oc8051_idata_n2378,
         oc8051_ram_top1_oc8051_idata_n2377,
         oc8051_ram_top1_oc8051_idata_n2376,
         oc8051_ram_top1_oc8051_idata_n2375,
         oc8051_ram_top1_oc8051_idata_n2374,
         oc8051_ram_top1_oc8051_idata_n2373,
         oc8051_ram_top1_oc8051_idata_n2372,
         oc8051_ram_top1_oc8051_idata_n2371,
         oc8051_ram_top1_oc8051_idata_n2370,
         oc8051_ram_top1_oc8051_idata_n2369,
         oc8051_ram_top1_oc8051_idata_n2368,
         oc8051_ram_top1_oc8051_idata_n2367,
         oc8051_ram_top1_oc8051_idata_n2366,
         oc8051_ram_top1_oc8051_idata_n2365,
         oc8051_ram_top1_oc8051_idata_n2364,
         oc8051_ram_top1_oc8051_idata_n2363,
         oc8051_ram_top1_oc8051_idata_n2362,
         oc8051_ram_top1_oc8051_idata_n2361,
         oc8051_ram_top1_oc8051_idata_n2360,
         oc8051_ram_top1_oc8051_idata_n2359,
         oc8051_ram_top1_oc8051_idata_n2358,
         oc8051_ram_top1_oc8051_idata_n2357,
         oc8051_ram_top1_oc8051_idata_n2356,
         oc8051_ram_top1_oc8051_idata_n2355,
         oc8051_ram_top1_oc8051_idata_n2354,
         oc8051_ram_top1_oc8051_idata_n2353,
         oc8051_ram_top1_oc8051_idata_n2352,
         oc8051_ram_top1_oc8051_idata_n2351,
         oc8051_ram_top1_oc8051_idata_n2350,
         oc8051_ram_top1_oc8051_idata_n2349,
         oc8051_ram_top1_oc8051_idata_n2348,
         oc8051_ram_top1_oc8051_idata_n2347,
         oc8051_ram_top1_oc8051_idata_n2346,
         oc8051_ram_top1_oc8051_idata_n2345,
         oc8051_ram_top1_oc8051_idata_n2344,
         oc8051_ram_top1_oc8051_idata_n2343,
         oc8051_ram_top1_oc8051_idata_n2342,
         oc8051_ram_top1_oc8051_idata_n2341,
         oc8051_ram_top1_oc8051_idata_n2340,
         oc8051_ram_top1_oc8051_idata_n2339,
         oc8051_ram_top1_oc8051_idata_n2338,
         oc8051_ram_top1_oc8051_idata_n2337,
         oc8051_ram_top1_oc8051_idata_n2336,
         oc8051_ram_top1_oc8051_idata_n2335,
         oc8051_ram_top1_oc8051_idata_n2334,
         oc8051_ram_top1_oc8051_idata_n2333,
         oc8051_ram_top1_oc8051_idata_n2332,
         oc8051_ram_top1_oc8051_idata_n2331,
         oc8051_ram_top1_oc8051_idata_n2330,
         oc8051_ram_top1_oc8051_idata_n2329,
         oc8051_ram_top1_oc8051_idata_n2328,
         oc8051_ram_top1_oc8051_idata_n2327,
         oc8051_ram_top1_oc8051_idata_n2326,
         oc8051_ram_top1_oc8051_idata_n2325,
         oc8051_ram_top1_oc8051_idata_n2324,
         oc8051_ram_top1_oc8051_idata_n2323,
         oc8051_ram_top1_oc8051_idata_n2322,
         oc8051_ram_top1_oc8051_idata_n2321,
         oc8051_ram_top1_oc8051_idata_n2320,
         oc8051_ram_top1_oc8051_idata_n2319,
         oc8051_ram_top1_oc8051_idata_n2318,
         oc8051_ram_top1_oc8051_idata_n2317,
         oc8051_ram_top1_oc8051_idata_n2316,
         oc8051_ram_top1_oc8051_idata_n2315,
         oc8051_ram_top1_oc8051_idata_n2314,
         oc8051_ram_top1_oc8051_idata_n2313,
         oc8051_ram_top1_oc8051_idata_n2312,
         oc8051_ram_top1_oc8051_idata_n2311,
         oc8051_ram_top1_oc8051_idata_n2310,
         oc8051_ram_top1_oc8051_idata_n2309,
         oc8051_ram_top1_oc8051_idata_n2308,
         oc8051_ram_top1_oc8051_idata_n2307,
         oc8051_ram_top1_oc8051_idata_n2306,
         oc8051_ram_top1_oc8051_idata_n2305,
         oc8051_ram_top1_oc8051_idata_n2304,
         oc8051_ram_top1_oc8051_idata_n2303,
         oc8051_ram_top1_oc8051_idata_n2302,
         oc8051_ram_top1_oc8051_idata_n2301,
         oc8051_ram_top1_oc8051_idata_n2300,
         oc8051_ram_top1_oc8051_idata_n2299,
         oc8051_ram_top1_oc8051_idata_n2298,
         oc8051_ram_top1_oc8051_idata_n2297,
         oc8051_ram_top1_oc8051_idata_n2296,
         oc8051_ram_top1_oc8051_idata_n2295,
         oc8051_ram_top1_oc8051_idata_n2294,
         oc8051_ram_top1_oc8051_idata_n2293,
         oc8051_ram_top1_oc8051_idata_n2292,
         oc8051_ram_top1_oc8051_idata_n2291,
         oc8051_ram_top1_oc8051_idata_n2290,
         oc8051_ram_top1_oc8051_idata_n2289,
         oc8051_ram_top1_oc8051_idata_n2288,
         oc8051_ram_top1_oc8051_idata_n2287,
         oc8051_ram_top1_oc8051_idata_n2286,
         oc8051_ram_top1_oc8051_idata_n2285,
         oc8051_ram_top1_oc8051_idata_n2284,
         oc8051_ram_top1_oc8051_idata_n2283,
         oc8051_ram_top1_oc8051_idata_n2282,
         oc8051_ram_top1_oc8051_idata_n2281,
         oc8051_ram_top1_oc8051_idata_n2280,
         oc8051_ram_top1_oc8051_idata_n2279,
         oc8051_ram_top1_oc8051_idata_n2278,
         oc8051_ram_top1_oc8051_idata_n2277,
         oc8051_ram_top1_oc8051_idata_n2276,
         oc8051_ram_top1_oc8051_idata_n2275,
         oc8051_ram_top1_oc8051_idata_n2274,
         oc8051_ram_top1_oc8051_idata_n2273,
         oc8051_ram_top1_oc8051_idata_n2272,
         oc8051_ram_top1_oc8051_idata_n2271,
         oc8051_ram_top1_oc8051_idata_n2270,
         oc8051_ram_top1_oc8051_idata_n2269,
         oc8051_ram_top1_oc8051_idata_n2268,
         oc8051_ram_top1_oc8051_idata_n2267,
         oc8051_ram_top1_oc8051_idata_n2266,
         oc8051_ram_top1_oc8051_idata_n2265,
         oc8051_ram_top1_oc8051_idata_n2264,
         oc8051_ram_top1_oc8051_idata_n2263,
         oc8051_ram_top1_oc8051_idata_n2262,
         oc8051_ram_top1_oc8051_idata_n2261,
         oc8051_ram_top1_oc8051_idata_n2260,
         oc8051_ram_top1_oc8051_idata_n2259,
         oc8051_ram_top1_oc8051_idata_n2258,
         oc8051_ram_top1_oc8051_idata_n2257,
         oc8051_ram_top1_oc8051_idata_n2256,
         oc8051_ram_top1_oc8051_idata_n2255,
         oc8051_ram_top1_oc8051_idata_n2254,
         oc8051_ram_top1_oc8051_idata_n2253,
         oc8051_ram_top1_oc8051_idata_n2252,
         oc8051_ram_top1_oc8051_idata_n2251,
         oc8051_ram_top1_oc8051_idata_n2250,
         oc8051_ram_top1_oc8051_idata_n2249,
         oc8051_ram_top1_oc8051_idata_n2248,
         oc8051_ram_top1_oc8051_idata_n2247,
         oc8051_ram_top1_oc8051_idata_n2246,
         oc8051_ram_top1_oc8051_idata_n2245,
         oc8051_ram_top1_oc8051_idata_n2244,
         oc8051_ram_top1_oc8051_idata_n2243,
         oc8051_ram_top1_oc8051_idata_n2242,
         oc8051_ram_top1_oc8051_idata_n2241,
         oc8051_ram_top1_oc8051_idata_n2240,
         oc8051_ram_top1_oc8051_idata_n2239,
         oc8051_ram_top1_oc8051_idata_n2238,
         oc8051_ram_top1_oc8051_idata_n2237,
         oc8051_ram_top1_oc8051_idata_n2236,
         oc8051_ram_top1_oc8051_idata_n2235,
         oc8051_ram_top1_oc8051_idata_n2234,
         oc8051_ram_top1_oc8051_idata_n2233,
         oc8051_ram_top1_oc8051_idata_n2232,
         oc8051_ram_top1_oc8051_idata_n2231,
         oc8051_ram_top1_oc8051_idata_n2230,
         oc8051_ram_top1_oc8051_idata_n2229,
         oc8051_ram_top1_oc8051_idata_n2228,
         oc8051_ram_top1_oc8051_idata_n2227,
         oc8051_ram_top1_oc8051_idata_n2226,
         oc8051_ram_top1_oc8051_idata_n2225,
         oc8051_ram_top1_oc8051_idata_n2224,
         oc8051_ram_top1_oc8051_idata_n2223,
         oc8051_ram_top1_oc8051_idata_n2222,
         oc8051_ram_top1_oc8051_idata_n2221,
         oc8051_ram_top1_oc8051_idata_n2220,
         oc8051_ram_top1_oc8051_idata_n2219,
         oc8051_ram_top1_oc8051_idata_n2218,
         oc8051_ram_top1_oc8051_idata_n2217,
         oc8051_ram_top1_oc8051_idata_n2216,
         oc8051_ram_top1_oc8051_idata_n2215,
         oc8051_ram_top1_oc8051_idata_n2214,
         oc8051_ram_top1_oc8051_idata_n2213,
         oc8051_ram_top1_oc8051_idata_n2212,
         oc8051_ram_top1_oc8051_idata_n2211,
         oc8051_ram_top1_oc8051_idata_n2210,
         oc8051_ram_top1_oc8051_idata_n2209,
         oc8051_ram_top1_oc8051_idata_n2208,
         oc8051_ram_top1_oc8051_idata_n2207,
         oc8051_ram_top1_oc8051_idata_n2206,
         oc8051_ram_top1_oc8051_idata_n2205,
         oc8051_ram_top1_oc8051_idata_n2204,
         oc8051_ram_top1_oc8051_idata_n2203,
         oc8051_ram_top1_oc8051_idata_n2202,
         oc8051_ram_top1_oc8051_idata_n2201,
         oc8051_ram_top1_oc8051_idata_n2200,
         oc8051_ram_top1_oc8051_idata_n2199,
         oc8051_ram_top1_oc8051_idata_n2198,
         oc8051_ram_top1_oc8051_idata_n2197,
         oc8051_ram_top1_oc8051_idata_n2196,
         oc8051_ram_top1_oc8051_idata_n2195,
         oc8051_ram_top1_oc8051_idata_n2194,
         oc8051_ram_top1_oc8051_idata_n2193,
         oc8051_ram_top1_oc8051_idata_n2192,
         oc8051_ram_top1_oc8051_idata_n2191,
         oc8051_ram_top1_oc8051_idata_n2190,
         oc8051_ram_top1_oc8051_idata_n2189,
         oc8051_ram_top1_oc8051_idata_n2188,
         oc8051_ram_top1_oc8051_idata_n2187,
         oc8051_ram_top1_oc8051_idata_n2186,
         oc8051_ram_top1_oc8051_idata_n2185,
         oc8051_ram_top1_oc8051_idata_n2184,
         oc8051_ram_top1_oc8051_idata_n2183,
         oc8051_ram_top1_oc8051_idata_n2182,
         oc8051_ram_top1_oc8051_idata_n2181,
         oc8051_ram_top1_oc8051_idata_n2180,
         oc8051_ram_top1_oc8051_idata_n2179,
         oc8051_ram_top1_oc8051_idata_n2178,
         oc8051_ram_top1_oc8051_idata_n2177,
         oc8051_ram_top1_oc8051_idata_n2176,
         oc8051_ram_top1_oc8051_idata_n2175,
         oc8051_ram_top1_oc8051_idata_n2174,
         oc8051_ram_top1_oc8051_idata_n2173,
         oc8051_ram_top1_oc8051_idata_n2172,
         oc8051_ram_top1_oc8051_idata_n2171,
         oc8051_ram_top1_oc8051_idata_n2170,
         oc8051_ram_top1_oc8051_idata_n2169,
         oc8051_ram_top1_oc8051_idata_n2168,
         oc8051_ram_top1_oc8051_idata_n2167,
         oc8051_ram_top1_oc8051_idata_n2166,
         oc8051_ram_top1_oc8051_idata_n2165,
         oc8051_ram_top1_oc8051_idata_n2164,
         oc8051_ram_top1_oc8051_idata_n2163,
         oc8051_ram_top1_oc8051_idata_n2162,
         oc8051_ram_top1_oc8051_idata_n2161,
         oc8051_ram_top1_oc8051_idata_n2160,
         oc8051_ram_top1_oc8051_idata_n2159,
         oc8051_ram_top1_oc8051_idata_n2158,
         oc8051_ram_top1_oc8051_idata_n2157,
         oc8051_ram_top1_oc8051_idata_n2156,
         oc8051_ram_top1_oc8051_idata_n2155,
         oc8051_ram_top1_oc8051_idata_n2154,
         oc8051_ram_top1_oc8051_idata_n2153,
         oc8051_ram_top1_oc8051_idata_n2152,
         oc8051_ram_top1_oc8051_idata_n2151,
         oc8051_ram_top1_oc8051_idata_n2150,
         oc8051_ram_top1_oc8051_idata_n2149,
         oc8051_ram_top1_oc8051_idata_n2148,
         oc8051_ram_top1_oc8051_idata_n2147,
         oc8051_ram_top1_oc8051_idata_n2146,
         oc8051_ram_top1_oc8051_idata_n2145,
         oc8051_ram_top1_oc8051_idata_n2144,
         oc8051_ram_top1_oc8051_idata_n2143,
         oc8051_ram_top1_oc8051_idata_n2142,
         oc8051_ram_top1_oc8051_idata_n2141,
         oc8051_ram_top1_oc8051_idata_n2140,
         oc8051_ram_top1_oc8051_idata_n2139,
         oc8051_ram_top1_oc8051_idata_n2138,
         oc8051_ram_top1_oc8051_idata_n2137,
         oc8051_ram_top1_oc8051_idata_n2136,
         oc8051_ram_top1_oc8051_idata_n2135,
         oc8051_ram_top1_oc8051_idata_n2134,
         oc8051_ram_top1_oc8051_idata_n2133,
         oc8051_ram_top1_oc8051_idata_n2132,
         oc8051_ram_top1_oc8051_idata_n2131,
         oc8051_ram_top1_oc8051_idata_n2130,
         oc8051_ram_top1_oc8051_idata_n2129,
         oc8051_ram_top1_oc8051_idata_n2128,
         oc8051_ram_top1_oc8051_idata_n2127,
         oc8051_ram_top1_oc8051_idata_n2126,
         oc8051_ram_top1_oc8051_idata_n2125,
         oc8051_ram_top1_oc8051_idata_n2124,
         oc8051_ram_top1_oc8051_idata_n2123,
         oc8051_ram_top1_oc8051_idata_n2122,
         oc8051_ram_top1_oc8051_idata_n2121,
         oc8051_ram_top1_oc8051_idata_n2120,
         oc8051_ram_top1_oc8051_idata_n2119,
         oc8051_ram_top1_oc8051_idata_n2118,
         oc8051_ram_top1_oc8051_idata_n2117,
         oc8051_ram_top1_oc8051_idata_n2116,
         oc8051_ram_top1_oc8051_idata_n2115,
         oc8051_ram_top1_oc8051_idata_n2114,
         oc8051_ram_top1_oc8051_idata_n2113,
         oc8051_ram_top1_oc8051_idata_n2112,
         oc8051_ram_top1_oc8051_idata_n2111,
         oc8051_ram_top1_oc8051_idata_n2110,
         oc8051_ram_top1_oc8051_idata_n2109,
         oc8051_ram_top1_oc8051_idata_n2108,
         oc8051_ram_top1_oc8051_idata_n2107,
         oc8051_ram_top1_oc8051_idata_n2106,
         oc8051_ram_top1_oc8051_idata_n2105,
         oc8051_ram_top1_oc8051_idata_n2104,
         oc8051_ram_top1_oc8051_idata_n2103,
         oc8051_ram_top1_oc8051_idata_n2102,
         oc8051_ram_top1_oc8051_idata_n2101,
         oc8051_ram_top1_oc8051_idata_n2100,
         oc8051_ram_top1_oc8051_idata_n2099,
         oc8051_ram_top1_oc8051_idata_n2098,
         oc8051_ram_top1_oc8051_idata_n2097,
         oc8051_ram_top1_oc8051_idata_n2096,
         oc8051_ram_top1_oc8051_idata_n2095,
         oc8051_ram_top1_oc8051_idata_n2094,
         oc8051_ram_top1_oc8051_idata_n2093,
         oc8051_ram_top1_oc8051_idata_n2092,
         oc8051_ram_top1_oc8051_idata_n2091,
         oc8051_ram_top1_oc8051_idata_n2090,
         oc8051_ram_top1_oc8051_idata_n2089,
         oc8051_ram_top1_oc8051_idata_n2088,
         oc8051_ram_top1_oc8051_idata_n2087,
         oc8051_ram_top1_oc8051_idata_n2086,
         oc8051_ram_top1_oc8051_idata_n2085,
         oc8051_ram_top1_oc8051_idata_n2084,
         oc8051_ram_top1_oc8051_idata_n2083,
         oc8051_ram_top1_oc8051_idata_n2082,
         oc8051_ram_top1_oc8051_idata_n2081,
         oc8051_ram_top1_oc8051_idata_n2080,
         oc8051_ram_top1_oc8051_idata_n2079,
         oc8051_ram_top1_oc8051_idata_n2078,
         oc8051_ram_top1_oc8051_idata_n2077,
         oc8051_ram_top1_oc8051_idata_n2076,
         oc8051_ram_top1_oc8051_idata_n2075,
         oc8051_ram_top1_oc8051_idata_n2074,
         oc8051_ram_top1_oc8051_idata_n2073,
         oc8051_ram_top1_oc8051_idata_n2072,
         oc8051_ram_top1_oc8051_idata_n2071,
         oc8051_ram_top1_oc8051_idata_n2070,
         oc8051_ram_top1_oc8051_idata_n2069,
         oc8051_ram_top1_oc8051_idata_n2068,
         oc8051_ram_top1_oc8051_idata_n2067,
         oc8051_ram_top1_oc8051_idata_n2066,
         oc8051_ram_top1_oc8051_idata_n2065,
         oc8051_ram_top1_oc8051_idata_n2064,
         oc8051_ram_top1_oc8051_idata_n2063,
         oc8051_ram_top1_oc8051_idata_n2062,
         oc8051_ram_top1_oc8051_idata_n2061,
         oc8051_ram_top1_oc8051_idata_n2060,
         oc8051_ram_top1_oc8051_idata_n2059,
         oc8051_ram_top1_oc8051_idata_n2058,
         oc8051_ram_top1_oc8051_idata_n2057,
         oc8051_ram_top1_oc8051_idata_n2056,
         oc8051_ram_top1_oc8051_idata_n2055,
         oc8051_ram_top1_oc8051_idata_n2054,
         oc8051_ram_top1_oc8051_idata_n2053,
         oc8051_ram_top1_oc8051_idata_n2052,
         oc8051_ram_top1_oc8051_idata_n2051,
         oc8051_ram_top1_oc8051_idata_n2050,
         oc8051_ram_top1_oc8051_idata_n2049,
         oc8051_ram_top1_oc8051_idata_n2048,
         oc8051_ram_top1_oc8051_idata_n2047,
         oc8051_ram_top1_oc8051_idata_n2046,
         oc8051_ram_top1_oc8051_idata_n2045,
         oc8051_ram_top1_oc8051_idata_n2044,
         oc8051_ram_top1_oc8051_idata_n2043,
         oc8051_ram_top1_oc8051_idata_n2042,
         oc8051_ram_top1_oc8051_idata_n2041,
         oc8051_ram_top1_oc8051_idata_n2040,
         oc8051_ram_top1_oc8051_idata_n2039,
         oc8051_ram_top1_oc8051_idata_n2038,
         oc8051_ram_top1_oc8051_idata_n2037,
         oc8051_ram_top1_oc8051_idata_n2036,
         oc8051_ram_top1_oc8051_idata_n2035,
         oc8051_ram_top1_oc8051_idata_n2034,
         oc8051_ram_top1_oc8051_idata_n2033,
         oc8051_ram_top1_oc8051_idata_n2032,
         oc8051_ram_top1_oc8051_idata_n2031,
         oc8051_ram_top1_oc8051_idata_n2030,
         oc8051_ram_top1_oc8051_idata_n2029,
         oc8051_ram_top1_oc8051_idata_n2028,
         oc8051_ram_top1_oc8051_idata_n2027,
         oc8051_ram_top1_oc8051_idata_n2026,
         oc8051_ram_top1_oc8051_idata_n2025,
         oc8051_ram_top1_oc8051_idata_n2024,
         oc8051_ram_top1_oc8051_idata_n2023,
         oc8051_ram_top1_oc8051_idata_n2022,
         oc8051_ram_top1_oc8051_idata_n2021,
         oc8051_ram_top1_oc8051_idata_n2020,
         oc8051_ram_top1_oc8051_idata_n2019,
         oc8051_ram_top1_oc8051_idata_n2018,
         oc8051_ram_top1_oc8051_idata_n2017,
         oc8051_ram_top1_oc8051_idata_n2016,
         oc8051_ram_top1_oc8051_idata_n2015,
         oc8051_ram_top1_oc8051_idata_n2014,
         oc8051_ram_top1_oc8051_idata_n2013,
         oc8051_ram_top1_oc8051_idata_n2012,
         oc8051_ram_top1_oc8051_idata_n2011,
         oc8051_ram_top1_oc8051_idata_n2010,
         oc8051_ram_top1_oc8051_idata_n2009,
         oc8051_ram_top1_oc8051_idata_n2008,
         oc8051_ram_top1_oc8051_idata_n2007,
         oc8051_ram_top1_oc8051_idata_n2006,
         oc8051_ram_top1_oc8051_idata_n2005,
         oc8051_ram_top1_oc8051_idata_n2004,
         oc8051_ram_top1_oc8051_idata_n2003,
         oc8051_ram_top1_oc8051_idata_n2002,
         oc8051_ram_top1_oc8051_idata_n2001,
         oc8051_ram_top1_oc8051_idata_n2000,
         oc8051_ram_top1_oc8051_idata_n1999,
         oc8051_ram_top1_oc8051_idata_n1998,
         oc8051_ram_top1_oc8051_idata_n1997,
         oc8051_ram_top1_oc8051_idata_n1996,
         oc8051_ram_top1_oc8051_idata_n1995,
         oc8051_ram_top1_oc8051_idata_n1994,
         oc8051_ram_top1_oc8051_idata_n1993,
         oc8051_ram_top1_oc8051_idata_n1992,
         oc8051_ram_top1_oc8051_idata_n1991,
         oc8051_ram_top1_oc8051_idata_n1990,
         oc8051_ram_top1_oc8051_idata_n1989,
         oc8051_ram_top1_oc8051_idata_n1988,
         oc8051_ram_top1_oc8051_idata_n1987,
         oc8051_ram_top1_oc8051_idata_n1986,
         oc8051_ram_top1_oc8051_idata_n1985,
         oc8051_ram_top1_oc8051_idata_n1984,
         oc8051_ram_top1_oc8051_idata_n1983,
         oc8051_ram_top1_oc8051_idata_n1982,
         oc8051_ram_top1_oc8051_idata_n1981,
         oc8051_ram_top1_oc8051_idata_n1980,
         oc8051_ram_top1_oc8051_idata_n1979,
         oc8051_ram_top1_oc8051_idata_n1978,
         oc8051_ram_top1_oc8051_idata_n1977,
         oc8051_ram_top1_oc8051_idata_n1976,
         oc8051_ram_top1_oc8051_idata_n1975,
         oc8051_ram_top1_oc8051_idata_n1974,
         oc8051_ram_top1_oc8051_idata_n1973,
         oc8051_ram_top1_oc8051_idata_n1972,
         oc8051_ram_top1_oc8051_idata_n1971,
         oc8051_ram_top1_oc8051_idata_n1970,
         oc8051_ram_top1_oc8051_idata_n1969,
         oc8051_ram_top1_oc8051_idata_n1968,
         oc8051_ram_top1_oc8051_idata_n1967,
         oc8051_ram_top1_oc8051_idata_n1966,
         oc8051_ram_top1_oc8051_idata_n1965,
         oc8051_ram_top1_oc8051_idata_n1964,
         oc8051_ram_top1_oc8051_idata_n1963,
         oc8051_ram_top1_oc8051_idata_n1962,
         oc8051_ram_top1_oc8051_idata_n1961,
         oc8051_ram_top1_oc8051_idata_n1960,
         oc8051_ram_top1_oc8051_idata_n1959,
         oc8051_ram_top1_oc8051_idata_n1958,
         oc8051_ram_top1_oc8051_idata_n1957,
         oc8051_ram_top1_oc8051_idata_n1956,
         oc8051_ram_top1_oc8051_idata_n1955,
         oc8051_ram_top1_oc8051_idata_n1954,
         oc8051_ram_top1_oc8051_idata_n1953,
         oc8051_ram_top1_oc8051_idata_n1952,
         oc8051_ram_top1_oc8051_idata_n1951,
         oc8051_ram_top1_oc8051_idata_n1950,
         oc8051_ram_top1_oc8051_idata_n1949,
         oc8051_ram_top1_oc8051_idata_n1948,
         oc8051_ram_top1_oc8051_idata_n1947,
         oc8051_ram_top1_oc8051_idata_n1946,
         oc8051_ram_top1_oc8051_idata_n1945,
         oc8051_ram_top1_oc8051_idata_n1944,
         oc8051_ram_top1_oc8051_idata_n1943,
         oc8051_ram_top1_oc8051_idata_n1942,
         oc8051_ram_top1_oc8051_idata_n1941,
         oc8051_ram_top1_oc8051_idata_n1940,
         oc8051_ram_top1_oc8051_idata_n1939,
         oc8051_ram_top1_oc8051_idata_n1938,
         oc8051_ram_top1_oc8051_idata_n1937,
         oc8051_ram_top1_oc8051_idata_n1936,
         oc8051_ram_top1_oc8051_idata_n1935,
         oc8051_ram_top1_oc8051_idata_n1934,
         oc8051_ram_top1_oc8051_idata_n1933,
         oc8051_ram_top1_oc8051_idata_n1932,
         oc8051_ram_top1_oc8051_idata_n1931,
         oc8051_ram_top1_oc8051_idata_n1930,
         oc8051_ram_top1_oc8051_idata_n1929,
         oc8051_ram_top1_oc8051_idata_n1928,
         oc8051_ram_top1_oc8051_idata_n1927,
         oc8051_ram_top1_oc8051_idata_n1926,
         oc8051_ram_top1_oc8051_idata_n1925,
         oc8051_ram_top1_oc8051_idata_n1924,
         oc8051_ram_top1_oc8051_idata_n1923,
         oc8051_ram_top1_oc8051_idata_n1922,
         oc8051_ram_top1_oc8051_idata_n1921,
         oc8051_ram_top1_oc8051_idata_n1920,
         oc8051_ram_top1_oc8051_idata_n1919,
         oc8051_ram_top1_oc8051_idata_n1918,
         oc8051_ram_top1_oc8051_idata_n1917,
         oc8051_ram_top1_oc8051_idata_n1916,
         oc8051_ram_top1_oc8051_idata_n1915,
         oc8051_ram_top1_oc8051_idata_n1914,
         oc8051_ram_top1_oc8051_idata_n1913,
         oc8051_ram_top1_oc8051_idata_n1912,
         oc8051_ram_top1_oc8051_idata_n1911,
         oc8051_ram_top1_oc8051_idata_n1910,
         oc8051_ram_top1_oc8051_idata_n1909,
         oc8051_ram_top1_oc8051_idata_n1908,
         oc8051_ram_top1_oc8051_idata_n1907,
         oc8051_ram_top1_oc8051_idata_n1906,
         oc8051_ram_top1_oc8051_idata_n1905,
         oc8051_ram_top1_oc8051_idata_n1904,
         oc8051_ram_top1_oc8051_idata_n1903,
         oc8051_ram_top1_oc8051_idata_n1902,
         oc8051_ram_top1_oc8051_idata_n1901,
         oc8051_ram_top1_oc8051_idata_n1900,
         oc8051_ram_top1_oc8051_idata_n1899,
         oc8051_ram_top1_oc8051_idata_n1898,
         oc8051_ram_top1_oc8051_idata_n1897,
         oc8051_ram_top1_oc8051_idata_n1896,
         oc8051_ram_top1_oc8051_idata_n1895,
         oc8051_ram_top1_oc8051_idata_n1894,
         oc8051_ram_top1_oc8051_idata_n1893,
         oc8051_ram_top1_oc8051_idata_n1892,
         oc8051_ram_top1_oc8051_idata_n1891,
         oc8051_ram_top1_oc8051_idata_n1890,
         oc8051_ram_top1_oc8051_idata_n1889,
         oc8051_ram_top1_oc8051_idata_n1888,
         oc8051_ram_top1_oc8051_idata_n1887,
         oc8051_ram_top1_oc8051_idata_n1886,
         oc8051_ram_top1_oc8051_idata_n1885,
         oc8051_ram_top1_oc8051_idata_n1884,
         oc8051_ram_top1_oc8051_idata_n1883,
         oc8051_ram_top1_oc8051_idata_n1882,
         oc8051_ram_top1_oc8051_idata_n1881,
         oc8051_ram_top1_oc8051_idata_n1880,
         oc8051_ram_top1_oc8051_idata_n1879,
         oc8051_ram_top1_oc8051_idata_n1878,
         oc8051_ram_top1_oc8051_idata_n1877,
         oc8051_ram_top1_oc8051_idata_n1876,
         oc8051_ram_top1_oc8051_idata_n1875,
         oc8051_ram_top1_oc8051_idata_n1874,
         oc8051_ram_top1_oc8051_idata_n1873,
         oc8051_ram_top1_oc8051_idata_n1872,
         oc8051_ram_top1_oc8051_idata_n1871,
         oc8051_ram_top1_oc8051_idata_n1870,
         oc8051_ram_top1_oc8051_idata_n1869,
         oc8051_ram_top1_oc8051_idata_n1868,
         oc8051_ram_top1_oc8051_idata_n1867,
         oc8051_ram_top1_oc8051_idata_n1866,
         oc8051_ram_top1_oc8051_idata_n1865,
         oc8051_ram_top1_oc8051_idata_n1864,
         oc8051_ram_top1_oc8051_idata_n1863,
         oc8051_ram_top1_oc8051_idata_n1862,
         oc8051_ram_top1_oc8051_idata_n1861,
         oc8051_ram_top1_oc8051_idata_n1860,
         oc8051_ram_top1_oc8051_idata_n1859,
         oc8051_ram_top1_oc8051_idata_n1858,
         oc8051_ram_top1_oc8051_idata_n1857,
         oc8051_ram_top1_oc8051_idata_n1856,
         oc8051_ram_top1_oc8051_idata_n1855,
         oc8051_ram_top1_oc8051_idata_n1854,
         oc8051_ram_top1_oc8051_idata_n1853,
         oc8051_ram_top1_oc8051_idata_n1852,
         oc8051_ram_top1_oc8051_idata_n1851,
         oc8051_ram_top1_oc8051_idata_n1850,
         oc8051_ram_top1_oc8051_idata_n1849,
         oc8051_ram_top1_oc8051_idata_n1848,
         oc8051_ram_top1_oc8051_idata_n1847,
         oc8051_ram_top1_oc8051_idata_n1846,
         oc8051_ram_top1_oc8051_idata_n1845,
         oc8051_ram_top1_oc8051_idata_n1844,
         oc8051_ram_top1_oc8051_idata_n1843,
         oc8051_ram_top1_oc8051_idata_n1842,
         oc8051_ram_top1_oc8051_idata_n1841,
         oc8051_ram_top1_oc8051_idata_n1840,
         oc8051_ram_top1_oc8051_idata_n1839,
         oc8051_ram_top1_oc8051_idata_n1838,
         oc8051_ram_top1_oc8051_idata_n1837,
         oc8051_ram_top1_oc8051_idata_n1836,
         oc8051_ram_top1_oc8051_idata_n1835,
         oc8051_ram_top1_oc8051_idata_n1834,
         oc8051_ram_top1_oc8051_idata_n1833,
         oc8051_ram_top1_oc8051_idata_n1832,
         oc8051_ram_top1_oc8051_idata_n1831,
         oc8051_ram_top1_oc8051_idata_n1830,
         oc8051_ram_top1_oc8051_idata_n1829,
         oc8051_ram_top1_oc8051_idata_n1828,
         oc8051_ram_top1_oc8051_idata_n1827,
         oc8051_ram_top1_oc8051_idata_n1826,
         oc8051_ram_top1_oc8051_idata_n1825,
         oc8051_ram_top1_oc8051_idata_n1824,
         oc8051_ram_top1_oc8051_idata_n1823,
         oc8051_ram_top1_oc8051_idata_n1822,
         oc8051_ram_top1_oc8051_idata_n1821,
         oc8051_ram_top1_oc8051_idata_n1820,
         oc8051_ram_top1_oc8051_idata_n1819,
         oc8051_ram_top1_oc8051_idata_n1818,
         oc8051_ram_top1_oc8051_idata_n1817,
         oc8051_ram_top1_oc8051_idata_n1816,
         oc8051_ram_top1_oc8051_idata_n1815,
         oc8051_ram_top1_oc8051_idata_n1814,
         oc8051_ram_top1_oc8051_idata_n1813,
         oc8051_ram_top1_oc8051_idata_n1812,
         oc8051_ram_top1_oc8051_idata_n1811,
         oc8051_ram_top1_oc8051_idata_n1810,
         oc8051_ram_top1_oc8051_idata_n1809,
         oc8051_ram_top1_oc8051_idata_n1808,
         oc8051_ram_top1_oc8051_idata_n1807,
         oc8051_ram_top1_oc8051_idata_n1806,
         oc8051_ram_top1_oc8051_idata_n1805,
         oc8051_ram_top1_oc8051_idata_n1804,
         oc8051_ram_top1_oc8051_idata_n1803,
         oc8051_ram_top1_oc8051_idata_n1802,
         oc8051_ram_top1_oc8051_idata_n1801,
         oc8051_ram_top1_oc8051_idata_n1800,
         oc8051_ram_top1_oc8051_idata_n1799,
         oc8051_ram_top1_oc8051_idata_n1798,
         oc8051_ram_top1_oc8051_idata_n1797,
         oc8051_ram_top1_oc8051_idata_n1796,
         oc8051_ram_top1_oc8051_idata_n1795,
         oc8051_ram_top1_oc8051_idata_n1794,
         oc8051_ram_top1_oc8051_idata_n1793,
         oc8051_ram_top1_oc8051_idata_n1792,
         oc8051_ram_top1_oc8051_idata_n1791,
         oc8051_ram_top1_oc8051_idata_n1790,
         oc8051_ram_top1_oc8051_idata_n1789,
         oc8051_ram_top1_oc8051_idata_n1788,
         oc8051_ram_top1_oc8051_idata_n1787,
         oc8051_ram_top1_oc8051_idata_n1786,
         oc8051_ram_top1_oc8051_idata_n1785,
         oc8051_ram_top1_oc8051_idata_n1784,
         oc8051_ram_top1_oc8051_idata_n1783,
         oc8051_ram_top1_oc8051_idata_n1782,
         oc8051_ram_top1_oc8051_idata_n1781,
         oc8051_ram_top1_oc8051_idata_n1780,
         oc8051_ram_top1_oc8051_idata_n1779,
         oc8051_ram_top1_oc8051_idata_n1778,
         oc8051_ram_top1_oc8051_idata_n1777,
         oc8051_ram_top1_oc8051_idata_n1776,
         oc8051_ram_top1_oc8051_idata_n1775,
         oc8051_ram_top1_oc8051_idata_n1774,
         oc8051_ram_top1_oc8051_idata_n1773,
         oc8051_ram_top1_oc8051_idata_n1772,
         oc8051_ram_top1_oc8051_idata_n1771,
         oc8051_ram_top1_oc8051_idata_n1770,
         oc8051_ram_top1_oc8051_idata_n1769,
         oc8051_ram_top1_oc8051_idata_n1768,
         oc8051_ram_top1_oc8051_idata_n1767,
         oc8051_ram_top1_oc8051_idata_n1766,
         oc8051_ram_top1_oc8051_idata_n1765,
         oc8051_ram_top1_oc8051_idata_n1764,
         oc8051_ram_top1_oc8051_idata_n1763,
         oc8051_ram_top1_oc8051_idata_n1762,
         oc8051_ram_top1_oc8051_idata_n1761,
         oc8051_ram_top1_oc8051_idata_n1760,
         oc8051_ram_top1_oc8051_idata_n1759,
         oc8051_ram_top1_oc8051_idata_n1758,
         oc8051_ram_top1_oc8051_idata_n1757,
         oc8051_ram_top1_oc8051_idata_n1756,
         oc8051_ram_top1_oc8051_idata_n1755,
         oc8051_ram_top1_oc8051_idata_n1754,
         oc8051_ram_top1_oc8051_idata_n1753,
         oc8051_ram_top1_oc8051_idata_n1752,
         oc8051_ram_top1_oc8051_idata_n1751,
         oc8051_ram_top1_oc8051_idata_n1750,
         oc8051_ram_top1_oc8051_idata_n1749,
         oc8051_ram_top1_oc8051_idata_n1748,
         oc8051_ram_top1_oc8051_idata_n1747,
         oc8051_ram_top1_oc8051_idata_n1746,
         oc8051_ram_top1_oc8051_idata_n1745,
         oc8051_ram_top1_oc8051_idata_n1744,
         oc8051_ram_top1_oc8051_idata_n1743,
         oc8051_ram_top1_oc8051_idata_n1742,
         oc8051_ram_top1_oc8051_idata_n1741,
         oc8051_ram_top1_oc8051_idata_n1740,
         oc8051_ram_top1_oc8051_idata_n1739,
         oc8051_ram_top1_oc8051_idata_n1738,
         oc8051_ram_top1_oc8051_idata_n1737,
         oc8051_ram_top1_oc8051_idata_n1736,
         oc8051_ram_top1_oc8051_idata_n1735,
         oc8051_ram_top1_oc8051_idata_n1734,
         oc8051_ram_top1_oc8051_idata_n1733,
         oc8051_ram_top1_oc8051_idata_n1732,
         oc8051_ram_top1_oc8051_idata_n1731,
         oc8051_ram_top1_oc8051_idata_n1730,
         oc8051_ram_top1_oc8051_idata_n1729,
         oc8051_ram_top1_oc8051_idata_n1728,
         oc8051_ram_top1_oc8051_idata_n1727,
         oc8051_ram_top1_oc8051_idata_n1726,
         oc8051_ram_top1_oc8051_idata_n1725,
         oc8051_ram_top1_oc8051_idata_n1724,
         oc8051_ram_top1_oc8051_idata_n1723,
         oc8051_ram_top1_oc8051_idata_n1722,
         oc8051_ram_top1_oc8051_idata_n1721,
         oc8051_ram_top1_oc8051_idata_n1720,
         oc8051_ram_top1_oc8051_idata_n1719,
         oc8051_ram_top1_oc8051_idata_n1718,
         oc8051_ram_top1_oc8051_idata_n1717,
         oc8051_ram_top1_oc8051_idata_n1716,
         oc8051_ram_top1_oc8051_idata_n1715,
         oc8051_ram_top1_oc8051_idata_n1714,
         oc8051_ram_top1_oc8051_idata_n1713,
         oc8051_ram_top1_oc8051_idata_n1712,
         oc8051_ram_top1_oc8051_idata_n1711,
         oc8051_ram_top1_oc8051_idata_n1710,
         oc8051_ram_top1_oc8051_idata_n1709,
         oc8051_ram_top1_oc8051_idata_n1708,
         oc8051_ram_top1_oc8051_idata_n1707,
         oc8051_ram_top1_oc8051_idata_n1706,
         oc8051_ram_top1_oc8051_idata_n1705,
         oc8051_ram_top1_oc8051_idata_n1704,
         oc8051_ram_top1_oc8051_idata_n1703,
         oc8051_ram_top1_oc8051_idata_n1702,
         oc8051_ram_top1_oc8051_idata_n1701,
         oc8051_ram_top1_oc8051_idata_n1700,
         oc8051_ram_top1_oc8051_idata_n1699,
         oc8051_ram_top1_oc8051_idata_n1698,
         oc8051_ram_top1_oc8051_idata_n1697,
         oc8051_ram_top1_oc8051_idata_n1696,
         oc8051_ram_top1_oc8051_idata_n1695,
         oc8051_ram_top1_oc8051_idata_n1694,
         oc8051_ram_top1_oc8051_idata_n1693,
         oc8051_ram_top1_oc8051_idata_n1692,
         oc8051_ram_top1_oc8051_idata_n1691,
         oc8051_ram_top1_oc8051_idata_n1690,
         oc8051_ram_top1_oc8051_idata_n1689,
         oc8051_ram_top1_oc8051_idata_n1688,
         oc8051_ram_top1_oc8051_idata_n1687,
         oc8051_ram_top1_oc8051_idata_n1686,
         oc8051_ram_top1_oc8051_idata_n1685,
         oc8051_ram_top1_oc8051_idata_n1684,
         oc8051_ram_top1_oc8051_idata_n1683,
         oc8051_ram_top1_oc8051_idata_n1682,
         oc8051_ram_top1_oc8051_idata_n1681,
         oc8051_ram_top1_oc8051_idata_n1680,
         oc8051_ram_top1_oc8051_idata_n1679,
         oc8051_ram_top1_oc8051_idata_n1678,
         oc8051_ram_top1_oc8051_idata_n1677,
         oc8051_ram_top1_oc8051_idata_n1676,
         oc8051_ram_top1_oc8051_idata_n1675,
         oc8051_ram_top1_oc8051_idata_n1674,
         oc8051_ram_top1_oc8051_idata_n1673,
         oc8051_ram_top1_oc8051_idata_n1672,
         oc8051_ram_top1_oc8051_idata_n1671,
         oc8051_ram_top1_oc8051_idata_n1670,
         oc8051_ram_top1_oc8051_idata_n1669,
         oc8051_ram_top1_oc8051_idata_n1668,
         oc8051_ram_top1_oc8051_idata_n1667,
         oc8051_ram_top1_oc8051_idata_n1666,
         oc8051_ram_top1_oc8051_idata_n1665,
         oc8051_ram_top1_oc8051_idata_n1664,
         oc8051_ram_top1_oc8051_idata_n1663,
         oc8051_ram_top1_oc8051_idata_n1662,
         oc8051_ram_top1_oc8051_idata_n1661,
         oc8051_ram_top1_oc8051_idata_n1660,
         oc8051_ram_top1_oc8051_idata_n1659,
         oc8051_ram_top1_oc8051_idata_n1658,
         oc8051_ram_top1_oc8051_idata_n1657,
         oc8051_ram_top1_oc8051_idata_n1656,
         oc8051_ram_top1_oc8051_idata_n1655,
         oc8051_ram_top1_oc8051_idata_n1654,
         oc8051_ram_top1_oc8051_idata_n1653,
         oc8051_ram_top1_oc8051_idata_n1652,
         oc8051_ram_top1_oc8051_idata_n1651,
         oc8051_ram_top1_oc8051_idata_n1650,
         oc8051_ram_top1_oc8051_idata_n1649,
         oc8051_ram_top1_oc8051_idata_n1648,
         oc8051_ram_top1_oc8051_idata_n1647,
         oc8051_ram_top1_oc8051_idata_n1646,
         oc8051_ram_top1_oc8051_idata_n1645,
         oc8051_ram_top1_oc8051_idata_n1644,
         oc8051_ram_top1_oc8051_idata_n1643,
         oc8051_ram_top1_oc8051_idata_n1642,
         oc8051_ram_top1_oc8051_idata_n1641,
         oc8051_ram_top1_oc8051_idata_n1640,
         oc8051_ram_top1_oc8051_idata_n1639,
         oc8051_ram_top1_oc8051_idata_n1638,
         oc8051_ram_top1_oc8051_idata_n1637,
         oc8051_ram_top1_oc8051_idata_n1636,
         oc8051_ram_top1_oc8051_idata_n1635,
         oc8051_ram_top1_oc8051_idata_n1634,
         oc8051_ram_top1_oc8051_idata_n1633,
         oc8051_ram_top1_oc8051_idata_n1632,
         oc8051_ram_top1_oc8051_idata_n1631,
         oc8051_ram_top1_oc8051_idata_n1630,
         oc8051_ram_top1_oc8051_idata_n1629,
         oc8051_ram_top1_oc8051_idata_n1628,
         oc8051_ram_top1_oc8051_idata_n1627,
         oc8051_ram_top1_oc8051_idata_n1626,
         oc8051_ram_top1_oc8051_idata_n1625,
         oc8051_ram_top1_oc8051_idata_n1624,
         oc8051_ram_top1_oc8051_idata_n1623,
         oc8051_ram_top1_oc8051_idata_n1622,
         oc8051_ram_top1_oc8051_idata_n1621,
         oc8051_ram_top1_oc8051_idata_n1620,
         oc8051_ram_top1_oc8051_idata_n1619,
         oc8051_ram_top1_oc8051_idata_n1618,
         oc8051_ram_top1_oc8051_idata_n1617,
         oc8051_ram_top1_oc8051_idata_n1616,
         oc8051_ram_top1_oc8051_idata_n1615,
         oc8051_ram_top1_oc8051_idata_n1614,
         oc8051_ram_top1_oc8051_idata_n1613,
         oc8051_ram_top1_oc8051_idata_n1612,
         oc8051_ram_top1_oc8051_idata_n1611,
         oc8051_ram_top1_oc8051_idata_n1610,
         oc8051_ram_top1_oc8051_idata_n1609,
         oc8051_ram_top1_oc8051_idata_n1608,
         oc8051_ram_top1_oc8051_idata_n1607,
         oc8051_ram_top1_oc8051_idata_n1606,
         oc8051_ram_top1_oc8051_idata_n1605,
         oc8051_ram_top1_oc8051_idata_n1604,
         oc8051_ram_top1_oc8051_idata_n1603,
         oc8051_ram_top1_oc8051_idata_n1602,
         oc8051_ram_top1_oc8051_idata_n1601,
         oc8051_ram_top1_oc8051_idata_n1600,
         oc8051_ram_top1_oc8051_idata_n1599,
         oc8051_ram_top1_oc8051_idata_n1598,
         oc8051_ram_top1_oc8051_idata_n1597,
         oc8051_ram_top1_oc8051_idata_n1596,
         oc8051_ram_top1_oc8051_idata_n1595,
         oc8051_ram_top1_oc8051_idata_n1594,
         oc8051_ram_top1_oc8051_idata_n1593,
         oc8051_ram_top1_oc8051_idata_n1592,
         oc8051_ram_top1_oc8051_idata_n1591,
         oc8051_ram_top1_oc8051_idata_n1590,
         oc8051_ram_top1_oc8051_idata_n1589,
         oc8051_ram_top1_oc8051_idata_n1588,
         oc8051_ram_top1_oc8051_idata_n1587,
         oc8051_ram_top1_oc8051_idata_n1586,
         oc8051_ram_top1_oc8051_idata_n1585,
         oc8051_ram_top1_oc8051_idata_n1584,
         oc8051_ram_top1_oc8051_idata_n1583,
         oc8051_ram_top1_oc8051_idata_n1582,
         oc8051_ram_top1_oc8051_idata_n1581,
         oc8051_ram_top1_oc8051_idata_n1580,
         oc8051_ram_top1_oc8051_idata_n1579,
         oc8051_ram_top1_oc8051_idata_n1578,
         oc8051_ram_top1_oc8051_idata_n1577,
         oc8051_ram_top1_oc8051_idata_n1576,
         oc8051_ram_top1_oc8051_idata_n1575,
         oc8051_ram_top1_oc8051_idata_n1574,
         oc8051_ram_top1_oc8051_idata_n1573,
         oc8051_ram_top1_oc8051_idata_n1572,
         oc8051_ram_top1_oc8051_idata_n1571,
         oc8051_ram_top1_oc8051_idata_n1570,
         oc8051_ram_top1_oc8051_idata_n1569,
         oc8051_ram_top1_oc8051_idata_n1568,
         oc8051_ram_top1_oc8051_idata_n1567,
         oc8051_ram_top1_oc8051_idata_n1566,
         oc8051_ram_top1_oc8051_idata_n1565,
         oc8051_ram_top1_oc8051_idata_n1564,
         oc8051_ram_top1_oc8051_idata_n1563,
         oc8051_ram_top1_oc8051_idata_n1562,
         oc8051_ram_top1_oc8051_idata_n1561,
         oc8051_ram_top1_oc8051_idata_n1560,
         oc8051_ram_top1_oc8051_idata_n1559,
         oc8051_ram_top1_oc8051_idata_n1558,
         oc8051_ram_top1_oc8051_idata_n1557,
         oc8051_ram_top1_oc8051_idata_n1556,
         oc8051_ram_top1_oc8051_idata_n1555,
         oc8051_ram_top1_oc8051_idata_n1554,
         oc8051_ram_top1_oc8051_idata_n1553,
         oc8051_ram_top1_oc8051_idata_n1552,
         oc8051_ram_top1_oc8051_idata_n1551,
         oc8051_ram_top1_oc8051_idata_n1550,
         oc8051_ram_top1_oc8051_idata_n1549,
         oc8051_ram_top1_oc8051_idata_n1548,
         oc8051_ram_top1_oc8051_idata_n1547,
         oc8051_ram_top1_oc8051_idata_n1546,
         oc8051_ram_top1_oc8051_idata_n1545,
         oc8051_ram_top1_oc8051_idata_n1544,
         oc8051_ram_top1_oc8051_idata_n1543,
         oc8051_ram_top1_oc8051_idata_n1542,
         oc8051_ram_top1_oc8051_idata_n1541,
         oc8051_ram_top1_oc8051_idata_n1540,
         oc8051_ram_top1_oc8051_idata_n1539,
         oc8051_ram_top1_oc8051_idata_n1538,
         oc8051_ram_top1_oc8051_idata_n1537,
         oc8051_ram_top1_oc8051_idata_n1536,
         oc8051_ram_top1_oc8051_idata_n1535,
         oc8051_ram_top1_oc8051_idata_n1534,
         oc8051_ram_top1_oc8051_idata_n1533,
         oc8051_ram_top1_oc8051_idata_n1532,
         oc8051_ram_top1_oc8051_idata_n1531,
         oc8051_ram_top1_oc8051_idata_n1530,
         oc8051_ram_top1_oc8051_idata_n1529,
         oc8051_ram_top1_oc8051_idata_n1528,
         oc8051_ram_top1_oc8051_idata_n1527,
         oc8051_ram_top1_oc8051_idata_n1526,
         oc8051_ram_top1_oc8051_idata_n1525,
         oc8051_ram_top1_oc8051_idata_n1524,
         oc8051_ram_top1_oc8051_idata_n1523,
         oc8051_ram_top1_oc8051_idata_n1522,
         oc8051_ram_top1_oc8051_idata_n1521,
         oc8051_ram_top1_oc8051_idata_n1520,
         oc8051_ram_top1_oc8051_idata_n1519,
         oc8051_ram_top1_oc8051_idata_n1518,
         oc8051_ram_top1_oc8051_idata_n1517,
         oc8051_ram_top1_oc8051_idata_n1516,
         oc8051_ram_top1_oc8051_idata_n1515,
         oc8051_ram_top1_oc8051_idata_n1514,
         oc8051_ram_top1_oc8051_idata_n1513,
         oc8051_ram_top1_oc8051_idata_n1512,
         oc8051_ram_top1_oc8051_idata_n1511,
         oc8051_ram_top1_oc8051_idata_n1510,
         oc8051_ram_top1_oc8051_idata_n1509,
         oc8051_ram_top1_oc8051_idata_n1508,
         oc8051_ram_top1_oc8051_idata_n1507,
         oc8051_ram_top1_oc8051_idata_n1506,
         oc8051_ram_top1_oc8051_idata_n1505,
         oc8051_ram_top1_oc8051_idata_n1504,
         oc8051_ram_top1_oc8051_idata_n1503,
         oc8051_ram_top1_oc8051_idata_n1502,
         oc8051_ram_top1_oc8051_idata_n1501,
         oc8051_ram_top1_oc8051_idata_n1500,
         oc8051_ram_top1_oc8051_idata_n1499,
         oc8051_ram_top1_oc8051_idata_n1498,
         oc8051_ram_top1_oc8051_idata_n1497,
         oc8051_ram_top1_oc8051_idata_n1496,
         oc8051_ram_top1_oc8051_idata_n1495,
         oc8051_ram_top1_oc8051_idata_n1494,
         oc8051_ram_top1_oc8051_idata_n1493,
         oc8051_ram_top1_oc8051_idata_n1492,
         oc8051_ram_top1_oc8051_idata_n1491,
         oc8051_ram_top1_oc8051_idata_n1490,
         oc8051_ram_top1_oc8051_idata_n1489,
         oc8051_ram_top1_oc8051_idata_n1488,
         oc8051_ram_top1_oc8051_idata_n1487,
         oc8051_ram_top1_oc8051_idata_n1486,
         oc8051_ram_top1_oc8051_idata_n1485,
         oc8051_ram_top1_oc8051_idata_n1484,
         oc8051_ram_top1_oc8051_idata_n1483,
         oc8051_ram_top1_oc8051_idata_n1482,
         oc8051_ram_top1_oc8051_idata_n1481,
         oc8051_ram_top1_oc8051_idata_n1480,
         oc8051_ram_top1_oc8051_idata_n1479,
         oc8051_ram_top1_oc8051_idata_n1478,
         oc8051_ram_top1_oc8051_idata_n1477,
         oc8051_ram_top1_oc8051_idata_n1476,
         oc8051_ram_top1_oc8051_idata_n1475,
         oc8051_ram_top1_oc8051_idata_n1474,
         oc8051_ram_top1_oc8051_idata_n1473,
         oc8051_ram_top1_oc8051_idata_n1472,
         oc8051_ram_top1_oc8051_idata_n1471,
         oc8051_ram_top1_oc8051_idata_n1470,
         oc8051_ram_top1_oc8051_idata_n1469,
         oc8051_ram_top1_oc8051_idata_n1468,
         oc8051_ram_top1_oc8051_idata_n1467,
         oc8051_ram_top1_oc8051_idata_n1466,
         oc8051_ram_top1_oc8051_idata_n1465,
         oc8051_ram_top1_oc8051_idata_n1464,
         oc8051_ram_top1_oc8051_idata_n1463,
         oc8051_ram_top1_oc8051_idata_n1462,
         oc8051_ram_top1_oc8051_idata_n1461,
         oc8051_ram_top1_oc8051_idata_n1460,
         oc8051_ram_top1_oc8051_idata_n1459,
         oc8051_ram_top1_oc8051_idata_n1458,
         oc8051_ram_top1_oc8051_idata_n1457,
         oc8051_ram_top1_oc8051_idata_n1456,
         oc8051_ram_top1_oc8051_idata_n1455,
         oc8051_ram_top1_oc8051_idata_n1454,
         oc8051_ram_top1_oc8051_idata_n1453,
         oc8051_ram_top1_oc8051_idata_n1452,
         oc8051_ram_top1_oc8051_idata_n1451,
         oc8051_ram_top1_oc8051_idata_n1450,
         oc8051_ram_top1_oc8051_idata_n1449,
         oc8051_ram_top1_oc8051_idata_n1448,
         oc8051_ram_top1_oc8051_idata_n1447,
         oc8051_ram_top1_oc8051_idata_n1446,
         oc8051_ram_top1_oc8051_idata_n1445,
         oc8051_ram_top1_oc8051_idata_n1444,
         oc8051_ram_top1_oc8051_idata_n1443,
         oc8051_ram_top1_oc8051_idata_n1442,
         oc8051_ram_top1_oc8051_idata_n1441,
         oc8051_ram_top1_oc8051_idata_n1440,
         oc8051_ram_top1_oc8051_idata_n1439,
         oc8051_ram_top1_oc8051_idata_n1438,
         oc8051_ram_top1_oc8051_idata_n1437,
         oc8051_ram_top1_oc8051_idata_n1436,
         oc8051_ram_top1_oc8051_idata_n1435,
         oc8051_ram_top1_oc8051_idata_n1434,
         oc8051_ram_top1_oc8051_idata_n1433,
         oc8051_ram_top1_oc8051_idata_n1432,
         oc8051_ram_top1_oc8051_idata_n1431,
         oc8051_ram_top1_oc8051_idata_n1430,
         oc8051_ram_top1_oc8051_idata_n1429,
         oc8051_ram_top1_oc8051_idata_n1428,
         oc8051_ram_top1_oc8051_idata_n1427,
         oc8051_ram_top1_oc8051_idata_n1426,
         oc8051_ram_top1_oc8051_idata_n1425,
         oc8051_ram_top1_oc8051_idata_n1424,
         oc8051_ram_top1_oc8051_idata_n1423,
         oc8051_ram_top1_oc8051_idata_n1422,
         oc8051_ram_top1_oc8051_idata_n1421,
         oc8051_ram_top1_oc8051_idata_n1420,
         oc8051_ram_top1_oc8051_idata_n1419,
         oc8051_ram_top1_oc8051_idata_n1418,
         oc8051_ram_top1_oc8051_idata_n1417,
         oc8051_ram_top1_oc8051_idata_n1416,
         oc8051_ram_top1_oc8051_idata_n1415,
         oc8051_ram_top1_oc8051_idata_n1414,
         oc8051_ram_top1_oc8051_idata_n1413,
         oc8051_ram_top1_oc8051_idata_n1412,
         oc8051_ram_top1_oc8051_idata_n1411,
         oc8051_ram_top1_oc8051_idata_n1410,
         oc8051_ram_top1_oc8051_idata_n1409,
         oc8051_ram_top1_oc8051_idata_n1408,
         oc8051_ram_top1_oc8051_idata_n1407,
         oc8051_ram_top1_oc8051_idata_n1406,
         oc8051_ram_top1_oc8051_idata_n1405,
         oc8051_ram_top1_oc8051_idata_n1404,
         oc8051_ram_top1_oc8051_idata_n1403,
         oc8051_ram_top1_oc8051_idata_n1402,
         oc8051_ram_top1_oc8051_idata_n1401,
         oc8051_ram_top1_oc8051_idata_n1400,
         oc8051_ram_top1_oc8051_idata_n1399,
         oc8051_ram_top1_oc8051_idata_n1398,
         oc8051_ram_top1_oc8051_idata_n1397,
         oc8051_ram_top1_oc8051_idata_n1396,
         oc8051_ram_top1_oc8051_idata_n1395,
         oc8051_ram_top1_oc8051_idata_n1394,
         oc8051_ram_top1_oc8051_idata_n1393,
         oc8051_ram_top1_oc8051_idata_n1392,
         oc8051_ram_top1_oc8051_idata_n1391,
         oc8051_ram_top1_oc8051_idata_n1390,
         oc8051_ram_top1_oc8051_idata_n1389,
         oc8051_ram_top1_oc8051_idata_n1388,
         oc8051_ram_top1_oc8051_idata_n1387,
         oc8051_ram_top1_oc8051_idata_n1386,
         oc8051_ram_top1_oc8051_idata_n1385,
         oc8051_ram_top1_oc8051_idata_n1384,
         oc8051_ram_top1_oc8051_idata_n1383,
         oc8051_ram_top1_oc8051_idata_n1382,
         oc8051_ram_top1_oc8051_idata_n1381,
         oc8051_ram_top1_oc8051_idata_n1380,
         oc8051_ram_top1_oc8051_idata_n1379,
         oc8051_ram_top1_oc8051_idata_n1378,
         oc8051_ram_top1_oc8051_idata_n1377,
         oc8051_ram_top1_oc8051_idata_n1376,
         oc8051_ram_top1_oc8051_idata_n1375,
         oc8051_ram_top1_oc8051_idata_n1374,
         oc8051_ram_top1_oc8051_idata_n1373,
         oc8051_ram_top1_oc8051_idata_n1372,
         oc8051_ram_top1_oc8051_idata_n1371,
         oc8051_ram_top1_oc8051_idata_n1370,
         oc8051_ram_top1_oc8051_idata_n1369,
         oc8051_ram_top1_oc8051_idata_n1368,
         oc8051_ram_top1_oc8051_idata_n1367,
         oc8051_ram_top1_oc8051_idata_n1366,
         oc8051_ram_top1_oc8051_idata_n1365,
         oc8051_ram_top1_oc8051_idata_n1364,
         oc8051_ram_top1_oc8051_idata_n1363,
         oc8051_ram_top1_oc8051_idata_n1362,
         oc8051_ram_top1_oc8051_idata_n1361,
         oc8051_ram_top1_oc8051_idata_n1360,
         oc8051_ram_top1_oc8051_idata_n1359,
         oc8051_ram_top1_oc8051_idata_n1358,
         oc8051_ram_top1_oc8051_idata_n1357,
         oc8051_ram_top1_oc8051_idata_n1356,
         oc8051_ram_top1_oc8051_idata_n1355,
         oc8051_ram_top1_oc8051_idata_n1354,
         oc8051_ram_top1_oc8051_idata_n1353,
         oc8051_ram_top1_oc8051_idata_n1352,
         oc8051_ram_top1_oc8051_idata_n1351,
         oc8051_ram_top1_oc8051_idata_n1350,
         oc8051_ram_top1_oc8051_idata_n1349,
         oc8051_ram_top1_oc8051_idata_n1348,
         oc8051_ram_top1_oc8051_idata_n1347,
         oc8051_ram_top1_oc8051_idata_n1346,
         oc8051_ram_top1_oc8051_idata_n1345,
         oc8051_ram_top1_oc8051_idata_n1344,
         oc8051_ram_top1_oc8051_idata_n1343,
         oc8051_ram_top1_oc8051_idata_n1342,
         oc8051_ram_top1_oc8051_idata_n1341,
         oc8051_ram_top1_oc8051_idata_n1340,
         oc8051_ram_top1_oc8051_idata_n1339,
         oc8051_ram_top1_oc8051_idata_n1338,
         oc8051_ram_top1_oc8051_idata_n1337,
         oc8051_ram_top1_oc8051_idata_n1336,
         oc8051_ram_top1_oc8051_idata_n1335,
         oc8051_ram_top1_oc8051_idata_n1334,
         oc8051_ram_top1_oc8051_idata_n1333,
         oc8051_ram_top1_oc8051_idata_n1332,
         oc8051_ram_top1_oc8051_idata_n1331,
         oc8051_ram_top1_oc8051_idata_n1330,
         oc8051_ram_top1_oc8051_idata_n1329,
         oc8051_ram_top1_oc8051_idata_n1328,
         oc8051_ram_top1_oc8051_idata_n1327,
         oc8051_ram_top1_oc8051_idata_n1326,
         oc8051_ram_top1_oc8051_idata_n1325,
         oc8051_ram_top1_oc8051_idata_n1324,
         oc8051_ram_top1_oc8051_idata_n1323,
         oc8051_ram_top1_oc8051_idata_n1322,
         oc8051_ram_top1_oc8051_idata_n1321,
         oc8051_ram_top1_oc8051_idata_n1320,
         oc8051_ram_top1_oc8051_idata_n1319,
         oc8051_ram_top1_oc8051_idata_n1318,
         oc8051_ram_top1_oc8051_idata_n1317,
         oc8051_ram_top1_oc8051_idata_n1316,
         oc8051_ram_top1_oc8051_idata_n1315,
         oc8051_ram_top1_oc8051_idata_n1314,
         oc8051_ram_top1_oc8051_idata_n1313,
         oc8051_ram_top1_oc8051_idata_n1312,
         oc8051_ram_top1_oc8051_idata_n1311,
         oc8051_ram_top1_oc8051_idata_n1310,
         oc8051_ram_top1_oc8051_idata_n1309,
         oc8051_ram_top1_oc8051_idata_n1308,
         oc8051_ram_top1_oc8051_idata_n1307,
         oc8051_ram_top1_oc8051_idata_n1306,
         oc8051_ram_top1_oc8051_idata_n1305,
         oc8051_ram_top1_oc8051_idata_n1304,
         oc8051_ram_top1_oc8051_idata_n1303,
         oc8051_ram_top1_oc8051_idata_n1302,
         oc8051_ram_top1_oc8051_idata_n1301,
         oc8051_ram_top1_oc8051_idata_n1300,
         oc8051_ram_top1_oc8051_idata_n1299,
         oc8051_ram_top1_oc8051_idata_n1298,
         oc8051_ram_top1_oc8051_idata_n1297,
         oc8051_ram_top1_oc8051_idata_n1296,
         oc8051_ram_top1_oc8051_idata_n1295,
         oc8051_ram_top1_oc8051_idata_n1294,
         oc8051_ram_top1_oc8051_idata_n1293,
         oc8051_ram_top1_oc8051_idata_n1292,
         oc8051_ram_top1_oc8051_idata_n1291,
         oc8051_ram_top1_oc8051_idata_n1290,
         oc8051_ram_top1_oc8051_idata_n1289,
         oc8051_ram_top1_oc8051_idata_n1288,
         oc8051_ram_top1_oc8051_idata_n1287,
         oc8051_ram_top1_oc8051_idata_n1286,
         oc8051_ram_top1_oc8051_idata_n1285,
         oc8051_ram_top1_oc8051_idata_n1284,
         oc8051_ram_top1_oc8051_idata_n1283,
         oc8051_ram_top1_oc8051_idata_n1282,
         oc8051_ram_top1_oc8051_idata_n1281,
         oc8051_ram_top1_oc8051_idata_n1280,
         oc8051_ram_top1_oc8051_idata_n1279,
         oc8051_ram_top1_oc8051_idata_n1278,
         oc8051_ram_top1_oc8051_idata_n1277,
         oc8051_ram_top1_oc8051_idata_n1276,
         oc8051_ram_top1_oc8051_idata_n1275,
         oc8051_ram_top1_oc8051_idata_n1274,
         oc8051_ram_top1_oc8051_idata_n1273,
         oc8051_ram_top1_oc8051_idata_n1272,
         oc8051_ram_top1_oc8051_idata_n1271,
         oc8051_ram_top1_oc8051_idata_n1270,
         oc8051_ram_top1_oc8051_idata_n1269,
         oc8051_ram_top1_oc8051_idata_n1268,
         oc8051_ram_top1_oc8051_idata_n1267,
         oc8051_ram_top1_oc8051_idata_n1266,
         oc8051_ram_top1_oc8051_idata_n1265,
         oc8051_ram_top1_oc8051_idata_n1264,
         oc8051_ram_top1_oc8051_idata_n1263,
         oc8051_ram_top1_oc8051_idata_n1262,
         oc8051_ram_top1_oc8051_idata_n1261,
         oc8051_ram_top1_oc8051_idata_n1260,
         oc8051_ram_top1_oc8051_idata_n1259,
         oc8051_ram_top1_oc8051_idata_n1258,
         oc8051_ram_top1_oc8051_idata_n1257,
         oc8051_ram_top1_oc8051_idata_n1256,
         oc8051_ram_top1_oc8051_idata_n1255,
         oc8051_ram_top1_oc8051_idata_n1254,
         oc8051_ram_top1_oc8051_idata_n1253,
         oc8051_ram_top1_oc8051_idata_n1252,
         oc8051_ram_top1_oc8051_idata_n1251,
         oc8051_ram_top1_oc8051_idata_n1250,
         oc8051_ram_top1_oc8051_idata_n1249,
         oc8051_ram_top1_oc8051_idata_n1248,
         oc8051_ram_top1_oc8051_idata_n1247,
         oc8051_ram_top1_oc8051_idata_n1246,
         oc8051_ram_top1_oc8051_idata_n1245,
         oc8051_ram_top1_oc8051_idata_n1244,
         oc8051_ram_top1_oc8051_idata_n1243,
         oc8051_ram_top1_oc8051_idata_n1242,
         oc8051_ram_top1_oc8051_idata_n1241,
         oc8051_ram_top1_oc8051_idata_n1240,
         oc8051_ram_top1_oc8051_idata_n1239,
         oc8051_ram_top1_oc8051_idata_n1238,
         oc8051_ram_top1_oc8051_idata_n1237,
         oc8051_ram_top1_oc8051_idata_n1236,
         oc8051_ram_top1_oc8051_idata_n1235,
         oc8051_ram_top1_oc8051_idata_n1234,
         oc8051_ram_top1_oc8051_idata_n1233,
         oc8051_ram_top1_oc8051_idata_n1232,
         oc8051_ram_top1_oc8051_idata_n1231,
         oc8051_ram_top1_oc8051_idata_n1230,
         oc8051_ram_top1_oc8051_idata_n1229,
         oc8051_ram_top1_oc8051_idata_n1228,
         oc8051_ram_top1_oc8051_idata_n1227,
         oc8051_ram_top1_oc8051_idata_n1226,
         oc8051_ram_top1_oc8051_idata_n1225,
         oc8051_ram_top1_oc8051_idata_n1224,
         oc8051_ram_top1_oc8051_idata_n1223,
         oc8051_ram_top1_oc8051_idata_n1222,
         oc8051_ram_top1_oc8051_idata_n1221,
         oc8051_ram_top1_oc8051_idata_n1220,
         oc8051_ram_top1_oc8051_idata_n1219,
         oc8051_ram_top1_oc8051_idata_n1218,
         oc8051_ram_top1_oc8051_idata_n1217,
         oc8051_ram_top1_oc8051_idata_n1216,
         oc8051_ram_top1_oc8051_idata_n1215,
         oc8051_ram_top1_oc8051_idata_n1214,
         oc8051_ram_top1_oc8051_idata_n1213,
         oc8051_ram_top1_oc8051_idata_n1212,
         oc8051_ram_top1_oc8051_idata_n1211,
         oc8051_ram_top1_oc8051_idata_n1210,
         oc8051_ram_top1_oc8051_idata_n1209,
         oc8051_ram_top1_oc8051_idata_n1208,
         oc8051_ram_top1_oc8051_idata_n1207,
         oc8051_ram_top1_oc8051_idata_n1206,
         oc8051_ram_top1_oc8051_idata_n1205,
         oc8051_ram_top1_oc8051_idata_n1204,
         oc8051_ram_top1_oc8051_idata_n1203,
         oc8051_ram_top1_oc8051_idata_n1202,
         oc8051_ram_top1_oc8051_idata_n1201,
         oc8051_ram_top1_oc8051_idata_n1200,
         oc8051_ram_top1_oc8051_idata_n1199,
         oc8051_ram_top1_oc8051_idata_n1198,
         oc8051_ram_top1_oc8051_idata_n1197,
         oc8051_ram_top1_oc8051_idata_n1196,
         oc8051_ram_top1_oc8051_idata_n1195,
         oc8051_ram_top1_oc8051_idata_n1194,
         oc8051_ram_top1_oc8051_idata_n1193,
         oc8051_ram_top1_oc8051_idata_n1192,
         oc8051_ram_top1_oc8051_idata_n1191,
         oc8051_ram_top1_oc8051_idata_n1190,
         oc8051_ram_top1_oc8051_idata_n1189,
         oc8051_ram_top1_oc8051_idata_n1188,
         oc8051_ram_top1_oc8051_idata_n1187,
         oc8051_ram_top1_oc8051_idata_n1186,
         oc8051_ram_top1_oc8051_idata_n1185,
         oc8051_ram_top1_oc8051_idata_n1184,
         oc8051_ram_top1_oc8051_idata_n1183,
         oc8051_ram_top1_oc8051_idata_n1182,
         oc8051_ram_top1_oc8051_idata_n1181,
         oc8051_ram_top1_oc8051_idata_n1180,
         oc8051_ram_top1_oc8051_idata_n1179,
         oc8051_ram_top1_oc8051_idata_n1178,
         oc8051_ram_top1_oc8051_idata_n1177,
         oc8051_ram_top1_oc8051_idata_n1176,
         oc8051_ram_top1_oc8051_idata_n1175,
         oc8051_ram_top1_oc8051_idata_n1174,
         oc8051_ram_top1_oc8051_idata_n1173,
         oc8051_ram_top1_oc8051_idata_n1172,
         oc8051_ram_top1_oc8051_idata_n1171,
         oc8051_ram_top1_oc8051_idata_n1170,
         oc8051_ram_top1_oc8051_idata_n1169,
         oc8051_ram_top1_oc8051_idata_n1168,
         oc8051_ram_top1_oc8051_idata_n1167,
         oc8051_ram_top1_oc8051_idata_n1166,
         oc8051_ram_top1_oc8051_idata_n1165,
         oc8051_ram_top1_oc8051_idata_n1164,
         oc8051_ram_top1_oc8051_idata_n1163,
         oc8051_ram_top1_oc8051_idata_n1162,
         oc8051_ram_top1_oc8051_idata_n1161,
         oc8051_ram_top1_oc8051_idata_n1160,
         oc8051_ram_top1_oc8051_idata_n1159,
         oc8051_ram_top1_oc8051_idata_n1158,
         oc8051_ram_top1_oc8051_idata_n1157,
         oc8051_ram_top1_oc8051_idata_n1156,
         oc8051_ram_top1_oc8051_idata_n1155,
         oc8051_ram_top1_oc8051_idata_n1154,
         oc8051_ram_top1_oc8051_idata_n1153,
         oc8051_ram_top1_oc8051_idata_n1152,
         oc8051_ram_top1_oc8051_idata_n1151,
         oc8051_ram_top1_oc8051_idata_n1150,
         oc8051_ram_top1_oc8051_idata_n1149,
         oc8051_ram_top1_oc8051_idata_n1148,
         oc8051_ram_top1_oc8051_idata_n1147,
         oc8051_ram_top1_oc8051_idata_n1146,
         oc8051_ram_top1_oc8051_idata_n1145,
         oc8051_ram_top1_oc8051_idata_n1144,
         oc8051_ram_top1_oc8051_idata_n1143,
         oc8051_ram_top1_oc8051_idata_n1142,
         oc8051_ram_top1_oc8051_idata_n1141,
         oc8051_ram_top1_oc8051_idata_n1140,
         oc8051_ram_top1_oc8051_idata_n1139,
         oc8051_ram_top1_oc8051_idata_n1138,
         oc8051_ram_top1_oc8051_idata_n1137,
         oc8051_ram_top1_oc8051_idata_n1136,
         oc8051_ram_top1_oc8051_idata_n1135,
         oc8051_ram_top1_oc8051_idata_n1134,
         oc8051_ram_top1_oc8051_idata_n1133,
         oc8051_ram_top1_oc8051_idata_n1132,
         oc8051_ram_top1_oc8051_idata_n1131,
         oc8051_ram_top1_oc8051_idata_n1130,
         oc8051_ram_top1_oc8051_idata_n1129,
         oc8051_ram_top1_oc8051_idata_n1128,
         oc8051_ram_top1_oc8051_idata_n1127,
         oc8051_ram_top1_oc8051_idata_n1126,
         oc8051_ram_top1_oc8051_idata_n1125,
         oc8051_ram_top1_oc8051_idata_n1124,
         oc8051_ram_top1_oc8051_idata_n1123,
         oc8051_ram_top1_oc8051_idata_n1122,
         oc8051_ram_top1_oc8051_idata_n1121,
         oc8051_ram_top1_oc8051_idata_n1120,
         oc8051_ram_top1_oc8051_idata_n1119,
         oc8051_ram_top1_oc8051_idata_n1118,
         oc8051_ram_top1_oc8051_idata_n1117,
         oc8051_ram_top1_oc8051_idata_n1116,
         oc8051_ram_top1_oc8051_idata_n1115,
         oc8051_ram_top1_oc8051_idata_n1114,
         oc8051_ram_top1_oc8051_idata_n1113,
         oc8051_ram_top1_oc8051_idata_n1112,
         oc8051_ram_top1_oc8051_idata_n1111,
         oc8051_ram_top1_oc8051_idata_n1110,
         oc8051_ram_top1_oc8051_idata_n1109,
         oc8051_ram_top1_oc8051_idata_n1108,
         oc8051_ram_top1_oc8051_idata_n1107,
         oc8051_ram_top1_oc8051_idata_n1106,
         oc8051_ram_top1_oc8051_idata_n1105,
         oc8051_ram_top1_oc8051_idata_n1104,
         oc8051_ram_top1_oc8051_idata_n1103,
         oc8051_ram_top1_oc8051_idata_n1102,
         oc8051_ram_top1_oc8051_idata_n1101,
         oc8051_ram_top1_oc8051_idata_n1100,
         oc8051_ram_top1_oc8051_idata_n1099,
         oc8051_ram_top1_oc8051_idata_n1098,
         oc8051_ram_top1_oc8051_idata_n1097,
         oc8051_ram_top1_oc8051_idata_n1096,
         oc8051_ram_top1_oc8051_idata_n1095,
         oc8051_ram_top1_oc8051_idata_n1094,
         oc8051_ram_top1_oc8051_idata_n1093,
         oc8051_ram_top1_oc8051_idata_n1092,
         oc8051_ram_top1_oc8051_idata_n1091,
         oc8051_ram_top1_oc8051_idata_n1090,
         oc8051_ram_top1_oc8051_idata_n1089,
         oc8051_ram_top1_oc8051_idata_n1088,
         oc8051_ram_top1_oc8051_idata_n1087,
         oc8051_ram_top1_oc8051_idata_n1086,
         oc8051_ram_top1_oc8051_idata_n1085,
         oc8051_ram_top1_oc8051_idata_n1084,
         oc8051_ram_top1_oc8051_idata_n1083,
         oc8051_ram_top1_oc8051_idata_n1082,
         oc8051_ram_top1_oc8051_idata_n1081,
         oc8051_ram_top1_oc8051_idata_n1080,
         oc8051_ram_top1_oc8051_idata_n1079,
         oc8051_ram_top1_oc8051_idata_n1078,
         oc8051_ram_top1_oc8051_idata_n1077,
         oc8051_ram_top1_oc8051_idata_n1076,
         oc8051_ram_top1_oc8051_idata_n1075,
         oc8051_ram_top1_oc8051_idata_n1074,
         oc8051_ram_top1_oc8051_idata_n1073,
         oc8051_ram_top1_oc8051_idata_n1072,
         oc8051_ram_top1_oc8051_idata_n1071,
         oc8051_ram_top1_oc8051_idata_n1070,
         oc8051_ram_top1_oc8051_idata_n1069,
         oc8051_ram_top1_oc8051_idata_n1068,
         oc8051_ram_top1_oc8051_idata_n1067,
         oc8051_ram_top1_oc8051_idata_n1066,
         oc8051_ram_top1_oc8051_idata_n1065,
         oc8051_ram_top1_oc8051_idata_n1064,
         oc8051_ram_top1_oc8051_idata_n1063,
         oc8051_ram_top1_oc8051_idata_n1062,
         oc8051_ram_top1_oc8051_idata_n1061,
         oc8051_ram_top1_oc8051_idata_n1060,
         oc8051_ram_top1_oc8051_idata_n1059,
         oc8051_ram_top1_oc8051_idata_n1058,
         oc8051_ram_top1_oc8051_idata_n1057,
         oc8051_ram_top1_oc8051_idata_n1056,
         oc8051_ram_top1_oc8051_idata_n1055,
         oc8051_ram_top1_oc8051_idata_n1054,
         oc8051_ram_top1_oc8051_idata_n1053,
         oc8051_ram_top1_oc8051_idata_n1052,
         oc8051_ram_top1_oc8051_idata_n1051,
         oc8051_ram_top1_oc8051_idata_n1050,
         oc8051_ram_top1_oc8051_idata_n1049,
         oc8051_ram_top1_oc8051_idata_n1048,
         oc8051_ram_top1_oc8051_idata_n1047,
         oc8051_ram_top1_oc8051_idata_n1046,
         oc8051_ram_top1_oc8051_idata_n1045,
         oc8051_ram_top1_oc8051_idata_n1044,
         oc8051_ram_top1_oc8051_idata_n1043,
         oc8051_ram_top1_oc8051_idata_n1042,
         oc8051_ram_top1_oc8051_idata_n1041,
         oc8051_ram_top1_oc8051_idata_n1040,
         oc8051_ram_top1_oc8051_idata_n1039,
         oc8051_ram_top1_oc8051_idata_n1038,
         oc8051_ram_top1_oc8051_idata_n1037,
         oc8051_ram_top1_oc8051_idata_n1036,
         oc8051_ram_top1_oc8051_idata_n1035,
         oc8051_ram_top1_oc8051_idata_n1034,
         oc8051_ram_top1_oc8051_idata_n1033,
         oc8051_ram_top1_oc8051_idata_n1032,
         oc8051_ram_top1_oc8051_idata_n1031,
         oc8051_ram_top1_oc8051_idata_n1030,
         oc8051_ram_top1_oc8051_idata_n1029,
         oc8051_ram_top1_oc8051_idata_n1028,
         oc8051_ram_top1_oc8051_idata_n1027,
         oc8051_ram_top1_oc8051_idata_n1026,
         oc8051_ram_top1_oc8051_idata_n1025,
         oc8051_ram_top1_oc8051_idata_n1024,
         oc8051_ram_top1_oc8051_idata_n1023,
         oc8051_ram_top1_oc8051_idata_n1022,
         oc8051_ram_top1_oc8051_idata_n1021,
         oc8051_ram_top1_oc8051_idata_n1020,
         oc8051_ram_top1_oc8051_idata_n1019,
         oc8051_ram_top1_oc8051_idata_n1018,
         oc8051_ram_top1_oc8051_idata_n1017,
         oc8051_ram_top1_oc8051_idata_n1016,
         oc8051_ram_top1_oc8051_idata_n1015,
         oc8051_ram_top1_oc8051_idata_n1014,
         oc8051_ram_top1_oc8051_idata_n1013,
         oc8051_ram_top1_oc8051_idata_n1012,
         oc8051_ram_top1_oc8051_idata_n1011,
         oc8051_ram_top1_oc8051_idata_n1010,
         oc8051_ram_top1_oc8051_idata_n1009,
         oc8051_ram_top1_oc8051_idata_n1008,
         oc8051_ram_top1_oc8051_idata_n1007,
         oc8051_ram_top1_oc8051_idata_n1006,
         oc8051_ram_top1_oc8051_idata_n1005,
         oc8051_ram_top1_oc8051_idata_n1004,
         oc8051_ram_top1_oc8051_idata_n1003,
         oc8051_ram_top1_oc8051_idata_n1002,
         oc8051_ram_top1_oc8051_idata_n1001,
         oc8051_ram_top1_oc8051_idata_n1000, oc8051_ram_top1_oc8051_idata_n999,
         oc8051_ram_top1_oc8051_idata_n998, oc8051_ram_top1_oc8051_idata_n997,
         oc8051_ram_top1_oc8051_idata_n996, oc8051_ram_top1_oc8051_idata_n995,
         oc8051_ram_top1_oc8051_idata_n994, oc8051_ram_top1_oc8051_idata_n993,
         oc8051_ram_top1_oc8051_idata_n992, oc8051_ram_top1_oc8051_idata_n991,
         oc8051_ram_top1_oc8051_idata_n990, oc8051_ram_top1_oc8051_idata_n989,
         oc8051_ram_top1_oc8051_idata_n988, oc8051_ram_top1_oc8051_idata_n987,
         oc8051_ram_top1_oc8051_idata_n986, oc8051_ram_top1_oc8051_idata_n985,
         oc8051_ram_top1_oc8051_idata_n984, oc8051_ram_top1_oc8051_idata_n983,
         oc8051_ram_top1_oc8051_idata_n982, oc8051_ram_top1_oc8051_idata_n981,
         oc8051_ram_top1_oc8051_idata_n980, oc8051_ram_top1_oc8051_idata_n979,
         oc8051_ram_top1_oc8051_idata_n978, oc8051_ram_top1_oc8051_idata_n977,
         oc8051_ram_top1_oc8051_idata_n976, oc8051_ram_top1_oc8051_idata_n975,
         oc8051_ram_top1_oc8051_idata_n974, oc8051_ram_top1_oc8051_idata_n973,
         oc8051_ram_top1_oc8051_idata_n972, oc8051_ram_top1_oc8051_idata_n971,
         oc8051_ram_top1_oc8051_idata_n970, oc8051_ram_top1_oc8051_idata_n969,
         oc8051_ram_top1_oc8051_idata_n968, oc8051_ram_top1_oc8051_idata_n967,
         oc8051_ram_top1_oc8051_idata_n966, oc8051_ram_top1_oc8051_idata_n965,
         oc8051_ram_top1_oc8051_idata_n964, oc8051_ram_top1_oc8051_idata_n963,
         oc8051_ram_top1_oc8051_idata_n962, oc8051_ram_top1_oc8051_idata_n961,
         oc8051_ram_top1_oc8051_idata_n960, oc8051_ram_top1_oc8051_idata_n959,
         oc8051_ram_top1_oc8051_idata_n958, oc8051_ram_top1_oc8051_idata_n957,
         oc8051_ram_top1_oc8051_idata_n956, oc8051_ram_top1_oc8051_idata_n955,
         oc8051_ram_top1_oc8051_idata_n954, oc8051_ram_top1_oc8051_idata_n953,
         oc8051_ram_top1_oc8051_idata_n952, oc8051_ram_top1_oc8051_idata_n951,
         oc8051_ram_top1_oc8051_idata_n950, oc8051_ram_top1_oc8051_idata_n949,
         oc8051_ram_top1_oc8051_idata_n948, oc8051_ram_top1_oc8051_idata_n947,
         oc8051_ram_top1_oc8051_idata_n946, oc8051_ram_top1_oc8051_idata_n945,
         oc8051_ram_top1_oc8051_idata_n944, oc8051_ram_top1_oc8051_idata_n943,
         oc8051_ram_top1_oc8051_idata_n942, oc8051_ram_top1_oc8051_idata_n941,
         oc8051_ram_top1_oc8051_idata_n940, oc8051_ram_top1_oc8051_idata_n939,
         oc8051_ram_top1_oc8051_idata_n938, oc8051_ram_top1_oc8051_idata_n937,
         oc8051_ram_top1_oc8051_idata_n936, oc8051_ram_top1_oc8051_idata_n935,
         oc8051_ram_top1_oc8051_idata_n934, oc8051_ram_top1_oc8051_idata_n933,
         oc8051_ram_top1_oc8051_idata_n932, oc8051_ram_top1_oc8051_idata_n931,
         oc8051_ram_top1_oc8051_idata_n930, oc8051_ram_top1_oc8051_idata_n929,
         oc8051_ram_top1_oc8051_idata_n928, oc8051_ram_top1_oc8051_idata_n927,
         oc8051_ram_top1_oc8051_idata_n926, oc8051_ram_top1_oc8051_idata_n925,
         oc8051_ram_top1_oc8051_idata_n924, oc8051_ram_top1_oc8051_idata_n923,
         oc8051_ram_top1_oc8051_idata_n922, oc8051_ram_top1_oc8051_idata_n921,
         oc8051_ram_top1_oc8051_idata_n920, oc8051_ram_top1_oc8051_idata_n919,
         oc8051_ram_top1_oc8051_idata_n918, oc8051_ram_top1_oc8051_idata_n917,
         oc8051_ram_top1_oc8051_idata_n916, oc8051_ram_top1_oc8051_idata_n915,
         oc8051_ram_top1_oc8051_idata_n914, oc8051_ram_top1_oc8051_idata_n913,
         oc8051_ram_top1_oc8051_idata_n912, oc8051_ram_top1_oc8051_idata_n911,
         oc8051_ram_top1_oc8051_idata_n910, oc8051_ram_top1_oc8051_idata_n909,
         oc8051_ram_top1_oc8051_idata_n908, oc8051_ram_top1_oc8051_idata_n907,
         oc8051_ram_top1_oc8051_idata_n906, oc8051_ram_top1_oc8051_idata_n905,
         oc8051_ram_top1_oc8051_idata_n904, oc8051_ram_top1_oc8051_idata_n903,
         oc8051_ram_top1_oc8051_idata_n902, oc8051_ram_top1_oc8051_idata_n901,
         oc8051_ram_top1_oc8051_idata_n900, oc8051_ram_top1_oc8051_idata_n899,
         oc8051_ram_top1_oc8051_idata_n898, oc8051_ram_top1_oc8051_idata_n897,
         oc8051_ram_top1_oc8051_idata_n896, oc8051_ram_top1_oc8051_idata_n895,
         oc8051_ram_top1_oc8051_idata_n894, oc8051_ram_top1_oc8051_idata_n893,
         oc8051_ram_top1_oc8051_idata_n892, oc8051_ram_top1_oc8051_idata_n891,
         oc8051_ram_top1_oc8051_idata_n890, oc8051_ram_top1_oc8051_idata_n889,
         oc8051_ram_top1_oc8051_idata_n888, oc8051_ram_top1_oc8051_idata_n887,
         oc8051_ram_top1_oc8051_idata_n886, oc8051_ram_top1_oc8051_idata_n885,
         oc8051_ram_top1_oc8051_idata_n884, oc8051_ram_top1_oc8051_idata_n883,
         oc8051_ram_top1_oc8051_idata_n882, oc8051_ram_top1_oc8051_idata_n881,
         oc8051_ram_top1_oc8051_idata_n880, oc8051_ram_top1_oc8051_idata_n879,
         oc8051_ram_top1_oc8051_idata_n878, oc8051_ram_top1_oc8051_idata_n877,
         oc8051_ram_top1_oc8051_idata_n876, oc8051_ram_top1_oc8051_idata_n875,
         oc8051_ram_top1_oc8051_idata_n874, oc8051_ram_top1_oc8051_idata_n873,
         oc8051_ram_top1_oc8051_idata_n872, oc8051_ram_top1_oc8051_idata_n871,
         oc8051_ram_top1_oc8051_idata_n870, oc8051_ram_top1_oc8051_idata_n869,
         oc8051_ram_top1_oc8051_idata_n868, oc8051_ram_top1_oc8051_idata_n867,
         oc8051_ram_top1_oc8051_idata_n866, oc8051_ram_top1_oc8051_idata_n865,
         oc8051_ram_top1_oc8051_idata_n864, oc8051_ram_top1_oc8051_idata_n863,
         oc8051_ram_top1_oc8051_idata_n862, oc8051_ram_top1_oc8051_idata_n861,
         oc8051_ram_top1_oc8051_idata_n860, oc8051_ram_top1_oc8051_idata_n859,
         oc8051_ram_top1_oc8051_idata_n858, oc8051_ram_top1_oc8051_idata_n857,
         oc8051_ram_top1_oc8051_idata_n856, oc8051_ram_top1_oc8051_idata_n855,
         oc8051_ram_top1_oc8051_idata_n854, oc8051_ram_top1_oc8051_idata_n853,
         oc8051_ram_top1_oc8051_idata_n852, oc8051_ram_top1_oc8051_idata_n851,
         oc8051_ram_top1_oc8051_idata_n850, oc8051_ram_top1_oc8051_idata_n849,
         oc8051_ram_top1_oc8051_idata_n848, oc8051_ram_top1_oc8051_idata_n847,
         oc8051_ram_top1_oc8051_idata_n846, oc8051_ram_top1_oc8051_idata_n845,
         oc8051_ram_top1_oc8051_idata_n844, oc8051_ram_top1_oc8051_idata_n843,
         oc8051_ram_top1_oc8051_idata_n842, oc8051_ram_top1_oc8051_idata_n841,
         oc8051_ram_top1_oc8051_idata_n840, oc8051_ram_top1_oc8051_idata_n839,
         oc8051_ram_top1_oc8051_idata_n838, oc8051_ram_top1_oc8051_idata_n837,
         oc8051_ram_top1_oc8051_idata_n836, oc8051_ram_top1_oc8051_idata_n835,
         oc8051_ram_top1_oc8051_idata_n834, oc8051_ram_top1_oc8051_idata_n833,
         oc8051_ram_top1_oc8051_idata_n832, oc8051_ram_top1_oc8051_idata_n831,
         oc8051_ram_top1_oc8051_idata_n830, oc8051_ram_top1_oc8051_idata_n829,
         oc8051_ram_top1_oc8051_idata_n828, oc8051_ram_top1_oc8051_idata_n827,
         oc8051_ram_top1_oc8051_idata_n826, oc8051_ram_top1_oc8051_idata_n825,
         oc8051_ram_top1_oc8051_idata_n824, oc8051_ram_top1_oc8051_idata_n823,
         oc8051_ram_top1_oc8051_idata_n822, oc8051_ram_top1_oc8051_idata_n821,
         oc8051_ram_top1_oc8051_idata_n820, oc8051_ram_top1_oc8051_idata_n819,
         oc8051_ram_top1_oc8051_idata_n818, oc8051_ram_top1_oc8051_idata_n817,
         oc8051_ram_top1_oc8051_idata_n816, oc8051_ram_top1_oc8051_idata_n815,
         oc8051_ram_top1_oc8051_idata_n814, oc8051_ram_top1_oc8051_idata_n813,
         oc8051_ram_top1_oc8051_idata_n812, oc8051_ram_top1_oc8051_idata_n811,
         oc8051_ram_top1_oc8051_idata_n810, oc8051_ram_top1_oc8051_idata_n809,
         oc8051_ram_top1_oc8051_idata_n808, oc8051_ram_top1_oc8051_idata_n807,
         oc8051_ram_top1_oc8051_idata_n806, oc8051_ram_top1_oc8051_idata_n805,
         oc8051_ram_top1_oc8051_idata_n804, oc8051_ram_top1_oc8051_idata_n803,
         oc8051_ram_top1_oc8051_idata_n802, oc8051_ram_top1_oc8051_idata_n801,
         oc8051_ram_top1_oc8051_idata_n800, oc8051_ram_top1_oc8051_idata_n799,
         oc8051_ram_top1_oc8051_idata_n798, oc8051_ram_top1_oc8051_idata_n797,
         oc8051_ram_top1_oc8051_idata_n796, oc8051_ram_top1_oc8051_idata_n795,
         oc8051_ram_top1_oc8051_idata_n794, oc8051_ram_top1_oc8051_idata_n793,
         oc8051_ram_top1_oc8051_idata_n792, oc8051_ram_top1_oc8051_idata_n791,
         oc8051_ram_top1_oc8051_idata_n790, oc8051_ram_top1_oc8051_idata_n789,
         oc8051_ram_top1_oc8051_idata_n788, oc8051_ram_top1_oc8051_idata_n787,
         oc8051_ram_top1_oc8051_idata_n786, oc8051_ram_top1_oc8051_idata_n785,
         oc8051_ram_top1_oc8051_idata_n784, oc8051_ram_top1_oc8051_idata_n783,
         oc8051_ram_top1_oc8051_idata_n782, oc8051_ram_top1_oc8051_idata_n781,
         oc8051_ram_top1_oc8051_idata_n780, oc8051_ram_top1_oc8051_idata_n779,
         oc8051_ram_top1_oc8051_idata_n778, oc8051_ram_top1_oc8051_idata_n777,
         oc8051_ram_top1_oc8051_idata_n776, oc8051_ram_top1_oc8051_idata_n775,
         oc8051_ram_top1_oc8051_idata_n774, oc8051_ram_top1_oc8051_idata_n773,
         oc8051_ram_top1_oc8051_idata_n772, oc8051_ram_top1_oc8051_idata_n771,
         oc8051_ram_top1_oc8051_idata_n770, oc8051_ram_top1_oc8051_idata_n769,
         oc8051_ram_top1_oc8051_idata_n768, oc8051_ram_top1_oc8051_idata_n767,
         oc8051_ram_top1_oc8051_idata_n766, oc8051_ram_top1_oc8051_idata_n765,
         oc8051_ram_top1_oc8051_idata_n764, oc8051_ram_top1_oc8051_idata_n763,
         oc8051_ram_top1_oc8051_idata_n762, oc8051_ram_top1_oc8051_idata_n761,
         oc8051_ram_top1_oc8051_idata_n760, oc8051_ram_top1_oc8051_idata_n759,
         oc8051_ram_top1_oc8051_idata_n758, oc8051_ram_top1_oc8051_idata_n757,
         oc8051_ram_top1_oc8051_idata_n756, oc8051_ram_top1_oc8051_idata_n755,
         oc8051_ram_top1_oc8051_idata_n754, oc8051_ram_top1_oc8051_idata_n753,
         oc8051_ram_top1_oc8051_idata_n752, oc8051_ram_top1_oc8051_idata_n751,
         oc8051_ram_top1_oc8051_idata_n750, oc8051_ram_top1_oc8051_idata_n749,
         oc8051_ram_top1_oc8051_idata_n748, oc8051_ram_top1_oc8051_idata_n747,
         oc8051_ram_top1_oc8051_idata_n746, oc8051_ram_top1_oc8051_idata_n745,
         oc8051_ram_top1_oc8051_idata_n744, oc8051_ram_top1_oc8051_idata_n743,
         oc8051_ram_top1_oc8051_idata_n742, oc8051_ram_top1_oc8051_idata_n741,
         oc8051_ram_top1_oc8051_idata_n740, oc8051_ram_top1_oc8051_idata_n739,
         oc8051_ram_top1_oc8051_idata_n738, oc8051_ram_top1_oc8051_idata_n737,
         oc8051_ram_top1_oc8051_idata_n736, oc8051_ram_top1_oc8051_idata_n735,
         oc8051_ram_top1_oc8051_idata_n734, oc8051_ram_top1_oc8051_idata_n733,
         oc8051_ram_top1_oc8051_idata_n732, oc8051_ram_top1_oc8051_idata_n731,
         oc8051_ram_top1_oc8051_idata_n730, oc8051_ram_top1_oc8051_idata_n729,
         oc8051_ram_top1_oc8051_idata_n728, oc8051_ram_top1_oc8051_idata_n727,
         oc8051_ram_top1_oc8051_idata_n726, oc8051_ram_top1_oc8051_idata_n725,
         oc8051_ram_top1_oc8051_idata_n724, oc8051_ram_top1_oc8051_idata_n723,
         oc8051_ram_top1_oc8051_idata_n722, oc8051_ram_top1_oc8051_idata_n721,
         oc8051_ram_top1_oc8051_idata_n720, oc8051_ram_top1_oc8051_idata_n719,
         oc8051_ram_top1_oc8051_idata_n718, oc8051_ram_top1_oc8051_idata_n717,
         oc8051_ram_top1_oc8051_idata_n716, oc8051_ram_top1_oc8051_idata_n715,
         oc8051_ram_top1_oc8051_idata_n714, oc8051_ram_top1_oc8051_idata_n713,
         oc8051_ram_top1_oc8051_idata_n712, oc8051_ram_top1_oc8051_idata_n711,
         oc8051_ram_top1_oc8051_idata_n710, oc8051_ram_top1_oc8051_idata_n709,
         oc8051_ram_top1_oc8051_idata_n708, oc8051_ram_top1_oc8051_idata_n707,
         oc8051_ram_top1_oc8051_idata_n706, oc8051_ram_top1_oc8051_idata_n705,
         oc8051_ram_top1_oc8051_idata_n704, oc8051_ram_top1_oc8051_idata_n703,
         oc8051_ram_top1_oc8051_idata_n702, oc8051_ram_top1_oc8051_idata_n701,
         oc8051_ram_top1_oc8051_idata_n700, oc8051_ram_top1_oc8051_idata_n699,
         oc8051_ram_top1_oc8051_idata_n698, oc8051_ram_top1_oc8051_idata_n697,
         oc8051_ram_top1_oc8051_idata_n696, oc8051_ram_top1_oc8051_idata_n695,
         oc8051_ram_top1_oc8051_idata_n694, oc8051_ram_top1_oc8051_idata_n693,
         oc8051_ram_top1_oc8051_idata_n692, oc8051_ram_top1_oc8051_idata_n691,
         oc8051_ram_top1_oc8051_idata_n690, oc8051_ram_top1_oc8051_idata_n689,
         oc8051_ram_top1_oc8051_idata_n688, oc8051_ram_top1_oc8051_idata_n687,
         oc8051_ram_top1_oc8051_idata_n686, oc8051_ram_top1_oc8051_idata_n685,
         oc8051_ram_top1_oc8051_idata_n684, oc8051_ram_top1_oc8051_idata_n683,
         oc8051_ram_top1_oc8051_idata_n682, oc8051_ram_top1_oc8051_idata_n681,
         oc8051_ram_top1_oc8051_idata_n680, oc8051_ram_top1_oc8051_idata_n679,
         oc8051_ram_top1_oc8051_idata_n678, oc8051_ram_top1_oc8051_idata_n677,
         oc8051_ram_top1_oc8051_idata_n676, oc8051_ram_top1_oc8051_idata_n675,
         oc8051_ram_top1_oc8051_idata_n674, oc8051_ram_top1_oc8051_idata_n673,
         oc8051_ram_top1_oc8051_idata_n672, oc8051_ram_top1_oc8051_idata_n671,
         oc8051_ram_top1_oc8051_idata_n670, oc8051_ram_top1_oc8051_idata_n669,
         oc8051_ram_top1_oc8051_idata_n668, oc8051_ram_top1_oc8051_idata_n667,
         oc8051_ram_top1_oc8051_idata_n666, oc8051_ram_top1_oc8051_idata_n665,
         oc8051_ram_top1_oc8051_idata_n664, oc8051_ram_top1_oc8051_idata_n663,
         oc8051_ram_top1_oc8051_idata_n662, oc8051_ram_top1_oc8051_idata_n661,
         oc8051_ram_top1_oc8051_idata_n660, oc8051_ram_top1_oc8051_idata_n659,
         oc8051_ram_top1_oc8051_idata_n658, oc8051_ram_top1_oc8051_idata_n657,
         oc8051_ram_top1_oc8051_idata_n656, oc8051_ram_top1_oc8051_idata_n655,
         oc8051_ram_top1_oc8051_idata_n654, oc8051_ram_top1_oc8051_idata_n653,
         oc8051_ram_top1_oc8051_idata_n652, oc8051_ram_top1_oc8051_idata_n651,
         oc8051_ram_top1_oc8051_idata_n650, oc8051_ram_top1_oc8051_idata_n649,
         oc8051_ram_top1_oc8051_idata_n648, oc8051_ram_top1_oc8051_idata_n647,
         oc8051_ram_top1_oc8051_idata_n646, oc8051_ram_top1_oc8051_idata_n645,
         oc8051_ram_top1_oc8051_idata_n644, oc8051_ram_top1_oc8051_idata_n643,
         oc8051_ram_top1_oc8051_idata_n642, oc8051_ram_top1_oc8051_idata_n641,
         oc8051_ram_top1_oc8051_idata_n640, oc8051_ram_top1_oc8051_idata_n639,
         oc8051_ram_top1_oc8051_idata_n638, oc8051_ram_top1_oc8051_idata_n637,
         oc8051_ram_top1_oc8051_idata_n636, oc8051_ram_top1_oc8051_idata_n635,
         oc8051_ram_top1_oc8051_idata_n634, oc8051_ram_top1_oc8051_idata_n633,
         oc8051_ram_top1_oc8051_idata_n632, oc8051_ram_top1_oc8051_idata_n631,
         oc8051_ram_top1_oc8051_idata_n630, oc8051_ram_top1_oc8051_idata_n629,
         oc8051_ram_top1_oc8051_idata_n628, oc8051_ram_top1_oc8051_idata_n627,
         oc8051_ram_top1_oc8051_idata_n626, oc8051_ram_top1_oc8051_idata_n625,
         oc8051_ram_top1_oc8051_idata_n624, oc8051_ram_top1_oc8051_idata_n623,
         oc8051_ram_top1_oc8051_idata_n622, oc8051_ram_top1_oc8051_idata_n621,
         oc8051_ram_top1_oc8051_idata_n620, oc8051_ram_top1_oc8051_idata_n619,
         oc8051_ram_top1_oc8051_idata_n618, oc8051_ram_top1_oc8051_idata_n617,
         oc8051_ram_top1_oc8051_idata_n616, oc8051_ram_top1_oc8051_idata_n615,
         oc8051_ram_top1_oc8051_idata_n614, oc8051_ram_top1_oc8051_idata_n613,
         oc8051_ram_top1_oc8051_idata_n612, oc8051_ram_top1_oc8051_idata_n611,
         oc8051_ram_top1_oc8051_idata_n610, oc8051_ram_top1_oc8051_idata_n609,
         oc8051_ram_top1_oc8051_idata_n608, oc8051_ram_top1_oc8051_idata_n607,
         oc8051_ram_top1_oc8051_idata_n606, oc8051_ram_top1_oc8051_idata_n605,
         oc8051_ram_top1_oc8051_idata_n604, oc8051_ram_top1_oc8051_idata_n603,
         oc8051_ram_top1_oc8051_idata_n602, oc8051_ram_top1_oc8051_idata_n601,
         oc8051_ram_top1_oc8051_idata_n600, oc8051_ram_top1_oc8051_idata_n599,
         oc8051_ram_top1_oc8051_idata_n598, oc8051_ram_top1_oc8051_idata_n597,
         oc8051_ram_top1_oc8051_idata_n596, oc8051_ram_top1_oc8051_idata_n595,
         oc8051_ram_top1_oc8051_idata_n594, oc8051_ram_top1_oc8051_idata_n593,
         oc8051_ram_top1_oc8051_idata_n592, oc8051_ram_top1_oc8051_idata_n591,
         oc8051_ram_top1_oc8051_idata_n590, oc8051_ram_top1_oc8051_idata_n589,
         oc8051_ram_top1_oc8051_idata_n588, oc8051_ram_top1_oc8051_idata_n587,
         oc8051_ram_top1_oc8051_idata_n586, oc8051_ram_top1_oc8051_idata_n585,
         oc8051_ram_top1_oc8051_idata_n584, oc8051_ram_top1_oc8051_idata_n583,
         oc8051_ram_top1_oc8051_idata_n582, oc8051_ram_top1_oc8051_idata_n581,
         oc8051_ram_top1_oc8051_idata_n580, oc8051_ram_top1_oc8051_idata_n579,
         oc8051_ram_top1_oc8051_idata_n578, oc8051_ram_top1_oc8051_idata_n577,
         oc8051_ram_top1_oc8051_idata_n576, oc8051_ram_top1_oc8051_idata_n575,
         oc8051_ram_top1_oc8051_idata_n574, oc8051_ram_top1_oc8051_idata_n573,
         oc8051_ram_top1_oc8051_idata_n572, oc8051_ram_top1_oc8051_idata_n571,
         oc8051_ram_top1_oc8051_idata_n570, oc8051_ram_top1_oc8051_idata_n569,
         oc8051_ram_top1_oc8051_idata_n568, oc8051_ram_top1_oc8051_idata_n567,
         oc8051_ram_top1_oc8051_idata_n566, oc8051_ram_top1_oc8051_idata_n565,
         oc8051_ram_top1_oc8051_idata_n564, oc8051_ram_top1_oc8051_idata_n563,
         oc8051_ram_top1_oc8051_idata_n562, oc8051_ram_top1_oc8051_idata_n561,
         oc8051_ram_top1_oc8051_idata_n560, oc8051_ram_top1_oc8051_idata_n559,
         oc8051_ram_top1_oc8051_idata_n558, oc8051_ram_top1_oc8051_idata_n557,
         oc8051_ram_top1_oc8051_idata_n556, oc8051_ram_top1_oc8051_idata_n555,
         oc8051_ram_top1_oc8051_idata_n554, oc8051_ram_top1_oc8051_idata_n553,
         oc8051_ram_top1_oc8051_idata_n552, oc8051_ram_top1_oc8051_idata_n551,
         oc8051_ram_top1_oc8051_idata_n550, oc8051_ram_top1_oc8051_idata_n549,
         oc8051_ram_top1_oc8051_idata_n548, oc8051_ram_top1_oc8051_idata_n547,
         oc8051_ram_top1_oc8051_idata_n546, oc8051_ram_top1_oc8051_idata_n545,
         oc8051_ram_top1_oc8051_idata_n544, oc8051_ram_top1_oc8051_idata_n543,
         oc8051_ram_top1_oc8051_idata_n542, oc8051_ram_top1_oc8051_idata_n541,
         oc8051_ram_top1_oc8051_idata_n540, oc8051_ram_top1_oc8051_idata_n539,
         oc8051_ram_top1_oc8051_idata_n538, oc8051_ram_top1_oc8051_idata_n537,
         oc8051_ram_top1_oc8051_idata_n536, oc8051_ram_top1_oc8051_idata_n535,
         oc8051_ram_top1_oc8051_idata_n534, oc8051_ram_top1_oc8051_idata_n533,
         oc8051_ram_top1_oc8051_idata_n532, oc8051_ram_top1_oc8051_idata_n531,
         oc8051_ram_top1_oc8051_idata_n530, oc8051_ram_top1_oc8051_idata_n529,
         oc8051_ram_top1_oc8051_idata_n528, oc8051_ram_top1_oc8051_idata_n527,
         oc8051_ram_top1_oc8051_idata_n526, oc8051_ram_top1_oc8051_idata_n525,
         oc8051_ram_top1_oc8051_idata_n524, oc8051_ram_top1_oc8051_idata_n523,
         oc8051_ram_top1_oc8051_idata_n522, oc8051_ram_top1_oc8051_idata_n521,
         oc8051_ram_top1_oc8051_idata_n520, oc8051_ram_top1_oc8051_idata_n519,
         oc8051_ram_top1_oc8051_idata_n518, oc8051_ram_top1_oc8051_idata_n517,
         oc8051_ram_top1_oc8051_idata_n516, oc8051_ram_top1_oc8051_idata_n3,
         oc8051_ram_top1_oc8051_idata_n2, oc8051_ram_top1_oc8051_idata_n1,
         oc8051_ram_top1_oc8051_idata_n4530,
         oc8051_ram_top1_oc8051_idata_n4529,
         oc8051_ram_top1_oc8051_idata_n4528,
         oc8051_ram_top1_oc8051_idata_n4527,
         oc8051_ram_top1_oc8051_idata_n4526,
         oc8051_ram_top1_oc8051_idata_n4525,
         oc8051_ram_top1_oc8051_idata_n4524,
         oc8051_ram_top1_oc8051_idata_n4523,
         oc8051_ram_top1_oc8051_idata_n4522,
         oc8051_ram_top1_oc8051_idata_n4521,
         oc8051_ram_top1_oc8051_idata_n4520,
         oc8051_ram_top1_oc8051_idata_n4519,
         oc8051_ram_top1_oc8051_idata_n4518,
         oc8051_ram_top1_oc8051_idata_n4517,
         oc8051_ram_top1_oc8051_idata_n4516,
         oc8051_ram_top1_oc8051_idata_n4515,
         oc8051_ram_top1_oc8051_idata_n4514,
         oc8051_ram_top1_oc8051_idata_n4513,
         oc8051_ram_top1_oc8051_idata_n4512,
         oc8051_ram_top1_oc8051_idata_n4511,
         oc8051_ram_top1_oc8051_idata_n4510,
         oc8051_ram_top1_oc8051_idata_n4509,
         oc8051_ram_top1_oc8051_idata_n4508,
         oc8051_ram_top1_oc8051_idata_n4507,
         oc8051_ram_top1_oc8051_idata_n4506,
         oc8051_ram_top1_oc8051_idata_n4505,
         oc8051_ram_top1_oc8051_idata_n4504,
         oc8051_ram_top1_oc8051_idata_n4503,
         oc8051_ram_top1_oc8051_idata_n4502,
         oc8051_ram_top1_oc8051_idata_n4501,
         oc8051_ram_top1_oc8051_idata_n4500,
         oc8051_ram_top1_oc8051_idata_n4499,
         oc8051_ram_top1_oc8051_idata_n4498,
         oc8051_ram_top1_oc8051_idata_n4497,
         oc8051_ram_top1_oc8051_idata_n4496,
         oc8051_ram_top1_oc8051_idata_n4495,
         oc8051_ram_top1_oc8051_idata_n4494,
         oc8051_ram_top1_oc8051_idata_n4493,
         oc8051_ram_top1_oc8051_idata_n4492,
         oc8051_ram_top1_oc8051_idata_n4491,
         oc8051_ram_top1_oc8051_idata_n4490,
         oc8051_ram_top1_oc8051_idata_n4489,
         oc8051_ram_top1_oc8051_idata_n4488,
         oc8051_ram_top1_oc8051_idata_n4487,
         oc8051_ram_top1_oc8051_idata_n4486,
         oc8051_ram_top1_oc8051_idata_n4485,
         oc8051_ram_top1_oc8051_idata_n4484,
         oc8051_ram_top1_oc8051_idata_n4483,
         oc8051_ram_top1_oc8051_idata_n4482,
         oc8051_ram_top1_oc8051_idata_n4481,
         oc8051_ram_top1_oc8051_idata_n4480,
         oc8051_ram_top1_oc8051_idata_n4479,
         oc8051_ram_top1_oc8051_idata_n4478,
         oc8051_ram_top1_oc8051_idata_n4477,
         oc8051_ram_top1_oc8051_idata_n4476,
         oc8051_ram_top1_oc8051_idata_n4475,
         oc8051_ram_top1_oc8051_idata_n4474,
         oc8051_ram_top1_oc8051_idata_n4473,
         oc8051_ram_top1_oc8051_idata_n4472,
         oc8051_ram_top1_oc8051_idata_n4471,
         oc8051_ram_top1_oc8051_idata_n4470,
         oc8051_ram_top1_oc8051_idata_n4469,
         oc8051_ram_top1_oc8051_idata_n4468,
         oc8051_ram_top1_oc8051_idata_n4467,
         oc8051_ram_top1_oc8051_idata_n4466,
         oc8051_ram_top1_oc8051_idata_n4465,
         oc8051_ram_top1_oc8051_idata_n4464,
         oc8051_ram_top1_oc8051_idata_n4463,
         oc8051_ram_top1_oc8051_idata_n4462,
         oc8051_ram_top1_oc8051_idata_n4461,
         oc8051_ram_top1_oc8051_idata_n4460,
         oc8051_ram_top1_oc8051_idata_n4459,
         oc8051_ram_top1_oc8051_idata_n4458,
         oc8051_ram_top1_oc8051_idata_n4457,
         oc8051_ram_top1_oc8051_idata_n4456,
         oc8051_ram_top1_oc8051_idata_n4455,
         oc8051_ram_top1_oc8051_idata_n4454,
         oc8051_ram_top1_oc8051_idata_n4453,
         oc8051_ram_top1_oc8051_idata_n4452,
         oc8051_ram_top1_oc8051_idata_n4451,
         oc8051_ram_top1_oc8051_idata_n4450,
         oc8051_ram_top1_oc8051_idata_n4449,
         oc8051_ram_top1_oc8051_idata_n4448,
         oc8051_ram_top1_oc8051_idata_n4447,
         oc8051_ram_top1_oc8051_idata_n4446,
         oc8051_ram_top1_oc8051_idata_n4445,
         oc8051_ram_top1_oc8051_idata_n4444,
         oc8051_ram_top1_oc8051_idata_n4443,
         oc8051_ram_top1_oc8051_idata_n4442,
         oc8051_ram_top1_oc8051_idata_n4441,
         oc8051_ram_top1_oc8051_idata_n4440,
         oc8051_ram_top1_oc8051_idata_n4439,
         oc8051_ram_top1_oc8051_idata_n4438,
         oc8051_ram_top1_oc8051_idata_n4437,
         oc8051_ram_top1_oc8051_idata_n4436,
         oc8051_ram_top1_oc8051_idata_n4435,
         oc8051_ram_top1_oc8051_idata_n4434,
         oc8051_ram_top1_oc8051_idata_n4433,
         oc8051_ram_top1_oc8051_idata_n4432,
         oc8051_ram_top1_oc8051_idata_n4431,
         oc8051_ram_top1_oc8051_idata_n4430,
         oc8051_ram_top1_oc8051_idata_n4429,
         oc8051_ram_top1_oc8051_idata_n4428,
         oc8051_ram_top1_oc8051_idata_n4427,
         oc8051_ram_top1_oc8051_idata_n4426,
         oc8051_ram_top1_oc8051_idata_n4425,
         oc8051_ram_top1_oc8051_idata_n4424,
         oc8051_ram_top1_oc8051_idata_n4423,
         oc8051_ram_top1_oc8051_idata_n4422,
         oc8051_ram_top1_oc8051_idata_n4421,
         oc8051_ram_top1_oc8051_idata_n4420,
         oc8051_ram_top1_oc8051_idata_n4419,
         oc8051_ram_top1_oc8051_idata_n4418,
         oc8051_ram_top1_oc8051_idata_n4417,
         oc8051_ram_top1_oc8051_idata_n4416,
         oc8051_ram_top1_oc8051_idata_n4415,
         oc8051_ram_top1_oc8051_idata_n4414,
         oc8051_ram_top1_oc8051_idata_n4413,
         oc8051_ram_top1_oc8051_idata_n4412,
         oc8051_ram_top1_oc8051_idata_n4411,
         oc8051_ram_top1_oc8051_idata_n4410,
         oc8051_ram_top1_oc8051_idata_n4409,
         oc8051_ram_top1_oc8051_idata_n4408,
         oc8051_ram_top1_oc8051_idata_n4407,
         oc8051_ram_top1_oc8051_idata_n4406,
         oc8051_ram_top1_oc8051_idata_n4405,
         oc8051_ram_top1_oc8051_idata_n4404,
         oc8051_ram_top1_oc8051_idata_n4403,
         oc8051_ram_top1_oc8051_idata_n4402,
         oc8051_ram_top1_oc8051_idata_n4401,
         oc8051_ram_top1_oc8051_idata_n4400,
         oc8051_ram_top1_oc8051_idata_n4399,
         oc8051_ram_top1_oc8051_idata_n4398,
         oc8051_ram_top1_oc8051_idata_n4397,
         oc8051_ram_top1_oc8051_idata_n4396,
         oc8051_ram_top1_oc8051_idata_n4395,
         oc8051_ram_top1_oc8051_idata_n4394,
         oc8051_ram_top1_oc8051_idata_n4393,
         oc8051_ram_top1_oc8051_idata_n4392,
         oc8051_ram_top1_oc8051_idata_n4391,
         oc8051_ram_top1_oc8051_idata_n4390,
         oc8051_ram_top1_oc8051_idata_n4389,
         oc8051_ram_top1_oc8051_idata_n4388,
         oc8051_ram_top1_oc8051_idata_n4387,
         oc8051_ram_top1_oc8051_idata_n4386,
         oc8051_ram_top1_oc8051_idata_n4385,
         oc8051_ram_top1_oc8051_idata_n4384,
         oc8051_ram_top1_oc8051_idata_n4383,
         oc8051_ram_top1_oc8051_idata_n4382,
         oc8051_ram_top1_oc8051_idata_n4381,
         oc8051_ram_top1_oc8051_idata_n4380,
         oc8051_ram_top1_oc8051_idata_n4379,
         oc8051_ram_top1_oc8051_idata_n4378,
         oc8051_ram_top1_oc8051_idata_n4377,
         oc8051_ram_top1_oc8051_idata_n4376,
         oc8051_ram_top1_oc8051_idata_n4375,
         oc8051_ram_top1_oc8051_idata_n4374,
         oc8051_ram_top1_oc8051_idata_n4373,
         oc8051_ram_top1_oc8051_idata_n4372,
         oc8051_ram_top1_oc8051_idata_n4371,
         oc8051_ram_top1_oc8051_idata_n4370,
         oc8051_ram_top1_oc8051_idata_n4369,
         oc8051_ram_top1_oc8051_idata_n4368,
         oc8051_ram_top1_oc8051_idata_n4367,
         oc8051_ram_top1_oc8051_idata_n4366,
         oc8051_ram_top1_oc8051_idata_n4365,
         oc8051_ram_top1_oc8051_idata_n4364,
         oc8051_ram_top1_oc8051_idata_n4363,
         oc8051_ram_top1_oc8051_idata_n4362,
         oc8051_ram_top1_oc8051_idata_n4361,
         oc8051_ram_top1_oc8051_idata_n4360,
         oc8051_ram_top1_oc8051_idata_n4359,
         oc8051_ram_top1_oc8051_idata_n4358,
         oc8051_ram_top1_oc8051_idata_n4357,
         oc8051_ram_top1_oc8051_idata_n4356,
         oc8051_ram_top1_oc8051_idata_n4355,
         oc8051_ram_top1_oc8051_idata_n4354,
         oc8051_ram_top1_oc8051_idata_n4353,
         oc8051_ram_top1_oc8051_idata_n4352,
         oc8051_ram_top1_oc8051_idata_n4351,
         oc8051_ram_top1_oc8051_idata_n4350,
         oc8051_ram_top1_oc8051_idata_n4349,
         oc8051_ram_top1_oc8051_idata_n4348,
         oc8051_ram_top1_oc8051_idata_n4347,
         oc8051_ram_top1_oc8051_idata_n4346,
         oc8051_ram_top1_oc8051_idata_n4345,
         oc8051_ram_top1_oc8051_idata_n4344,
         oc8051_ram_top1_oc8051_idata_n4343,
         oc8051_ram_top1_oc8051_idata_n4342,
         oc8051_ram_top1_oc8051_idata_n4341,
         oc8051_ram_top1_oc8051_idata_n4340,
         oc8051_ram_top1_oc8051_idata_n4339,
         oc8051_ram_top1_oc8051_idata_n4338,
         oc8051_ram_top1_oc8051_idata_n4337,
         oc8051_ram_top1_oc8051_idata_n4336,
         oc8051_ram_top1_oc8051_idata_n4335,
         oc8051_ram_top1_oc8051_idata_n4334,
         oc8051_ram_top1_oc8051_idata_n4333,
         oc8051_ram_top1_oc8051_idata_n4332,
         oc8051_ram_top1_oc8051_idata_n4331,
         oc8051_ram_top1_oc8051_idata_n4330,
         oc8051_ram_top1_oc8051_idata_n4329,
         oc8051_ram_top1_oc8051_idata_n4328,
         oc8051_ram_top1_oc8051_idata_n4327,
         oc8051_ram_top1_oc8051_idata_n4326,
         oc8051_ram_top1_oc8051_idata_n4325,
         oc8051_ram_top1_oc8051_idata_n4324,
         oc8051_ram_top1_oc8051_idata_n4323,
         oc8051_ram_top1_oc8051_idata_n4322,
         oc8051_ram_top1_oc8051_idata_n4321,
         oc8051_ram_top1_oc8051_idata_n4320,
         oc8051_ram_top1_oc8051_idata_n4319,
         oc8051_ram_top1_oc8051_idata_n4318,
         oc8051_ram_top1_oc8051_idata_n4317,
         oc8051_ram_top1_oc8051_idata_n4316,
         oc8051_ram_top1_oc8051_idata_n4315,
         oc8051_ram_top1_oc8051_idata_n4314,
         oc8051_ram_top1_oc8051_idata_n4313,
         oc8051_ram_top1_oc8051_idata_n4312,
         oc8051_ram_top1_oc8051_idata_n4311,
         oc8051_ram_top1_oc8051_idata_n4310,
         oc8051_ram_top1_oc8051_idata_n4309,
         oc8051_ram_top1_oc8051_idata_n4308,
         oc8051_ram_top1_oc8051_idata_n4307,
         oc8051_ram_top1_oc8051_idata_n4306,
         oc8051_ram_top1_oc8051_idata_n4305,
         oc8051_ram_top1_oc8051_idata_n4304,
         oc8051_ram_top1_oc8051_idata_n4303,
         oc8051_ram_top1_oc8051_idata_n4302,
         oc8051_ram_top1_oc8051_idata_n4301,
         oc8051_ram_top1_oc8051_idata_n4300,
         oc8051_ram_top1_oc8051_idata_n4299,
         oc8051_ram_top1_oc8051_idata_n4298,
         oc8051_ram_top1_oc8051_idata_n4297,
         oc8051_ram_top1_oc8051_idata_n4296,
         oc8051_ram_top1_oc8051_idata_n4295,
         oc8051_ram_top1_oc8051_idata_n4294,
         oc8051_ram_top1_oc8051_idata_n4293,
         oc8051_ram_top1_oc8051_idata_n4292,
         oc8051_ram_top1_oc8051_idata_n4291,
         oc8051_ram_top1_oc8051_idata_n4290,
         oc8051_ram_top1_oc8051_idata_n4289,
         oc8051_ram_top1_oc8051_idata_n4288,
         oc8051_ram_top1_oc8051_idata_n4287,
         oc8051_ram_top1_oc8051_idata_n4286,
         oc8051_ram_top1_oc8051_idata_n4285,
         oc8051_ram_top1_oc8051_idata_n4284,
         oc8051_ram_top1_oc8051_idata_n4283,
         oc8051_ram_top1_oc8051_idata_n4282,
         oc8051_ram_top1_oc8051_idata_n4281,
         oc8051_ram_top1_oc8051_idata_n4280,
         oc8051_ram_top1_oc8051_idata_n4279,
         oc8051_ram_top1_oc8051_idata_n4278,
         oc8051_ram_top1_oc8051_idata_n4277,
         oc8051_ram_top1_oc8051_idata_n4276,
         oc8051_ram_top1_oc8051_idata_n4275,
         oc8051_ram_top1_oc8051_idata_n4274,
         oc8051_ram_top1_oc8051_idata_n4273,
         oc8051_ram_top1_oc8051_idata_n4272,
         oc8051_ram_top1_oc8051_idata_n4271,
         oc8051_ram_top1_oc8051_idata_n4270,
         oc8051_ram_top1_oc8051_idata_n4269,
         oc8051_ram_top1_oc8051_idata_n4268,
         oc8051_ram_top1_oc8051_idata_n4267,
         oc8051_ram_top1_oc8051_idata_n4266,
         oc8051_ram_top1_oc8051_idata_n4265,
         oc8051_ram_top1_oc8051_idata_n4264,
         oc8051_ram_top1_oc8051_idata_n4263,
         oc8051_ram_top1_oc8051_idata_n4262,
         oc8051_ram_top1_oc8051_idata_n4261,
         oc8051_ram_top1_oc8051_idata_n4260,
         oc8051_ram_top1_oc8051_idata_n4259,
         oc8051_ram_top1_oc8051_idata_n4258,
         oc8051_ram_top1_oc8051_idata_n4257,
         oc8051_ram_top1_oc8051_idata_n4256,
         oc8051_ram_top1_oc8051_idata_n4255,
         oc8051_ram_top1_oc8051_idata_n4254,
         oc8051_ram_top1_oc8051_idata_n4253,
         oc8051_ram_top1_oc8051_idata_n4252,
         oc8051_ram_top1_oc8051_idata_n4251,
         oc8051_ram_top1_oc8051_idata_n4250,
         oc8051_ram_top1_oc8051_idata_n4249,
         oc8051_ram_top1_oc8051_idata_n4248,
         oc8051_ram_top1_oc8051_idata_n4247,
         oc8051_ram_top1_oc8051_idata_n4246,
         oc8051_ram_top1_oc8051_idata_n4245,
         oc8051_ram_top1_oc8051_idata_n4244,
         oc8051_ram_top1_oc8051_idata_n4243,
         oc8051_ram_top1_oc8051_idata_n4242,
         oc8051_ram_top1_oc8051_idata_n4241,
         oc8051_ram_top1_oc8051_idata_n4240,
         oc8051_ram_top1_oc8051_idata_n4239,
         oc8051_ram_top1_oc8051_idata_n4238,
         oc8051_ram_top1_oc8051_idata_n4237,
         oc8051_ram_top1_oc8051_idata_n4236,
         oc8051_ram_top1_oc8051_idata_n4235,
         oc8051_ram_top1_oc8051_idata_n4234,
         oc8051_ram_top1_oc8051_idata_n4233,
         oc8051_ram_top1_oc8051_idata_n4232,
         oc8051_ram_top1_oc8051_idata_n4231,
         oc8051_ram_top1_oc8051_idata_n4230,
         oc8051_ram_top1_oc8051_idata_n4229,
         oc8051_ram_top1_oc8051_idata_n4228,
         oc8051_ram_top1_oc8051_idata_n4227,
         oc8051_ram_top1_oc8051_idata_n4226,
         oc8051_ram_top1_oc8051_idata_n4225,
         oc8051_ram_top1_oc8051_idata_n4224,
         oc8051_ram_top1_oc8051_idata_n4223,
         oc8051_ram_top1_oc8051_idata_n4222,
         oc8051_ram_top1_oc8051_idata_n4221,
         oc8051_ram_top1_oc8051_idata_n4220,
         oc8051_ram_top1_oc8051_idata_n4219,
         oc8051_ram_top1_oc8051_idata_n4218,
         oc8051_ram_top1_oc8051_idata_n4217,
         oc8051_ram_top1_oc8051_idata_n4216,
         oc8051_ram_top1_oc8051_idata_n4215,
         oc8051_ram_top1_oc8051_idata_n4214,
         oc8051_ram_top1_oc8051_idata_n4213,
         oc8051_ram_top1_oc8051_idata_n4212,
         oc8051_ram_top1_oc8051_idata_n4211,
         oc8051_ram_top1_oc8051_idata_n4210,
         oc8051_ram_top1_oc8051_idata_n4209,
         oc8051_ram_top1_oc8051_idata_n4208,
         oc8051_ram_top1_oc8051_idata_n4207,
         oc8051_ram_top1_oc8051_idata_n4206,
         oc8051_ram_top1_oc8051_idata_n4205,
         oc8051_ram_top1_oc8051_idata_n4204,
         oc8051_ram_top1_oc8051_idata_n4203,
         oc8051_ram_top1_oc8051_idata_n4202,
         oc8051_ram_top1_oc8051_idata_n4201,
         oc8051_ram_top1_oc8051_idata_n4200,
         oc8051_ram_top1_oc8051_idata_n4199,
         oc8051_ram_top1_oc8051_idata_n4198,
         oc8051_ram_top1_oc8051_idata_n4197,
         oc8051_ram_top1_oc8051_idata_n4196,
         oc8051_ram_top1_oc8051_idata_n4195,
         oc8051_ram_top1_oc8051_idata_n4194,
         oc8051_ram_top1_oc8051_idata_n4193,
         oc8051_ram_top1_oc8051_idata_n4192,
         oc8051_ram_top1_oc8051_idata_n4191,
         oc8051_ram_top1_oc8051_idata_n4190,
         oc8051_ram_top1_oc8051_idata_n4189,
         oc8051_ram_top1_oc8051_idata_n4188,
         oc8051_ram_top1_oc8051_idata_n4187,
         oc8051_ram_top1_oc8051_idata_n4186,
         oc8051_ram_top1_oc8051_idata_n4185,
         oc8051_ram_top1_oc8051_idata_n4184,
         oc8051_ram_top1_oc8051_idata_n4183,
         oc8051_ram_top1_oc8051_idata_n4182,
         oc8051_ram_top1_oc8051_idata_n4181,
         oc8051_ram_top1_oc8051_idata_n4180,
         oc8051_ram_top1_oc8051_idata_n4179,
         oc8051_ram_top1_oc8051_idata_n4178,
         oc8051_ram_top1_oc8051_idata_n4177,
         oc8051_ram_top1_oc8051_idata_n4176,
         oc8051_ram_top1_oc8051_idata_n4175,
         oc8051_ram_top1_oc8051_idata_n4174,
         oc8051_ram_top1_oc8051_idata_n4173,
         oc8051_ram_top1_oc8051_idata_n4172,
         oc8051_ram_top1_oc8051_idata_n4171,
         oc8051_ram_top1_oc8051_idata_n4170,
         oc8051_ram_top1_oc8051_idata_n4169,
         oc8051_ram_top1_oc8051_idata_n4168,
         oc8051_ram_top1_oc8051_idata_n4167,
         oc8051_ram_top1_oc8051_idata_n4166,
         oc8051_ram_top1_oc8051_idata_n4165,
         oc8051_ram_top1_oc8051_idata_n4164,
         oc8051_ram_top1_oc8051_idata_n4163,
         oc8051_ram_top1_oc8051_idata_n4162,
         oc8051_ram_top1_oc8051_idata_n4161,
         oc8051_ram_top1_oc8051_idata_n4160,
         oc8051_ram_top1_oc8051_idata_n4159,
         oc8051_ram_top1_oc8051_idata_n4158,
         oc8051_ram_top1_oc8051_idata_n4157,
         oc8051_ram_top1_oc8051_idata_n4156,
         oc8051_ram_top1_oc8051_idata_n4155,
         oc8051_ram_top1_oc8051_idata_n4154,
         oc8051_ram_top1_oc8051_idata_n4153,
         oc8051_ram_top1_oc8051_idata_n4152,
         oc8051_ram_top1_oc8051_idata_n4151,
         oc8051_ram_top1_oc8051_idata_n4150,
         oc8051_ram_top1_oc8051_idata_n4149,
         oc8051_ram_top1_oc8051_idata_n4148,
         oc8051_ram_top1_oc8051_idata_n4147,
         oc8051_ram_top1_oc8051_idata_n4146,
         oc8051_ram_top1_oc8051_idata_n4145,
         oc8051_ram_top1_oc8051_idata_n4144,
         oc8051_ram_top1_oc8051_idata_n4143,
         oc8051_ram_top1_oc8051_idata_n4142,
         oc8051_ram_top1_oc8051_idata_n4141,
         oc8051_ram_top1_oc8051_idata_n4140,
         oc8051_ram_top1_oc8051_idata_n4139,
         oc8051_ram_top1_oc8051_idata_n4138,
         oc8051_ram_top1_oc8051_idata_n4137,
         oc8051_ram_top1_oc8051_idata_n4136,
         oc8051_ram_top1_oc8051_idata_n4135,
         oc8051_ram_top1_oc8051_idata_n4134,
         oc8051_ram_top1_oc8051_idata_n4133,
         oc8051_ram_top1_oc8051_idata_n4132,
         oc8051_ram_top1_oc8051_idata_n4131,
         oc8051_ram_top1_oc8051_idata_n4130,
         oc8051_ram_top1_oc8051_idata_n4129,
         oc8051_ram_top1_oc8051_idata_n4128,
         oc8051_ram_top1_oc8051_idata_n4127,
         oc8051_ram_top1_oc8051_idata_n4126,
         oc8051_ram_top1_oc8051_idata_n4125,
         oc8051_ram_top1_oc8051_idata_n4124,
         oc8051_ram_top1_oc8051_idata_n4123,
         oc8051_ram_top1_oc8051_idata_n4122,
         oc8051_ram_top1_oc8051_idata_n4121,
         oc8051_ram_top1_oc8051_idata_n4120,
         oc8051_ram_top1_oc8051_idata_n4119,
         oc8051_ram_top1_oc8051_idata_n4118,
         oc8051_ram_top1_oc8051_idata_n4117,
         oc8051_ram_top1_oc8051_idata_n4116,
         oc8051_ram_top1_oc8051_idata_n4115,
         oc8051_ram_top1_oc8051_idata_n4114,
         oc8051_ram_top1_oc8051_idata_n4113,
         oc8051_ram_top1_oc8051_idata_n4112,
         oc8051_ram_top1_oc8051_idata_n4111,
         oc8051_ram_top1_oc8051_idata_n4110,
         oc8051_ram_top1_oc8051_idata_n4109,
         oc8051_ram_top1_oc8051_idata_n4108,
         oc8051_ram_top1_oc8051_idata_n4107,
         oc8051_ram_top1_oc8051_idata_n4106,
         oc8051_ram_top1_oc8051_idata_n4105,
         oc8051_ram_top1_oc8051_idata_n4104,
         oc8051_ram_top1_oc8051_idata_n4103,
         oc8051_ram_top1_oc8051_idata_n4102,
         oc8051_ram_top1_oc8051_idata_n4101,
         oc8051_ram_top1_oc8051_idata_n4100,
         oc8051_ram_top1_oc8051_idata_n4099,
         oc8051_ram_top1_oc8051_idata_n4098,
         oc8051_ram_top1_oc8051_idata_n4097,
         oc8051_ram_top1_oc8051_idata_n4096,
         oc8051_ram_top1_oc8051_idata_n4095,
         oc8051_ram_top1_oc8051_idata_n4094,
         oc8051_ram_top1_oc8051_idata_n4093,
         oc8051_ram_top1_oc8051_idata_n4092,
         oc8051_ram_top1_oc8051_idata_n4091,
         oc8051_ram_top1_oc8051_idata_n4090,
         oc8051_ram_top1_oc8051_idata_n4089,
         oc8051_ram_top1_oc8051_idata_n4088,
         oc8051_ram_top1_oc8051_idata_n4087,
         oc8051_ram_top1_oc8051_idata_n4086,
         oc8051_ram_top1_oc8051_idata_n4085,
         oc8051_ram_top1_oc8051_idata_n4084,
         oc8051_ram_top1_oc8051_idata_n4083,
         oc8051_ram_top1_oc8051_idata_n4082,
         oc8051_ram_top1_oc8051_idata_n4081,
         oc8051_ram_top1_oc8051_idata_n4080,
         oc8051_ram_top1_oc8051_idata_n4079,
         oc8051_ram_top1_oc8051_idata_n4078,
         oc8051_ram_top1_oc8051_idata_n4077,
         oc8051_ram_top1_oc8051_idata_n4076,
         oc8051_ram_top1_oc8051_idata_n4075,
         oc8051_ram_top1_oc8051_idata_n4074,
         oc8051_ram_top1_oc8051_idata_n4073,
         oc8051_ram_top1_oc8051_idata_n4072,
         oc8051_ram_top1_oc8051_idata_n4071,
         oc8051_ram_top1_oc8051_idata_n4070,
         oc8051_ram_top1_oc8051_idata_n4069,
         oc8051_ram_top1_oc8051_idata_n4068,
         oc8051_ram_top1_oc8051_idata_n4067,
         oc8051_ram_top1_oc8051_idata_n4066,
         oc8051_ram_top1_oc8051_idata_n4065,
         oc8051_ram_top1_oc8051_idata_n4064,
         oc8051_ram_top1_oc8051_idata_n4063,
         oc8051_ram_top1_oc8051_idata_n4062,
         oc8051_ram_top1_oc8051_idata_n4061,
         oc8051_ram_top1_oc8051_idata_n4060,
         oc8051_ram_top1_oc8051_idata_n4059,
         oc8051_ram_top1_oc8051_idata_n4058,
         oc8051_ram_top1_oc8051_idata_n4057,
         oc8051_ram_top1_oc8051_idata_n4056,
         oc8051_ram_top1_oc8051_idata_n4055,
         oc8051_ram_top1_oc8051_idata_n4054,
         oc8051_ram_top1_oc8051_idata_n4053,
         oc8051_ram_top1_oc8051_idata_n4052,
         oc8051_ram_top1_oc8051_idata_n4051,
         oc8051_ram_top1_oc8051_idata_n4050,
         oc8051_ram_top1_oc8051_idata_n4049,
         oc8051_ram_top1_oc8051_idata_n4048,
         oc8051_ram_top1_oc8051_idata_n4047,
         oc8051_ram_top1_oc8051_idata_n4046,
         oc8051_ram_top1_oc8051_idata_n4045,
         oc8051_ram_top1_oc8051_idata_n4044,
         oc8051_ram_top1_oc8051_idata_n4043,
         oc8051_ram_top1_oc8051_idata_n4042,
         oc8051_ram_top1_oc8051_idata_n4041,
         oc8051_ram_top1_oc8051_idata_n4040,
         oc8051_ram_top1_oc8051_idata_n4039,
         oc8051_ram_top1_oc8051_idata_n4038,
         oc8051_ram_top1_oc8051_idata_n4037,
         oc8051_ram_top1_oc8051_idata_n4036,
         oc8051_ram_top1_oc8051_idata_n4035,
         oc8051_ram_top1_oc8051_idata_n4034,
         oc8051_ram_top1_oc8051_idata_n4033,
         oc8051_ram_top1_oc8051_idata_n4032,
         oc8051_ram_top1_oc8051_idata_n4031,
         oc8051_ram_top1_oc8051_idata_n4030,
         oc8051_ram_top1_oc8051_idata_n4029,
         oc8051_ram_top1_oc8051_idata_n4028,
         oc8051_ram_top1_oc8051_idata_n4027,
         oc8051_ram_top1_oc8051_idata_n4026,
         oc8051_ram_top1_oc8051_idata_n4025,
         oc8051_ram_top1_oc8051_idata_n4024,
         oc8051_ram_top1_oc8051_idata_n4023,
         oc8051_ram_top1_oc8051_idata_n4022,
         oc8051_ram_top1_oc8051_idata_n4021,
         oc8051_ram_top1_oc8051_idata_n4020,
         oc8051_ram_top1_oc8051_idata_n4019,
         oc8051_ram_top1_oc8051_idata_n4018,
         oc8051_ram_top1_oc8051_idata_n4017,
         oc8051_ram_top1_oc8051_idata_n4016,
         oc8051_ram_top1_oc8051_idata_n4015,
         oc8051_ram_top1_oc8051_idata_n4014,
         oc8051_ram_top1_oc8051_idata_n4013,
         oc8051_ram_top1_oc8051_idata_n4012,
         oc8051_ram_top1_oc8051_idata_n4011,
         oc8051_ram_top1_oc8051_idata_n4010,
         oc8051_ram_top1_oc8051_idata_n4009,
         oc8051_ram_top1_oc8051_idata_n4008,
         oc8051_ram_top1_oc8051_idata_n4007,
         oc8051_ram_top1_oc8051_idata_n4006,
         oc8051_ram_top1_oc8051_idata_n4005,
         oc8051_ram_top1_oc8051_idata_n4004,
         oc8051_ram_top1_oc8051_idata_n4003,
         oc8051_ram_top1_oc8051_idata_n4002,
         oc8051_ram_top1_oc8051_idata_n4001,
         oc8051_ram_top1_oc8051_idata_n4000,
         oc8051_ram_top1_oc8051_idata_n3999,
         oc8051_ram_top1_oc8051_idata_n3998,
         oc8051_ram_top1_oc8051_idata_n3997,
         oc8051_ram_top1_oc8051_idata_n3996,
         oc8051_ram_top1_oc8051_idata_n3995,
         oc8051_ram_top1_oc8051_idata_n3994,
         oc8051_ram_top1_oc8051_idata_n3993,
         oc8051_ram_top1_oc8051_idata_n3992,
         oc8051_ram_top1_oc8051_idata_n3991,
         oc8051_ram_top1_oc8051_idata_n3990,
         oc8051_ram_top1_oc8051_idata_n3989,
         oc8051_ram_top1_oc8051_idata_n3988,
         oc8051_ram_top1_oc8051_idata_n3987,
         oc8051_ram_top1_oc8051_idata_n3986,
         oc8051_ram_top1_oc8051_idata_n3985,
         oc8051_ram_top1_oc8051_idata_n3984,
         oc8051_ram_top1_oc8051_idata_n3983,
         oc8051_ram_top1_oc8051_idata_n3982,
         oc8051_ram_top1_oc8051_idata_n3981,
         oc8051_ram_top1_oc8051_idata_n3980,
         oc8051_ram_top1_oc8051_idata_n3979,
         oc8051_ram_top1_oc8051_idata_n3978,
         oc8051_ram_top1_oc8051_idata_n3977,
         oc8051_ram_top1_oc8051_idata_n3976,
         oc8051_ram_top1_oc8051_idata_n3975,
         oc8051_ram_top1_oc8051_idata_n3974,
         oc8051_ram_top1_oc8051_idata_n3973,
         oc8051_ram_top1_oc8051_idata_n3972,
         oc8051_ram_top1_oc8051_idata_n3971,
         oc8051_ram_top1_oc8051_idata_n3970,
         oc8051_ram_top1_oc8051_idata_n3969,
         oc8051_ram_top1_oc8051_idata_n3968,
         oc8051_ram_top1_oc8051_idata_n3967,
         oc8051_ram_top1_oc8051_idata_n3966,
         oc8051_ram_top1_oc8051_idata_n3965,
         oc8051_ram_top1_oc8051_idata_n3964,
         oc8051_ram_top1_oc8051_idata_n3963,
         oc8051_ram_top1_oc8051_idata_n3962,
         oc8051_ram_top1_oc8051_idata_n3961,
         oc8051_ram_top1_oc8051_idata_n3960,
         oc8051_ram_top1_oc8051_idata_n3959,
         oc8051_ram_top1_oc8051_idata_n3958,
         oc8051_ram_top1_oc8051_idata_n3957,
         oc8051_ram_top1_oc8051_idata_n3956,
         oc8051_ram_top1_oc8051_idata_n3955,
         oc8051_ram_top1_oc8051_idata_n3954,
         oc8051_ram_top1_oc8051_idata_n3953,
         oc8051_ram_top1_oc8051_idata_n3952,
         oc8051_ram_top1_oc8051_idata_n3951,
         oc8051_ram_top1_oc8051_idata_n3950,
         oc8051_ram_top1_oc8051_idata_n3949,
         oc8051_ram_top1_oc8051_idata_n3948,
         oc8051_ram_top1_oc8051_idata_n3947,
         oc8051_ram_top1_oc8051_idata_n3946,
         oc8051_ram_top1_oc8051_idata_n3945,
         oc8051_ram_top1_oc8051_idata_n3944,
         oc8051_ram_top1_oc8051_idata_n3943,
         oc8051_ram_top1_oc8051_idata_n3942,
         oc8051_ram_top1_oc8051_idata_n3941,
         oc8051_ram_top1_oc8051_idata_n3940,
         oc8051_ram_top1_oc8051_idata_n3939,
         oc8051_ram_top1_oc8051_idata_n3938,
         oc8051_ram_top1_oc8051_idata_n3937,
         oc8051_ram_top1_oc8051_idata_n3936,
         oc8051_ram_top1_oc8051_idata_n3935,
         oc8051_ram_top1_oc8051_idata_n3934,
         oc8051_ram_top1_oc8051_idata_n3933,
         oc8051_ram_top1_oc8051_idata_n3932,
         oc8051_ram_top1_oc8051_idata_n3931,
         oc8051_ram_top1_oc8051_idata_n3930,
         oc8051_ram_top1_oc8051_idata_n3929,
         oc8051_ram_top1_oc8051_idata_n3928,
         oc8051_ram_top1_oc8051_idata_n3927,
         oc8051_ram_top1_oc8051_idata_n3926,
         oc8051_ram_top1_oc8051_idata_n3925,
         oc8051_ram_top1_oc8051_idata_n3924,
         oc8051_ram_top1_oc8051_idata_n3923,
         oc8051_ram_top1_oc8051_idata_n3922,
         oc8051_ram_top1_oc8051_idata_n3921,
         oc8051_ram_top1_oc8051_idata_n3920,
         oc8051_ram_top1_oc8051_idata_n3919,
         oc8051_ram_top1_oc8051_idata_n3918,
         oc8051_ram_top1_oc8051_idata_n3917,
         oc8051_ram_top1_oc8051_idata_n3916,
         oc8051_ram_top1_oc8051_idata_n3915,
         oc8051_ram_top1_oc8051_idata_n3914,
         oc8051_ram_top1_oc8051_idata_n3913,
         oc8051_ram_top1_oc8051_idata_n3912,
         oc8051_ram_top1_oc8051_idata_n3911,
         oc8051_ram_top1_oc8051_idata_n3910,
         oc8051_ram_top1_oc8051_idata_n3909,
         oc8051_ram_top1_oc8051_idata_n3908,
         oc8051_ram_top1_oc8051_idata_n3907,
         oc8051_ram_top1_oc8051_idata_n3906,
         oc8051_ram_top1_oc8051_idata_n3905,
         oc8051_ram_top1_oc8051_idata_n3904,
         oc8051_ram_top1_oc8051_idata_n3903,
         oc8051_ram_top1_oc8051_idata_n3902,
         oc8051_ram_top1_oc8051_idata_n3901,
         oc8051_ram_top1_oc8051_idata_n3900,
         oc8051_ram_top1_oc8051_idata_n3899,
         oc8051_ram_top1_oc8051_idata_n3898,
         oc8051_ram_top1_oc8051_idata_n3897,
         oc8051_ram_top1_oc8051_idata_n3896,
         oc8051_ram_top1_oc8051_idata_n3895,
         oc8051_ram_top1_oc8051_idata_n3894,
         oc8051_ram_top1_oc8051_idata_n3893,
         oc8051_ram_top1_oc8051_idata_n3892,
         oc8051_ram_top1_oc8051_idata_n3891,
         oc8051_ram_top1_oc8051_idata_n3890,
         oc8051_ram_top1_oc8051_idata_n3889,
         oc8051_ram_top1_oc8051_idata_n3888,
         oc8051_ram_top1_oc8051_idata_n3887,
         oc8051_ram_top1_oc8051_idata_n3886,
         oc8051_ram_top1_oc8051_idata_n3885,
         oc8051_ram_top1_oc8051_idata_n3884,
         oc8051_ram_top1_oc8051_idata_n3883,
         oc8051_ram_top1_oc8051_idata_n3882,
         oc8051_ram_top1_oc8051_idata_n3881,
         oc8051_ram_top1_oc8051_idata_n3880,
         oc8051_ram_top1_oc8051_idata_n3879,
         oc8051_ram_top1_oc8051_idata_n3878,
         oc8051_ram_top1_oc8051_idata_n3877,
         oc8051_ram_top1_oc8051_idata_n3876,
         oc8051_ram_top1_oc8051_idata_n3875,
         oc8051_ram_top1_oc8051_idata_n3874,
         oc8051_ram_top1_oc8051_idata_n3873,
         oc8051_ram_top1_oc8051_idata_n3872,
         oc8051_ram_top1_oc8051_idata_n3871,
         oc8051_ram_top1_oc8051_idata_n3870,
         oc8051_ram_top1_oc8051_idata_n3869,
         oc8051_ram_top1_oc8051_idata_n3868,
         oc8051_ram_top1_oc8051_idata_n3867,
         oc8051_ram_top1_oc8051_idata_n3866,
         oc8051_ram_top1_oc8051_idata_n3865,
         oc8051_ram_top1_oc8051_idata_n3864,
         oc8051_ram_top1_oc8051_idata_n3863,
         oc8051_ram_top1_oc8051_idata_n3862,
         oc8051_ram_top1_oc8051_idata_n3861,
         oc8051_ram_top1_oc8051_idata_n3860,
         oc8051_ram_top1_oc8051_idata_n3859,
         oc8051_ram_top1_oc8051_idata_n3858,
         oc8051_ram_top1_oc8051_idata_n3857,
         oc8051_ram_top1_oc8051_idata_n3856,
         oc8051_ram_top1_oc8051_idata_n3855,
         oc8051_ram_top1_oc8051_idata_n3854,
         oc8051_ram_top1_oc8051_idata_n3853,
         oc8051_ram_top1_oc8051_idata_n3852,
         oc8051_ram_top1_oc8051_idata_n3851,
         oc8051_ram_top1_oc8051_idata_n3850,
         oc8051_ram_top1_oc8051_idata_n3849,
         oc8051_ram_top1_oc8051_idata_n3848,
         oc8051_ram_top1_oc8051_idata_n3847,
         oc8051_ram_top1_oc8051_idata_n3846,
         oc8051_ram_top1_oc8051_idata_n3845,
         oc8051_ram_top1_oc8051_idata_n3844,
         oc8051_ram_top1_oc8051_idata_n3843,
         oc8051_ram_top1_oc8051_idata_n3842,
         oc8051_ram_top1_oc8051_idata_n3841,
         oc8051_ram_top1_oc8051_idata_n3840,
         oc8051_ram_top1_oc8051_idata_n3839,
         oc8051_ram_top1_oc8051_idata_n3838,
         oc8051_ram_top1_oc8051_idata_n3837,
         oc8051_ram_top1_oc8051_idata_n3836,
         oc8051_ram_top1_oc8051_idata_n3835,
         oc8051_ram_top1_oc8051_idata_n3834,
         oc8051_ram_top1_oc8051_idata_n3833,
         oc8051_ram_top1_oc8051_idata_n3832,
         oc8051_ram_top1_oc8051_idata_n3831,
         oc8051_ram_top1_oc8051_idata_n3830,
         oc8051_ram_top1_oc8051_idata_n3829,
         oc8051_ram_top1_oc8051_idata_n3828,
         oc8051_ram_top1_oc8051_idata_n3827,
         oc8051_ram_top1_oc8051_idata_n3826,
         oc8051_ram_top1_oc8051_idata_n3825,
         oc8051_ram_top1_oc8051_idata_n3824,
         oc8051_ram_top1_oc8051_idata_n3823,
         oc8051_ram_top1_oc8051_idata_n3822,
         oc8051_ram_top1_oc8051_idata_n3821,
         oc8051_ram_top1_oc8051_idata_n3820,
         oc8051_ram_top1_oc8051_idata_n3819,
         oc8051_ram_top1_oc8051_idata_n3818,
         oc8051_ram_top1_oc8051_idata_n3817,
         oc8051_ram_top1_oc8051_idata_n3816,
         oc8051_ram_top1_oc8051_idata_n3815,
         oc8051_ram_top1_oc8051_idata_n3814,
         oc8051_ram_top1_oc8051_idata_n3813,
         oc8051_ram_top1_oc8051_idata_n3812,
         oc8051_ram_top1_oc8051_idata_n3811,
         oc8051_ram_top1_oc8051_idata_n3810,
         oc8051_ram_top1_oc8051_idata_n3809,
         oc8051_ram_top1_oc8051_idata_n3808,
         oc8051_ram_top1_oc8051_idata_n3807,
         oc8051_ram_top1_oc8051_idata_n3806,
         oc8051_ram_top1_oc8051_idata_n3805,
         oc8051_ram_top1_oc8051_idata_n3804,
         oc8051_ram_top1_oc8051_idata_n3803,
         oc8051_ram_top1_oc8051_idata_n3802,
         oc8051_ram_top1_oc8051_idata_n3801,
         oc8051_ram_top1_oc8051_idata_n3800,
         oc8051_ram_top1_oc8051_idata_n3799,
         oc8051_ram_top1_oc8051_idata_n3798,
         oc8051_ram_top1_oc8051_idata_n3797,
         oc8051_ram_top1_oc8051_idata_n3796,
         oc8051_ram_top1_oc8051_idata_n3795,
         oc8051_ram_top1_oc8051_idata_n3794,
         oc8051_ram_top1_oc8051_idata_n3793,
         oc8051_ram_top1_oc8051_idata_n3792,
         oc8051_ram_top1_oc8051_idata_n3791,
         oc8051_ram_top1_oc8051_idata_n3790,
         oc8051_ram_top1_oc8051_idata_n3789,
         oc8051_ram_top1_oc8051_idata_n3788,
         oc8051_ram_top1_oc8051_idata_n3787,
         oc8051_ram_top1_oc8051_idata_n3786,
         oc8051_ram_top1_oc8051_idata_n3785,
         oc8051_ram_top1_oc8051_idata_n3784,
         oc8051_ram_top1_oc8051_idata_n3783,
         oc8051_ram_top1_oc8051_idata_n3782,
         oc8051_ram_top1_oc8051_idata_n3781,
         oc8051_ram_top1_oc8051_idata_n3780,
         oc8051_ram_top1_oc8051_idata_n3779,
         oc8051_ram_top1_oc8051_idata_n3778,
         oc8051_ram_top1_oc8051_idata_n3777,
         oc8051_ram_top1_oc8051_idata_n3776,
         oc8051_ram_top1_oc8051_idata_n3775,
         oc8051_ram_top1_oc8051_idata_n3774,
         oc8051_ram_top1_oc8051_idata_n3773,
         oc8051_ram_top1_oc8051_idata_n3772,
         oc8051_ram_top1_oc8051_idata_n3771,
         oc8051_ram_top1_oc8051_idata_n3770,
         oc8051_ram_top1_oc8051_idata_n3769,
         oc8051_ram_top1_oc8051_idata_n3768,
         oc8051_ram_top1_oc8051_idata_n3767,
         oc8051_ram_top1_oc8051_idata_n3766,
         oc8051_ram_top1_oc8051_idata_n3765,
         oc8051_ram_top1_oc8051_idata_n3764,
         oc8051_ram_top1_oc8051_idata_n3763,
         oc8051_ram_top1_oc8051_idata_n3762,
         oc8051_ram_top1_oc8051_idata_n3761,
         oc8051_ram_top1_oc8051_idata_n3760,
         oc8051_ram_top1_oc8051_idata_n3759,
         oc8051_ram_top1_oc8051_idata_n3758,
         oc8051_ram_top1_oc8051_idata_n3757,
         oc8051_ram_top1_oc8051_idata_n3756,
         oc8051_ram_top1_oc8051_idata_n3755,
         oc8051_ram_top1_oc8051_idata_n3754,
         oc8051_ram_top1_oc8051_idata_n3753,
         oc8051_ram_top1_oc8051_idata_n3752,
         oc8051_ram_top1_oc8051_idata_n3751,
         oc8051_ram_top1_oc8051_idata_n3750,
         oc8051_ram_top1_oc8051_idata_n3749,
         oc8051_ram_top1_oc8051_idata_n3748,
         oc8051_ram_top1_oc8051_idata_n3747,
         oc8051_ram_top1_oc8051_idata_n3746,
         oc8051_ram_top1_oc8051_idata_n3745,
         oc8051_ram_top1_oc8051_idata_n3744,
         oc8051_ram_top1_oc8051_idata_n3743,
         oc8051_ram_top1_oc8051_idata_n3742,
         oc8051_ram_top1_oc8051_idata_n3741,
         oc8051_ram_top1_oc8051_idata_n3740,
         oc8051_ram_top1_oc8051_idata_n3739,
         oc8051_ram_top1_oc8051_idata_n3738,
         oc8051_ram_top1_oc8051_idata_n3737,
         oc8051_ram_top1_oc8051_idata_n3736,
         oc8051_ram_top1_oc8051_idata_n3735,
         oc8051_ram_top1_oc8051_idata_n3734,
         oc8051_ram_top1_oc8051_idata_n3733,
         oc8051_ram_top1_oc8051_idata_n3732,
         oc8051_ram_top1_oc8051_idata_n3731,
         oc8051_ram_top1_oc8051_idata_n3730,
         oc8051_ram_top1_oc8051_idata_n3729,
         oc8051_ram_top1_oc8051_idata_n3728,
         oc8051_ram_top1_oc8051_idata_n3727,
         oc8051_ram_top1_oc8051_idata_n3726,
         oc8051_ram_top1_oc8051_idata_n3725,
         oc8051_ram_top1_oc8051_idata_n3724,
         oc8051_ram_top1_oc8051_idata_n3723,
         oc8051_ram_top1_oc8051_idata_n3722,
         oc8051_ram_top1_oc8051_idata_n3721,
         oc8051_ram_top1_oc8051_idata_n3720,
         oc8051_ram_top1_oc8051_idata_n3719,
         oc8051_ram_top1_oc8051_idata_n3718,
         oc8051_ram_top1_oc8051_idata_n3717,
         oc8051_ram_top1_oc8051_idata_n3716,
         oc8051_ram_top1_oc8051_idata_n3715,
         oc8051_ram_top1_oc8051_idata_n3714,
         oc8051_ram_top1_oc8051_idata_n3713,
         oc8051_ram_top1_oc8051_idata_n3712,
         oc8051_ram_top1_oc8051_idata_n3711,
         oc8051_ram_top1_oc8051_idata_n3710,
         oc8051_ram_top1_oc8051_idata_n3709,
         oc8051_ram_top1_oc8051_idata_n3708,
         oc8051_ram_top1_oc8051_idata_n3707,
         oc8051_ram_top1_oc8051_idata_n3706,
         oc8051_ram_top1_oc8051_idata_n3705,
         oc8051_ram_top1_oc8051_idata_n3704,
         oc8051_ram_top1_oc8051_idata_n3703,
         oc8051_ram_top1_oc8051_idata_n3702,
         oc8051_ram_top1_oc8051_idata_n3701,
         oc8051_ram_top1_oc8051_idata_n3700,
         oc8051_ram_top1_oc8051_idata_n3699,
         oc8051_ram_top1_oc8051_idata_n3698,
         oc8051_ram_top1_oc8051_idata_n3697,
         oc8051_ram_top1_oc8051_idata_n3696,
         oc8051_ram_top1_oc8051_idata_n3695,
         oc8051_ram_top1_oc8051_idata_n3694,
         oc8051_ram_top1_oc8051_idata_n3693,
         oc8051_ram_top1_oc8051_idata_n3692,
         oc8051_ram_top1_oc8051_idata_n3691,
         oc8051_ram_top1_oc8051_idata_n3690,
         oc8051_ram_top1_oc8051_idata_n3689,
         oc8051_ram_top1_oc8051_idata_n3688,
         oc8051_ram_top1_oc8051_idata_n3687,
         oc8051_ram_top1_oc8051_idata_n3686,
         oc8051_ram_top1_oc8051_idata_n3685,
         oc8051_ram_top1_oc8051_idata_n3684,
         oc8051_ram_top1_oc8051_idata_n3683,
         oc8051_ram_top1_oc8051_idata_n3682,
         oc8051_ram_top1_oc8051_idata_n3681,
         oc8051_ram_top1_oc8051_idata_n3680,
         oc8051_ram_top1_oc8051_idata_n3679,
         oc8051_ram_top1_oc8051_idata_n3678,
         oc8051_ram_top1_oc8051_idata_n3677,
         oc8051_ram_top1_oc8051_idata_n3676,
         oc8051_ram_top1_oc8051_idata_n3675,
         oc8051_ram_top1_oc8051_idata_n3674,
         oc8051_ram_top1_oc8051_idata_n3673,
         oc8051_ram_top1_oc8051_idata_n3672,
         oc8051_ram_top1_oc8051_idata_n3671,
         oc8051_ram_top1_oc8051_idata_n3670,
         oc8051_ram_top1_oc8051_idata_n3669,
         oc8051_ram_top1_oc8051_idata_n3668,
         oc8051_ram_top1_oc8051_idata_n3667,
         oc8051_ram_top1_oc8051_idata_n3666,
         oc8051_ram_top1_oc8051_idata_n3665,
         oc8051_ram_top1_oc8051_idata_n3664,
         oc8051_ram_top1_oc8051_idata_n3663,
         oc8051_ram_top1_oc8051_idata_n3662,
         oc8051_ram_top1_oc8051_idata_n3661,
         oc8051_ram_top1_oc8051_idata_n3660,
         oc8051_ram_top1_oc8051_idata_n3659,
         oc8051_ram_top1_oc8051_idata_n3658,
         oc8051_ram_top1_oc8051_idata_n3657,
         oc8051_ram_top1_oc8051_idata_n3656,
         oc8051_ram_top1_oc8051_idata_n3655,
         oc8051_ram_top1_oc8051_idata_n3654,
         oc8051_ram_top1_oc8051_idata_n3653,
         oc8051_ram_top1_oc8051_idata_n3652,
         oc8051_ram_top1_oc8051_idata_n3651,
         oc8051_ram_top1_oc8051_idata_n3650,
         oc8051_ram_top1_oc8051_idata_n3649,
         oc8051_ram_top1_oc8051_idata_n3648,
         oc8051_ram_top1_oc8051_idata_n3647,
         oc8051_ram_top1_oc8051_idata_n3646,
         oc8051_ram_top1_oc8051_idata_n3645,
         oc8051_ram_top1_oc8051_idata_n3644,
         oc8051_ram_top1_oc8051_idata_n3643,
         oc8051_ram_top1_oc8051_idata_n3642,
         oc8051_ram_top1_oc8051_idata_n3641,
         oc8051_ram_top1_oc8051_idata_n3640,
         oc8051_ram_top1_oc8051_idata_n3639,
         oc8051_ram_top1_oc8051_idata_n3638,
         oc8051_ram_top1_oc8051_idata_n3637,
         oc8051_ram_top1_oc8051_idata_n3636,
         oc8051_ram_top1_oc8051_idata_n3635,
         oc8051_ram_top1_oc8051_idata_n3634,
         oc8051_ram_top1_oc8051_idata_n3633,
         oc8051_ram_top1_oc8051_idata_n3632,
         oc8051_ram_top1_oc8051_idata_n3631,
         oc8051_ram_top1_oc8051_idata_n3630,
         oc8051_ram_top1_oc8051_idata_n3629,
         oc8051_ram_top1_oc8051_idata_n3628,
         oc8051_ram_top1_oc8051_idata_n3627,
         oc8051_ram_top1_oc8051_idata_n3626,
         oc8051_ram_top1_oc8051_idata_n3625,
         oc8051_ram_top1_oc8051_idata_n3624,
         oc8051_ram_top1_oc8051_idata_n3623,
         oc8051_ram_top1_oc8051_idata_n3622,
         oc8051_ram_top1_oc8051_idata_n3621,
         oc8051_ram_top1_oc8051_idata_n3620,
         oc8051_ram_top1_oc8051_idata_n3619,
         oc8051_ram_top1_oc8051_idata_n3618,
         oc8051_ram_top1_oc8051_idata_n3617,
         oc8051_ram_top1_oc8051_idata_n3616,
         oc8051_ram_top1_oc8051_idata_n3615,
         oc8051_ram_top1_oc8051_idata_n3614,
         oc8051_ram_top1_oc8051_idata_n3613,
         oc8051_ram_top1_oc8051_idata_n3612,
         oc8051_ram_top1_oc8051_idata_n3611,
         oc8051_ram_top1_oc8051_idata_n3610,
         oc8051_ram_top1_oc8051_idata_n3609,
         oc8051_ram_top1_oc8051_idata_n3608,
         oc8051_ram_top1_oc8051_idata_n3607,
         oc8051_ram_top1_oc8051_idata_n3606,
         oc8051_ram_top1_oc8051_idata_n3605,
         oc8051_ram_top1_oc8051_idata_n3604,
         oc8051_ram_top1_oc8051_idata_n3603,
         oc8051_ram_top1_oc8051_idata_n3602,
         oc8051_ram_top1_oc8051_idata_n3601,
         oc8051_ram_top1_oc8051_idata_n3600,
         oc8051_ram_top1_oc8051_idata_n3599,
         oc8051_ram_top1_oc8051_idata_n3598,
         oc8051_ram_top1_oc8051_idata_n3597,
         oc8051_ram_top1_oc8051_idata_n3596,
         oc8051_ram_top1_oc8051_idata_n3595,
         oc8051_ram_top1_oc8051_idata_n3594,
         oc8051_ram_top1_oc8051_idata_n3593,
         oc8051_ram_top1_oc8051_idata_n3592,
         oc8051_ram_top1_oc8051_idata_n3591,
         oc8051_ram_top1_oc8051_idata_n3590,
         oc8051_ram_top1_oc8051_idata_n3589,
         oc8051_ram_top1_oc8051_idata_n3588,
         oc8051_ram_top1_oc8051_idata_n3587,
         oc8051_ram_top1_oc8051_idata_n3586,
         oc8051_ram_top1_oc8051_idata_n3585,
         oc8051_ram_top1_oc8051_idata_n3584,
         oc8051_ram_top1_oc8051_idata_n3583,
         oc8051_ram_top1_oc8051_idata_n3582,
         oc8051_ram_top1_oc8051_idata_n3581,
         oc8051_ram_top1_oc8051_idata_n3580,
         oc8051_ram_top1_oc8051_idata_n3579,
         oc8051_ram_top1_oc8051_idata_n3578,
         oc8051_ram_top1_oc8051_idata_n3577,
         oc8051_ram_top1_oc8051_idata_n3576,
         oc8051_ram_top1_oc8051_idata_n3575,
         oc8051_ram_top1_oc8051_idata_n3574,
         oc8051_ram_top1_oc8051_idata_n3573,
         oc8051_ram_top1_oc8051_idata_n3572,
         oc8051_ram_top1_oc8051_idata_n3571,
         oc8051_ram_top1_oc8051_idata_n3570,
         oc8051_ram_top1_oc8051_idata_n3569,
         oc8051_ram_top1_oc8051_idata_n3568,
         oc8051_ram_top1_oc8051_idata_n3567,
         oc8051_ram_top1_oc8051_idata_n3566,
         oc8051_ram_top1_oc8051_idata_n3565,
         oc8051_ram_top1_oc8051_idata_n3564,
         oc8051_ram_top1_oc8051_idata_n3563,
         oc8051_ram_top1_oc8051_idata_n3562,
         oc8051_ram_top1_oc8051_idata_n3561,
         oc8051_ram_top1_oc8051_idata_n3560,
         oc8051_ram_top1_oc8051_idata_n3559,
         oc8051_ram_top1_oc8051_idata_n3558,
         oc8051_ram_top1_oc8051_idata_n3557,
         oc8051_ram_top1_oc8051_idata_n3556,
         oc8051_ram_top1_oc8051_idata_n3555,
         oc8051_ram_top1_oc8051_idata_n3554,
         oc8051_ram_top1_oc8051_idata_n3553,
         oc8051_ram_top1_oc8051_idata_n3552,
         oc8051_ram_top1_oc8051_idata_n3551,
         oc8051_ram_top1_oc8051_idata_n3550,
         oc8051_ram_top1_oc8051_idata_n3549,
         oc8051_ram_top1_oc8051_idata_n3548,
         oc8051_ram_top1_oc8051_idata_n3547,
         oc8051_ram_top1_oc8051_idata_n3546,
         oc8051_ram_top1_oc8051_idata_n3545,
         oc8051_ram_top1_oc8051_idata_n3544,
         oc8051_ram_top1_oc8051_idata_n3543,
         oc8051_ram_top1_oc8051_idata_n3542,
         oc8051_ram_top1_oc8051_idata_n3541,
         oc8051_ram_top1_oc8051_idata_n3540,
         oc8051_ram_top1_oc8051_idata_n3539,
         oc8051_ram_top1_oc8051_idata_n3538,
         oc8051_ram_top1_oc8051_idata_n3537,
         oc8051_ram_top1_oc8051_idata_n3536,
         oc8051_ram_top1_oc8051_idata_n3535,
         oc8051_ram_top1_oc8051_idata_n3534,
         oc8051_ram_top1_oc8051_idata_n3533,
         oc8051_ram_top1_oc8051_idata_n3532,
         oc8051_ram_top1_oc8051_idata_n3531,
         oc8051_ram_top1_oc8051_idata_n3530,
         oc8051_ram_top1_oc8051_idata_n3529,
         oc8051_ram_top1_oc8051_idata_n3528,
         oc8051_ram_top1_oc8051_idata_n3527,
         oc8051_ram_top1_oc8051_idata_n3526,
         oc8051_ram_top1_oc8051_idata_n3525,
         oc8051_ram_top1_oc8051_idata_n3524,
         oc8051_ram_top1_oc8051_idata_n3523,
         oc8051_ram_top1_oc8051_idata_n3522,
         oc8051_ram_top1_oc8051_idata_n3521,
         oc8051_ram_top1_oc8051_idata_n3520,
         oc8051_ram_top1_oc8051_idata_n3519,
         oc8051_ram_top1_oc8051_idata_n3518,
         oc8051_ram_top1_oc8051_idata_n3517,
         oc8051_ram_top1_oc8051_idata_n3516,
         oc8051_ram_top1_oc8051_idata_n3515,
         oc8051_ram_top1_oc8051_idata_n3514,
         oc8051_ram_top1_oc8051_idata_n3513,
         oc8051_ram_top1_oc8051_idata_n3512,
         oc8051_ram_top1_oc8051_idata_n3511,
         oc8051_ram_top1_oc8051_idata_n3510,
         oc8051_ram_top1_oc8051_idata_n3509,
         oc8051_ram_top1_oc8051_idata_n3508,
         oc8051_ram_top1_oc8051_idata_n3507,
         oc8051_ram_top1_oc8051_idata_n3506,
         oc8051_ram_top1_oc8051_idata_n3505,
         oc8051_ram_top1_oc8051_idata_n3504,
         oc8051_ram_top1_oc8051_idata_n3503,
         oc8051_ram_top1_oc8051_idata_n3502,
         oc8051_ram_top1_oc8051_idata_n3501,
         oc8051_ram_top1_oc8051_idata_n3500,
         oc8051_ram_top1_oc8051_idata_n3499,
         oc8051_ram_top1_oc8051_idata_n3498,
         oc8051_ram_top1_oc8051_idata_n3497,
         oc8051_ram_top1_oc8051_idata_n3496,
         oc8051_ram_top1_oc8051_idata_n3495,
         oc8051_ram_top1_oc8051_idata_n3494,
         oc8051_ram_top1_oc8051_idata_n3493,
         oc8051_ram_top1_oc8051_idata_n3492,
         oc8051_ram_top1_oc8051_idata_n3491,
         oc8051_ram_top1_oc8051_idata_n3490,
         oc8051_ram_top1_oc8051_idata_n3489,
         oc8051_ram_top1_oc8051_idata_n3488,
         oc8051_ram_top1_oc8051_idata_n3487,
         oc8051_ram_top1_oc8051_idata_n3486,
         oc8051_ram_top1_oc8051_idata_n3485,
         oc8051_ram_top1_oc8051_idata_n3484,
         oc8051_ram_top1_oc8051_idata_n3483,
         oc8051_ram_top1_oc8051_idata_n3482,
         oc8051_ram_top1_oc8051_idata_n3481,
         oc8051_ram_top1_oc8051_idata_n3480,
         oc8051_ram_top1_oc8051_idata_n3479,
         oc8051_ram_top1_oc8051_idata_n3478,
         oc8051_ram_top1_oc8051_idata_n3477,
         oc8051_ram_top1_oc8051_idata_n3476,
         oc8051_ram_top1_oc8051_idata_n3475,
         oc8051_ram_top1_oc8051_idata_n3474,
         oc8051_ram_top1_oc8051_idata_n3473,
         oc8051_ram_top1_oc8051_idata_n3472,
         oc8051_ram_top1_oc8051_idata_n3471,
         oc8051_ram_top1_oc8051_idata_n3470,
         oc8051_ram_top1_oc8051_idata_n3469,
         oc8051_ram_top1_oc8051_idata_n3468,
         oc8051_ram_top1_oc8051_idata_n3467,
         oc8051_ram_top1_oc8051_idata_n3466,
         oc8051_ram_top1_oc8051_idata_n3465,
         oc8051_ram_top1_oc8051_idata_n3464,
         oc8051_ram_top1_oc8051_idata_n3463,
         oc8051_ram_top1_oc8051_idata_n3462,
         oc8051_ram_top1_oc8051_idata_n3461,
         oc8051_ram_top1_oc8051_idata_n3460,
         oc8051_ram_top1_oc8051_idata_n3459,
         oc8051_ram_top1_oc8051_idata_n3458,
         oc8051_ram_top1_oc8051_idata_n3457,
         oc8051_ram_top1_oc8051_idata_n3456,
         oc8051_ram_top1_oc8051_idata_n3455,
         oc8051_ram_top1_oc8051_idata_n3454,
         oc8051_ram_top1_oc8051_idata_n3453,
         oc8051_ram_top1_oc8051_idata_n3452,
         oc8051_ram_top1_oc8051_idata_n3451,
         oc8051_ram_top1_oc8051_idata_n3450,
         oc8051_ram_top1_oc8051_idata_n3449,
         oc8051_ram_top1_oc8051_idata_n3448,
         oc8051_ram_top1_oc8051_idata_n3447,
         oc8051_ram_top1_oc8051_idata_n3446,
         oc8051_ram_top1_oc8051_idata_n3445,
         oc8051_ram_top1_oc8051_idata_n3444,
         oc8051_ram_top1_oc8051_idata_n3443,
         oc8051_ram_top1_oc8051_idata_n3442,
         oc8051_ram_top1_oc8051_idata_n3441,
         oc8051_ram_top1_oc8051_idata_n3440,
         oc8051_ram_top1_oc8051_idata_n3439,
         oc8051_ram_top1_oc8051_idata_n3438,
         oc8051_ram_top1_oc8051_idata_n3437,
         oc8051_ram_top1_oc8051_idata_n3436,
         oc8051_ram_top1_oc8051_idata_n3435,
         oc8051_ram_top1_oc8051_idata_n3434,
         oc8051_ram_top1_oc8051_idata_n3433,
         oc8051_ram_top1_oc8051_idata_n3432,
         oc8051_ram_top1_oc8051_idata_n3431,
         oc8051_ram_top1_oc8051_idata_n3430,
         oc8051_ram_top1_oc8051_idata_n3429,
         oc8051_ram_top1_oc8051_idata_n3428,
         oc8051_ram_top1_oc8051_idata_n3427,
         oc8051_ram_top1_oc8051_idata_n3426,
         oc8051_ram_top1_oc8051_idata_n3425,
         oc8051_ram_top1_oc8051_idata_n3424,
         oc8051_ram_top1_oc8051_idata_n3423,
         oc8051_ram_top1_oc8051_idata_n3422,
         oc8051_ram_top1_oc8051_idata_n3421,
         oc8051_ram_top1_oc8051_idata_n3420,
         oc8051_ram_top1_oc8051_idata_n3419,
         oc8051_ram_top1_oc8051_idata_n3418,
         oc8051_ram_top1_oc8051_idata_n3417,
         oc8051_ram_top1_oc8051_idata_n3416,
         oc8051_ram_top1_oc8051_idata_n3415,
         oc8051_ram_top1_oc8051_idata_n3414,
         oc8051_ram_top1_oc8051_idata_n3413,
         oc8051_ram_top1_oc8051_idata_n3412,
         oc8051_ram_top1_oc8051_idata_n3411,
         oc8051_ram_top1_oc8051_idata_n3410,
         oc8051_ram_top1_oc8051_idata_n3409,
         oc8051_ram_top1_oc8051_idata_n3408,
         oc8051_ram_top1_oc8051_idata_n3407,
         oc8051_ram_top1_oc8051_idata_n3406,
         oc8051_ram_top1_oc8051_idata_n3405,
         oc8051_ram_top1_oc8051_idata_n3404,
         oc8051_ram_top1_oc8051_idata_n3403,
         oc8051_ram_top1_oc8051_idata_n3402,
         oc8051_ram_top1_oc8051_idata_n3401,
         oc8051_ram_top1_oc8051_idata_n3400,
         oc8051_ram_top1_oc8051_idata_n3399,
         oc8051_ram_top1_oc8051_idata_n3398,
         oc8051_ram_top1_oc8051_idata_n3397,
         oc8051_ram_top1_oc8051_idata_n3396,
         oc8051_ram_top1_oc8051_idata_n3395,
         oc8051_ram_top1_oc8051_idata_n3394,
         oc8051_ram_top1_oc8051_idata_n3393,
         oc8051_ram_top1_oc8051_idata_n3392,
         oc8051_ram_top1_oc8051_idata_n3391,
         oc8051_ram_top1_oc8051_idata_n3390,
         oc8051_ram_top1_oc8051_idata_n3389,
         oc8051_ram_top1_oc8051_idata_n3388,
         oc8051_ram_top1_oc8051_idata_n3387,
         oc8051_ram_top1_oc8051_idata_n3386,
         oc8051_ram_top1_oc8051_idata_n3385,
         oc8051_ram_top1_oc8051_idata_n3384,
         oc8051_ram_top1_oc8051_idata_n3383,
         oc8051_ram_top1_oc8051_idata_n3382,
         oc8051_ram_top1_oc8051_idata_n3381,
         oc8051_ram_top1_oc8051_idata_n3380,
         oc8051_ram_top1_oc8051_idata_n3379,
         oc8051_ram_top1_oc8051_idata_n3378,
         oc8051_ram_top1_oc8051_idata_n3377,
         oc8051_ram_top1_oc8051_idata_n3376,
         oc8051_ram_top1_oc8051_idata_n3375,
         oc8051_ram_top1_oc8051_idata_n3374,
         oc8051_ram_top1_oc8051_idata_n3373,
         oc8051_ram_top1_oc8051_idata_n3372,
         oc8051_ram_top1_oc8051_idata_n3371,
         oc8051_ram_top1_oc8051_idata_n3370,
         oc8051_ram_top1_oc8051_idata_n3369,
         oc8051_ram_top1_oc8051_idata_n3368,
         oc8051_ram_top1_oc8051_idata_n3367,
         oc8051_ram_top1_oc8051_idata_n3366,
         oc8051_ram_top1_oc8051_idata_n3365,
         oc8051_ram_top1_oc8051_idata_n3364,
         oc8051_ram_top1_oc8051_idata_n3363,
         oc8051_ram_top1_oc8051_idata_n3362,
         oc8051_ram_top1_oc8051_idata_n3361,
         oc8051_ram_top1_oc8051_idata_n3360,
         oc8051_ram_top1_oc8051_idata_n3359,
         oc8051_ram_top1_oc8051_idata_n3358,
         oc8051_ram_top1_oc8051_idata_n3357,
         oc8051_ram_top1_oc8051_idata_n3356,
         oc8051_ram_top1_oc8051_idata_n3355,
         oc8051_ram_top1_oc8051_idata_n3354,
         oc8051_ram_top1_oc8051_idata_n3353,
         oc8051_ram_top1_oc8051_idata_n3352,
         oc8051_ram_top1_oc8051_idata_n3351,
         oc8051_ram_top1_oc8051_idata_n3350,
         oc8051_ram_top1_oc8051_idata_n3349,
         oc8051_ram_top1_oc8051_idata_n3348,
         oc8051_ram_top1_oc8051_idata_n3347,
         oc8051_ram_top1_oc8051_idata_n3346,
         oc8051_ram_top1_oc8051_idata_n3345,
         oc8051_ram_top1_oc8051_idata_n3344,
         oc8051_ram_top1_oc8051_idata_n3343,
         oc8051_ram_top1_oc8051_idata_n3342,
         oc8051_ram_top1_oc8051_idata_n3341,
         oc8051_ram_top1_oc8051_idata_n3340,
         oc8051_ram_top1_oc8051_idata_n3339,
         oc8051_ram_top1_oc8051_idata_n3338,
         oc8051_ram_top1_oc8051_idata_n3337,
         oc8051_ram_top1_oc8051_idata_n3336,
         oc8051_ram_top1_oc8051_idata_n3335,
         oc8051_ram_top1_oc8051_idata_n3334,
         oc8051_ram_top1_oc8051_idata_n3333,
         oc8051_ram_top1_oc8051_idata_n3332,
         oc8051_ram_top1_oc8051_idata_n3331,
         oc8051_ram_top1_oc8051_idata_n3330,
         oc8051_ram_top1_oc8051_idata_n3329,
         oc8051_ram_top1_oc8051_idata_n3328,
         oc8051_ram_top1_oc8051_idata_n3327,
         oc8051_ram_top1_oc8051_idata_n3326,
         oc8051_ram_top1_oc8051_idata_n3325,
         oc8051_ram_top1_oc8051_idata_n3324,
         oc8051_ram_top1_oc8051_idata_n3323,
         oc8051_ram_top1_oc8051_idata_n3322,
         oc8051_ram_top1_oc8051_idata_n3321,
         oc8051_ram_top1_oc8051_idata_n3320,
         oc8051_ram_top1_oc8051_idata_n3319,
         oc8051_ram_top1_oc8051_idata_n3318,
         oc8051_ram_top1_oc8051_idata_n3317,
         oc8051_ram_top1_oc8051_idata_n3316,
         oc8051_ram_top1_oc8051_idata_n3315,
         oc8051_ram_top1_oc8051_idata_n3314,
         oc8051_ram_top1_oc8051_idata_n3313,
         oc8051_ram_top1_oc8051_idata_n3312,
         oc8051_ram_top1_oc8051_idata_n3311,
         oc8051_ram_top1_oc8051_idata_n3310,
         oc8051_ram_top1_oc8051_idata_n3309,
         oc8051_ram_top1_oc8051_idata_n3308,
         oc8051_ram_top1_oc8051_idata_n3307,
         oc8051_ram_top1_oc8051_idata_n3306,
         oc8051_ram_top1_oc8051_idata_n3305,
         oc8051_ram_top1_oc8051_idata_n3304,
         oc8051_ram_top1_oc8051_idata_n3303,
         oc8051_ram_top1_oc8051_idata_n3302,
         oc8051_ram_top1_oc8051_idata_n3301,
         oc8051_ram_top1_oc8051_idata_n3300,
         oc8051_ram_top1_oc8051_idata_n3299,
         oc8051_ram_top1_oc8051_idata_n3298,
         oc8051_ram_top1_oc8051_idata_n3297,
         oc8051_ram_top1_oc8051_idata_n3296,
         oc8051_ram_top1_oc8051_idata_n3295,
         oc8051_ram_top1_oc8051_idata_n3294,
         oc8051_ram_top1_oc8051_idata_n3293,
         oc8051_ram_top1_oc8051_idata_n3292,
         oc8051_ram_top1_oc8051_idata_n3291,
         oc8051_ram_top1_oc8051_idata_n3290,
         oc8051_ram_top1_oc8051_idata_n3289,
         oc8051_ram_top1_oc8051_idata_n3288,
         oc8051_ram_top1_oc8051_idata_n3287,
         oc8051_ram_top1_oc8051_idata_n3286,
         oc8051_ram_top1_oc8051_idata_n3285,
         oc8051_ram_top1_oc8051_idata_n3284,
         oc8051_ram_top1_oc8051_idata_n3283,
         oc8051_ram_top1_oc8051_idata_n3282,
         oc8051_ram_top1_oc8051_idata_n3281,
         oc8051_ram_top1_oc8051_idata_n3280,
         oc8051_ram_top1_oc8051_idata_n3279,
         oc8051_ram_top1_oc8051_idata_n3278,
         oc8051_ram_top1_oc8051_idata_n3277,
         oc8051_ram_top1_oc8051_idata_n3276,
         oc8051_ram_top1_oc8051_idata_n3275,
         oc8051_ram_top1_oc8051_idata_n3274,
         oc8051_ram_top1_oc8051_idata_n3273,
         oc8051_ram_top1_oc8051_idata_n3272,
         oc8051_ram_top1_oc8051_idata_n3271,
         oc8051_ram_top1_oc8051_idata_n3270,
         oc8051_ram_top1_oc8051_idata_n3269,
         oc8051_ram_top1_oc8051_idata_n3268,
         oc8051_ram_top1_oc8051_idata_n3267,
         oc8051_ram_top1_oc8051_idata_n3266,
         oc8051_ram_top1_oc8051_idata_n3265,
         oc8051_ram_top1_oc8051_idata_n3264,
         oc8051_ram_top1_oc8051_idata_n3263,
         oc8051_ram_top1_oc8051_idata_n3262,
         oc8051_ram_top1_oc8051_idata_n3261,
         oc8051_ram_top1_oc8051_idata_n3260,
         oc8051_ram_top1_oc8051_idata_n3259,
         oc8051_ram_top1_oc8051_idata_n3258,
         oc8051_ram_top1_oc8051_idata_n3257,
         oc8051_ram_top1_oc8051_idata_n3256,
         oc8051_ram_top1_oc8051_idata_n3255,
         oc8051_ram_top1_oc8051_idata_n3254,
         oc8051_ram_top1_oc8051_idata_n3253,
         oc8051_ram_top1_oc8051_idata_n3252,
         oc8051_ram_top1_oc8051_idata_n3251,
         oc8051_ram_top1_oc8051_idata_n3250,
         oc8051_ram_top1_oc8051_idata_n3249,
         oc8051_ram_top1_oc8051_idata_n3248,
         oc8051_ram_top1_oc8051_idata_n3247,
         oc8051_ram_top1_oc8051_idata_n3246,
         oc8051_ram_top1_oc8051_idata_n3245,
         oc8051_ram_top1_oc8051_idata_n3244,
         oc8051_ram_top1_oc8051_idata_n3243,
         oc8051_ram_top1_oc8051_idata_n3242,
         oc8051_ram_top1_oc8051_idata_n3241,
         oc8051_ram_top1_oc8051_idata_n3240,
         oc8051_ram_top1_oc8051_idata_n3239,
         oc8051_ram_top1_oc8051_idata_n3238,
         oc8051_ram_top1_oc8051_idata_n3237,
         oc8051_ram_top1_oc8051_idata_n3236,
         oc8051_ram_top1_oc8051_idata_n3235,
         oc8051_ram_top1_oc8051_idata_n3234,
         oc8051_ram_top1_oc8051_idata_n3233,
         oc8051_ram_top1_oc8051_idata_n3232,
         oc8051_ram_top1_oc8051_idata_n3231,
         oc8051_ram_top1_oc8051_idata_n3230,
         oc8051_ram_top1_oc8051_idata_n3229,
         oc8051_ram_top1_oc8051_idata_n3228,
         oc8051_ram_top1_oc8051_idata_n3227,
         oc8051_ram_top1_oc8051_idata_n3226,
         oc8051_ram_top1_oc8051_idata_n3225,
         oc8051_ram_top1_oc8051_idata_n3224,
         oc8051_ram_top1_oc8051_idata_n3223,
         oc8051_ram_top1_oc8051_idata_n3222,
         oc8051_ram_top1_oc8051_idata_n3221,
         oc8051_ram_top1_oc8051_idata_n3220,
         oc8051_ram_top1_oc8051_idata_n3219,
         oc8051_ram_top1_oc8051_idata_n3218,
         oc8051_ram_top1_oc8051_idata_n3217,
         oc8051_ram_top1_oc8051_idata_n3216,
         oc8051_ram_top1_oc8051_idata_n3215,
         oc8051_ram_top1_oc8051_idata_n3214,
         oc8051_ram_top1_oc8051_idata_n3213,
         oc8051_ram_top1_oc8051_idata_n3212,
         oc8051_ram_top1_oc8051_idata_n3211,
         oc8051_ram_top1_oc8051_idata_n3210,
         oc8051_ram_top1_oc8051_idata_n3209,
         oc8051_ram_top1_oc8051_idata_n3208,
         oc8051_ram_top1_oc8051_idata_n3207,
         oc8051_ram_top1_oc8051_idata_n3206,
         oc8051_ram_top1_oc8051_idata_n3205,
         oc8051_ram_top1_oc8051_idata_n3204,
         oc8051_ram_top1_oc8051_idata_n3203,
         oc8051_ram_top1_oc8051_idata_n3202,
         oc8051_ram_top1_oc8051_idata_n3201,
         oc8051_ram_top1_oc8051_idata_n3200,
         oc8051_ram_top1_oc8051_idata_n3199,
         oc8051_ram_top1_oc8051_idata_n3198,
         oc8051_ram_top1_oc8051_idata_n3197,
         oc8051_ram_top1_oc8051_idata_n3196,
         oc8051_ram_top1_oc8051_idata_n3195,
         oc8051_ram_top1_oc8051_idata_n3194,
         oc8051_ram_top1_oc8051_idata_n3193,
         oc8051_ram_top1_oc8051_idata_n3192,
         oc8051_ram_top1_oc8051_idata_n3191,
         oc8051_ram_top1_oc8051_idata_n3190,
         oc8051_ram_top1_oc8051_idata_n3189,
         oc8051_ram_top1_oc8051_idata_n3188,
         oc8051_ram_top1_oc8051_idata_n3187,
         oc8051_ram_top1_oc8051_idata_n3186,
         oc8051_ram_top1_oc8051_idata_n3185,
         oc8051_ram_top1_oc8051_idata_n3184,
         oc8051_ram_top1_oc8051_idata_n3183,
         oc8051_ram_top1_oc8051_idata_n3182,
         oc8051_ram_top1_oc8051_idata_n3181,
         oc8051_ram_top1_oc8051_idata_n3180,
         oc8051_ram_top1_oc8051_idata_n3179,
         oc8051_ram_top1_oc8051_idata_n3178,
         oc8051_ram_top1_oc8051_idata_n3177,
         oc8051_ram_top1_oc8051_idata_n3176,
         oc8051_ram_top1_oc8051_idata_n3175,
         oc8051_ram_top1_oc8051_idata_n3174,
         oc8051_ram_top1_oc8051_idata_n3173,
         oc8051_ram_top1_oc8051_idata_n3172,
         oc8051_ram_top1_oc8051_idata_n3171,
         oc8051_ram_top1_oc8051_idata_n3170,
         oc8051_ram_top1_oc8051_idata_n3169,
         oc8051_ram_top1_oc8051_idata_n3168,
         oc8051_ram_top1_oc8051_idata_n3167,
         oc8051_ram_top1_oc8051_idata_n3166,
         oc8051_ram_top1_oc8051_idata_n3165,
         oc8051_ram_top1_oc8051_idata_n3164,
         oc8051_ram_top1_oc8051_idata_n3163,
         oc8051_ram_top1_oc8051_idata_n3162,
         oc8051_ram_top1_oc8051_idata_n3161,
         oc8051_ram_top1_oc8051_idata_n3160,
         oc8051_ram_top1_oc8051_idata_n3159,
         oc8051_ram_top1_oc8051_idata_n3158,
         oc8051_ram_top1_oc8051_idata_n3157,
         oc8051_ram_top1_oc8051_idata_n3156,
         oc8051_ram_top1_oc8051_idata_n3155,
         oc8051_ram_top1_oc8051_idata_n3154,
         oc8051_ram_top1_oc8051_idata_n3153,
         oc8051_ram_top1_oc8051_idata_n3152,
         oc8051_ram_top1_oc8051_idata_n3151,
         oc8051_ram_top1_oc8051_idata_n3150,
         oc8051_ram_top1_oc8051_idata_n3149,
         oc8051_ram_top1_oc8051_idata_n3148,
         oc8051_ram_top1_oc8051_idata_n3147,
         oc8051_ram_top1_oc8051_idata_n3146,
         oc8051_ram_top1_oc8051_idata_n3145,
         oc8051_ram_top1_oc8051_idata_n3144,
         oc8051_ram_top1_oc8051_idata_n3143,
         oc8051_ram_top1_oc8051_idata_n3142,
         oc8051_ram_top1_oc8051_idata_n3141,
         oc8051_ram_top1_oc8051_idata_n3140,
         oc8051_ram_top1_oc8051_idata_n3139,
         oc8051_ram_top1_oc8051_idata_n3138,
         oc8051_ram_top1_oc8051_idata_n3137,
         oc8051_ram_top1_oc8051_idata_n3136,
         oc8051_ram_top1_oc8051_idata_n3135,
         oc8051_ram_top1_oc8051_idata_n3134,
         oc8051_ram_top1_oc8051_idata_n3133,
         oc8051_ram_top1_oc8051_idata_n3132,
         oc8051_ram_top1_oc8051_idata_n3131,
         oc8051_ram_top1_oc8051_idata_n3130,
         oc8051_ram_top1_oc8051_idata_n3129,
         oc8051_ram_top1_oc8051_idata_n3128,
         oc8051_ram_top1_oc8051_idata_n3127,
         oc8051_ram_top1_oc8051_idata_n3126,
         oc8051_ram_top1_oc8051_idata_n3125,
         oc8051_ram_top1_oc8051_idata_n3124,
         oc8051_ram_top1_oc8051_idata_n3123,
         oc8051_ram_top1_oc8051_idata_n3122,
         oc8051_ram_top1_oc8051_idata_n3121,
         oc8051_ram_top1_oc8051_idata_n3120,
         oc8051_ram_top1_oc8051_idata_n3119,
         oc8051_ram_top1_oc8051_idata_n3118,
         oc8051_ram_top1_oc8051_idata_n3117,
         oc8051_ram_top1_oc8051_idata_n3116,
         oc8051_ram_top1_oc8051_idata_n3115,
         oc8051_ram_top1_oc8051_idata_n3114,
         oc8051_ram_top1_oc8051_idata_n3113,
         oc8051_ram_top1_oc8051_idata_n3112,
         oc8051_ram_top1_oc8051_idata_n3111,
         oc8051_ram_top1_oc8051_idata_n3110,
         oc8051_ram_top1_oc8051_idata_n3109,
         oc8051_ram_top1_oc8051_idata_n3108,
         oc8051_ram_top1_oc8051_idata_n3107,
         oc8051_ram_top1_oc8051_idata_n3106,
         oc8051_ram_top1_oc8051_idata_n3105,
         oc8051_ram_top1_oc8051_idata_n3104,
         oc8051_ram_top1_oc8051_idata_n3103,
         oc8051_ram_top1_oc8051_idata_n3102,
         oc8051_ram_top1_oc8051_idata_n3101,
         oc8051_ram_top1_oc8051_idata_n3100,
         oc8051_ram_top1_oc8051_idata_n3099,
         oc8051_ram_top1_oc8051_idata_n3098,
         oc8051_ram_top1_oc8051_idata_n3097,
         oc8051_ram_top1_oc8051_idata_n3096,
         oc8051_ram_top1_oc8051_idata_n3095,
         oc8051_ram_top1_oc8051_idata_n3094,
         oc8051_ram_top1_oc8051_idata_n3093,
         oc8051_ram_top1_oc8051_idata_n3092,
         oc8051_ram_top1_oc8051_idata_n3091,
         oc8051_ram_top1_oc8051_idata_n3090,
         oc8051_ram_top1_oc8051_idata_n3089,
         oc8051_ram_top1_oc8051_idata_n3088,
         oc8051_ram_top1_oc8051_idata_n3087,
         oc8051_ram_top1_oc8051_idata_n3086,
         oc8051_ram_top1_oc8051_idata_n3085,
         oc8051_ram_top1_oc8051_idata_n3084,
         oc8051_ram_top1_oc8051_idata_n3083,
         oc8051_ram_top1_oc8051_idata_n3082,
         oc8051_ram_top1_oc8051_idata_n3081,
         oc8051_ram_top1_oc8051_idata_n3080,
         oc8051_ram_top1_oc8051_idata_n3079,
         oc8051_ram_top1_oc8051_idata_n3078,
         oc8051_ram_top1_oc8051_idata_n3077,
         oc8051_ram_top1_oc8051_idata_n3076,
         oc8051_ram_top1_oc8051_idata_n3075,
         oc8051_ram_top1_oc8051_idata_n3074,
         oc8051_ram_top1_oc8051_idata_n3073,
         oc8051_ram_top1_oc8051_idata_n3072,
         oc8051_ram_top1_oc8051_idata_n3071,
         oc8051_ram_top1_oc8051_idata_n3070,
         oc8051_ram_top1_oc8051_idata_n3069,
         oc8051_ram_top1_oc8051_idata_n3068,
         oc8051_ram_top1_oc8051_idata_n3067,
         oc8051_ram_top1_oc8051_idata_n3066,
         oc8051_ram_top1_oc8051_idata_n3065,
         oc8051_ram_top1_oc8051_idata_n3064,
         oc8051_ram_top1_oc8051_idata_n3063,
         oc8051_ram_top1_oc8051_idata_n3062,
         oc8051_ram_top1_oc8051_idata_n3061,
         oc8051_ram_top1_oc8051_idata_n3060,
         oc8051_ram_top1_oc8051_idata_n3059,
         oc8051_ram_top1_oc8051_idata_n3058,
         oc8051_ram_top1_oc8051_idata_n3057,
         oc8051_ram_top1_oc8051_idata_n3056,
         oc8051_ram_top1_oc8051_idata_n3055,
         oc8051_ram_top1_oc8051_idata_n3054,
         oc8051_ram_top1_oc8051_idata_n3053,
         oc8051_ram_top1_oc8051_idata_n3052,
         oc8051_ram_top1_oc8051_idata_n3051,
         oc8051_ram_top1_oc8051_idata_n3050,
         oc8051_ram_top1_oc8051_idata_n3049,
         oc8051_ram_top1_oc8051_idata_n3048,
         oc8051_ram_top1_oc8051_idata_n3047,
         oc8051_ram_top1_oc8051_idata_n3046,
         oc8051_ram_top1_oc8051_idata_n3045,
         oc8051_ram_top1_oc8051_idata_n3044,
         oc8051_ram_top1_oc8051_idata_n3043,
         oc8051_ram_top1_oc8051_idata_n3042,
         oc8051_ram_top1_oc8051_idata_n3041,
         oc8051_ram_top1_oc8051_idata_n3040,
         oc8051_ram_top1_oc8051_idata_n3039,
         oc8051_ram_top1_oc8051_idata_n3038,
         oc8051_ram_top1_oc8051_idata_n3037,
         oc8051_ram_top1_oc8051_idata_n3036,
         oc8051_ram_top1_oc8051_idata_n3035,
         oc8051_ram_top1_oc8051_idata_n3034,
         oc8051_ram_top1_oc8051_idata_n3033,
         oc8051_ram_top1_oc8051_idata_n3032,
         oc8051_ram_top1_oc8051_idata_n3031,
         oc8051_ram_top1_oc8051_idata_n3030,
         oc8051_ram_top1_oc8051_idata_n3029,
         oc8051_ram_top1_oc8051_idata_n3028,
         oc8051_ram_top1_oc8051_idata_n3027,
         oc8051_ram_top1_oc8051_idata_n3026,
         oc8051_ram_top1_oc8051_idata_n3025,
         oc8051_ram_top1_oc8051_idata_n3024,
         oc8051_ram_top1_oc8051_idata_n3023,
         oc8051_ram_top1_oc8051_idata_n3022,
         oc8051_ram_top1_oc8051_idata_n3021,
         oc8051_ram_top1_oc8051_idata_n3020,
         oc8051_ram_top1_oc8051_idata_n3019,
         oc8051_ram_top1_oc8051_idata_n3018,
         oc8051_ram_top1_oc8051_idata_n3017,
         oc8051_ram_top1_oc8051_idata_n3016,
         oc8051_ram_top1_oc8051_idata_n3015,
         oc8051_ram_top1_oc8051_idata_n3014,
         oc8051_ram_top1_oc8051_idata_n3013,
         oc8051_ram_top1_oc8051_idata_n3012,
         oc8051_ram_top1_oc8051_idata_n3011,
         oc8051_ram_top1_oc8051_idata_n3010,
         oc8051_ram_top1_oc8051_idata_n3009,
         oc8051_ram_top1_oc8051_idata_n3008,
         oc8051_ram_top1_oc8051_idata_n3007,
         oc8051_ram_top1_oc8051_idata_n3006,
         oc8051_ram_top1_oc8051_idata_n3005,
         oc8051_ram_top1_oc8051_idata_n3004,
         oc8051_ram_top1_oc8051_idata_n3003,
         oc8051_ram_top1_oc8051_idata_n3002,
         oc8051_ram_top1_oc8051_idata_n3001,
         oc8051_ram_top1_oc8051_idata_n3000,
         oc8051_ram_top1_oc8051_idata_n2999,
         oc8051_ram_top1_oc8051_idata_n2998,
         oc8051_ram_top1_oc8051_idata_n2997,
         oc8051_ram_top1_oc8051_idata_n2996,
         oc8051_ram_top1_oc8051_idata_n2995,
         oc8051_ram_top1_oc8051_idata_n2994,
         oc8051_ram_top1_oc8051_idata_n2993,
         oc8051_ram_top1_oc8051_idata_n2992,
         oc8051_ram_top1_oc8051_idata_n2991,
         oc8051_ram_top1_oc8051_idata_n2990,
         oc8051_ram_top1_oc8051_idata_n2989,
         oc8051_ram_top1_oc8051_idata_n2988,
         oc8051_ram_top1_oc8051_idata_n2987,
         oc8051_ram_top1_oc8051_idata_n2986,
         oc8051_ram_top1_oc8051_idata_n2985,
         oc8051_ram_top1_oc8051_idata_n2984,
         oc8051_ram_top1_oc8051_idata_n2983,
         oc8051_ram_top1_oc8051_idata_n2982,
         oc8051_ram_top1_oc8051_idata_n2981,
         oc8051_ram_top1_oc8051_idata_n2980,
         oc8051_ram_top1_oc8051_idata_n2979,
         oc8051_ram_top1_oc8051_idata_n2978,
         oc8051_ram_top1_oc8051_idata_n2977,
         oc8051_ram_top1_oc8051_idata_n2976,
         oc8051_ram_top1_oc8051_idata_n2975,
         oc8051_ram_top1_oc8051_idata_n2974,
         oc8051_ram_top1_oc8051_idata_n2973,
         oc8051_ram_top1_oc8051_idata_n2972,
         oc8051_ram_top1_oc8051_idata_n2971,
         oc8051_ram_top1_oc8051_idata_n2970,
         oc8051_ram_top1_oc8051_idata_n2969,
         oc8051_ram_top1_oc8051_idata_n2968,
         oc8051_ram_top1_oc8051_idata_n2967,
         oc8051_ram_top1_oc8051_idata_n2966,
         oc8051_ram_top1_oc8051_idata_n2965,
         oc8051_ram_top1_oc8051_idata_n2964,
         oc8051_ram_top1_oc8051_idata_n2963,
         oc8051_ram_top1_oc8051_idata_n2962,
         oc8051_ram_top1_oc8051_idata_n2961,
         oc8051_ram_top1_oc8051_idata_n2960,
         oc8051_ram_top1_oc8051_idata_n2959,
         oc8051_ram_top1_oc8051_idata_n2958,
         oc8051_ram_top1_oc8051_idata_n2957,
         oc8051_ram_top1_oc8051_idata_n2956,
         oc8051_ram_top1_oc8051_idata_n2955,
         oc8051_ram_top1_oc8051_idata_n2954,
         oc8051_ram_top1_oc8051_idata_n2953,
         oc8051_ram_top1_oc8051_idata_n2952,
         oc8051_ram_top1_oc8051_idata_n2951,
         oc8051_ram_top1_oc8051_idata_n2950,
         oc8051_ram_top1_oc8051_idata_n2949,
         oc8051_ram_top1_oc8051_idata_n2948,
         oc8051_ram_top1_oc8051_idata_n2947,
         oc8051_ram_top1_oc8051_idata_n2946,
         oc8051_ram_top1_oc8051_idata_n2945,
         oc8051_ram_top1_oc8051_idata_n2944,
         oc8051_ram_top1_oc8051_idata_n2943,
         oc8051_ram_top1_oc8051_idata_n2942,
         oc8051_ram_top1_oc8051_idata_n2941,
         oc8051_ram_top1_oc8051_idata_n2940,
         oc8051_ram_top1_oc8051_idata_n2939,
         oc8051_ram_top1_oc8051_idata_n2938,
         oc8051_ram_top1_oc8051_idata_n2937,
         oc8051_ram_top1_oc8051_idata_n2936,
         oc8051_ram_top1_oc8051_idata_n2935,
         oc8051_ram_top1_oc8051_idata_n2934,
         oc8051_ram_top1_oc8051_idata_n2933,
         oc8051_ram_top1_oc8051_idata_n2932,
         oc8051_ram_top1_oc8051_idata_n2931,
         oc8051_ram_top1_oc8051_idata_n2930,
         oc8051_ram_top1_oc8051_idata_n2929,
         oc8051_ram_top1_oc8051_idata_n2928,
         oc8051_ram_top1_oc8051_idata_n2927,
         oc8051_ram_top1_oc8051_idata_n2926,
         oc8051_ram_top1_oc8051_idata_n2925,
         oc8051_ram_top1_oc8051_idata_n2924,
         oc8051_ram_top1_oc8051_idata_n2923,
         oc8051_ram_top1_oc8051_idata_n2922,
         oc8051_ram_top1_oc8051_idata_n2921,
         oc8051_ram_top1_oc8051_idata_n2920,
         oc8051_ram_top1_oc8051_idata_n2919,
         oc8051_ram_top1_oc8051_idata_n2918,
         oc8051_ram_top1_oc8051_idata_n2917,
         oc8051_ram_top1_oc8051_idata_n2916,
         oc8051_ram_top1_oc8051_idata_n2915,
         oc8051_ram_top1_oc8051_idata_n2914,
         oc8051_ram_top1_oc8051_idata_n2913,
         oc8051_ram_top1_oc8051_idata_n2912,
         oc8051_ram_top1_oc8051_idata_n2911,
         oc8051_ram_top1_oc8051_idata_n2910,
         oc8051_ram_top1_oc8051_idata_n2909,
         oc8051_ram_top1_oc8051_idata_n2908,
         oc8051_ram_top1_oc8051_idata_n2907,
         oc8051_ram_top1_oc8051_idata_n2906,
         oc8051_ram_top1_oc8051_idata_n2905,
         oc8051_ram_top1_oc8051_idata_n2904,
         oc8051_ram_top1_oc8051_idata_n2903,
         oc8051_ram_top1_oc8051_idata_n2902,
         oc8051_ram_top1_oc8051_idata_n2901,
         oc8051_ram_top1_oc8051_idata_n2900,
         oc8051_ram_top1_oc8051_idata_n2899,
         oc8051_ram_top1_oc8051_idata_n2898,
         oc8051_ram_top1_oc8051_idata_n2897,
         oc8051_ram_top1_oc8051_idata_n2896,
         oc8051_ram_top1_oc8051_idata_n2895,
         oc8051_ram_top1_oc8051_idata_n2894,
         oc8051_ram_top1_oc8051_idata_n2893,
         oc8051_ram_top1_oc8051_idata_n2892,
         oc8051_ram_top1_oc8051_idata_n2891,
         oc8051_ram_top1_oc8051_idata_n2890,
         oc8051_ram_top1_oc8051_idata_n2889,
         oc8051_ram_top1_oc8051_idata_n2888,
         oc8051_ram_top1_oc8051_idata_n2887,
         oc8051_ram_top1_oc8051_idata_n2886,
         oc8051_ram_top1_oc8051_idata_n2885,
         oc8051_ram_top1_oc8051_idata_n2884,
         oc8051_ram_top1_oc8051_idata_n2883,
         oc8051_ram_top1_oc8051_idata_n2882,
         oc8051_ram_top1_oc8051_idata_n2881,
         oc8051_ram_top1_oc8051_idata_n2880,
         oc8051_ram_top1_oc8051_idata_n2879,
         oc8051_ram_top1_oc8051_idata_n2878,
         oc8051_ram_top1_oc8051_idata_n2877,
         oc8051_ram_top1_oc8051_idata_n2876,
         oc8051_ram_top1_oc8051_idata_n2875,
         oc8051_ram_top1_oc8051_idata_n2874,
         oc8051_ram_top1_oc8051_idata_n2873,
         oc8051_ram_top1_oc8051_idata_n2872,
         oc8051_ram_top1_oc8051_idata_n2871,
         oc8051_ram_top1_oc8051_idata_n2870,
         oc8051_ram_top1_oc8051_idata_n2869,
         oc8051_ram_top1_oc8051_idata_n2868,
         oc8051_ram_top1_oc8051_idata_n2867,
         oc8051_ram_top1_oc8051_idata_n2866,
         oc8051_ram_top1_oc8051_idata_n2865,
         oc8051_ram_top1_oc8051_idata_n2864,
         oc8051_ram_top1_oc8051_idata_n2863,
         oc8051_ram_top1_oc8051_idata_n2862,
         oc8051_ram_top1_oc8051_idata_n2861,
         oc8051_ram_top1_oc8051_idata_n2860,
         oc8051_ram_top1_oc8051_idata_n2859,
         oc8051_ram_top1_oc8051_idata_n2858,
         oc8051_ram_top1_oc8051_idata_n2857,
         oc8051_ram_top1_oc8051_idata_n2856,
         oc8051_ram_top1_oc8051_idata_n2855,
         oc8051_ram_top1_oc8051_idata_n2854,
         oc8051_ram_top1_oc8051_idata_n2853,
         oc8051_ram_top1_oc8051_idata_n2852,
         oc8051_ram_top1_oc8051_idata_n2851,
         oc8051_ram_top1_oc8051_idata_n2850,
         oc8051_ram_top1_oc8051_idata_n2849,
         oc8051_ram_top1_oc8051_idata_n2848,
         oc8051_ram_top1_oc8051_idata_n2847,
         oc8051_ram_top1_oc8051_idata_n2846,
         oc8051_ram_top1_oc8051_idata_n2845,
         oc8051_ram_top1_oc8051_idata_n2844,
         oc8051_ram_top1_oc8051_idata_n2843,
         oc8051_ram_top1_oc8051_idata_n2842,
         oc8051_ram_top1_oc8051_idata_n2841,
         oc8051_ram_top1_oc8051_idata_n2840,
         oc8051_ram_top1_oc8051_idata_n2839,
         oc8051_ram_top1_oc8051_idata_n2838,
         oc8051_ram_top1_oc8051_idata_n2837,
         oc8051_ram_top1_oc8051_idata_n2836,
         oc8051_ram_top1_oc8051_idata_n2835,
         oc8051_ram_top1_oc8051_idata_n2834,
         oc8051_ram_top1_oc8051_idata_n2833,
         oc8051_ram_top1_oc8051_idata_n2832,
         oc8051_ram_top1_oc8051_idata_n2831,
         oc8051_ram_top1_oc8051_idata_n2830,
         oc8051_ram_top1_oc8051_idata_n2829,
         oc8051_ram_top1_oc8051_idata_n2828,
         oc8051_ram_top1_oc8051_idata_n2827,
         oc8051_ram_top1_oc8051_idata_n2826,
         oc8051_ram_top1_oc8051_idata_n2825,
         oc8051_ram_top1_oc8051_idata_n2824,
         oc8051_ram_top1_oc8051_idata_n2823,
         oc8051_ram_top1_oc8051_idata_n2822,
         oc8051_ram_top1_oc8051_idata_n2821,
         oc8051_ram_top1_oc8051_idata_n2820,
         oc8051_ram_top1_oc8051_idata_n2819,
         oc8051_ram_top1_oc8051_idata_n2818,
         oc8051_ram_top1_oc8051_idata_n2817,
         oc8051_ram_top1_oc8051_idata_n2816,
         oc8051_ram_top1_oc8051_idata_n2815,
         oc8051_ram_top1_oc8051_idata_n2814,
         oc8051_ram_top1_oc8051_idata_n2813,
         oc8051_ram_top1_oc8051_idata_n2812,
         oc8051_ram_top1_oc8051_idata_n2811,
         oc8051_ram_top1_oc8051_idata_n2810,
         oc8051_ram_top1_oc8051_idata_n2809,
         oc8051_ram_top1_oc8051_idata_n2808,
         oc8051_ram_top1_oc8051_idata_n2807,
         oc8051_ram_top1_oc8051_idata_n2806,
         oc8051_ram_top1_oc8051_idata_n2805,
         oc8051_ram_top1_oc8051_idata_n2804,
         oc8051_ram_top1_oc8051_idata_n2803,
         oc8051_ram_top1_oc8051_idata_n2802,
         oc8051_ram_top1_oc8051_idata_n2801,
         oc8051_ram_top1_oc8051_idata_n2800,
         oc8051_ram_top1_oc8051_idata_n2799,
         oc8051_ram_top1_oc8051_idata_n2798,
         oc8051_ram_top1_oc8051_idata_n2797,
         oc8051_ram_top1_oc8051_idata_n2796,
         oc8051_ram_top1_oc8051_idata_n2795,
         oc8051_ram_top1_oc8051_idata_n2794,
         oc8051_ram_top1_oc8051_idata_n2793,
         oc8051_ram_top1_oc8051_idata_n2792,
         oc8051_ram_top1_oc8051_idata_n2791,
         oc8051_ram_top1_oc8051_idata_n2790,
         oc8051_ram_top1_oc8051_idata_n2789,
         oc8051_ram_top1_oc8051_idata_n2788,
         oc8051_ram_top1_oc8051_idata_n2787,
         oc8051_ram_top1_oc8051_idata_n2786,
         oc8051_ram_top1_oc8051_idata_n2785,
         oc8051_ram_top1_oc8051_idata_n2784,
         oc8051_ram_top1_oc8051_idata_n2783,
         oc8051_ram_top1_oc8051_idata_n2782,
         oc8051_ram_top1_oc8051_idata_n2781,
         oc8051_ram_top1_oc8051_idata_n2780,
         oc8051_ram_top1_oc8051_idata_n2779,
         oc8051_ram_top1_oc8051_idata_n2778,
         oc8051_ram_top1_oc8051_idata_n2777,
         oc8051_ram_top1_oc8051_idata_n2776,
         oc8051_ram_top1_oc8051_idata_n2775,
         oc8051_ram_top1_oc8051_idata_n2774,
         oc8051_ram_top1_oc8051_idata_n2773,
         oc8051_ram_top1_oc8051_idata_n2772,
         oc8051_ram_top1_oc8051_idata_n2771,
         oc8051_ram_top1_oc8051_idata_n2770,
         oc8051_ram_top1_oc8051_idata_n2769,
         oc8051_ram_top1_oc8051_idata_n2768,
         oc8051_ram_top1_oc8051_idata_n2767,
         oc8051_ram_top1_oc8051_idata_n2766,
         oc8051_ram_top1_oc8051_idata_n2765,
         oc8051_ram_top1_oc8051_idata_n2764,
         oc8051_ram_top1_oc8051_idata_n2763,
         oc8051_ram_top1_oc8051_idata_n2762,
         oc8051_ram_top1_oc8051_idata_n2761,
         oc8051_ram_top1_oc8051_idata_n2760,
         oc8051_ram_top1_oc8051_idata_n2759,
         oc8051_ram_top1_oc8051_idata_n2758,
         oc8051_ram_top1_oc8051_idata_n2757,
         oc8051_ram_top1_oc8051_idata_n2756,
         oc8051_ram_top1_oc8051_idata_n2755,
         oc8051_ram_top1_oc8051_idata_n2754,
         oc8051_ram_top1_oc8051_idata_n2753,
         oc8051_ram_top1_oc8051_idata_n2752,
         oc8051_ram_top1_oc8051_idata_n2751,
         oc8051_ram_top1_oc8051_idata_n2750,
         oc8051_ram_top1_oc8051_idata_n2749,
         oc8051_ram_top1_oc8051_idata_n2748,
         oc8051_ram_top1_oc8051_idata_n2747,
         oc8051_ram_top1_oc8051_idata_n2746,
         oc8051_ram_top1_oc8051_idata_n2745,
         oc8051_ram_top1_oc8051_idata_n2744,
         oc8051_ram_top1_oc8051_idata_n2743,
         oc8051_ram_top1_oc8051_idata_n2742,
         oc8051_ram_top1_oc8051_idata_n2741,
         oc8051_ram_top1_oc8051_idata_n2740,
         oc8051_ram_top1_oc8051_idata_n2739,
         oc8051_ram_top1_oc8051_idata_n2738,
         oc8051_ram_top1_oc8051_idata_n2737,
         oc8051_ram_top1_oc8051_idata_n2736,
         oc8051_ram_top1_oc8051_idata_n2735,
         oc8051_ram_top1_oc8051_idata_n2734,
         oc8051_ram_top1_oc8051_idata_n2733,
         oc8051_ram_top1_oc8051_idata_n2732,
         oc8051_ram_top1_oc8051_idata_n2731,
         oc8051_ram_top1_oc8051_idata_n2730,
         oc8051_ram_top1_oc8051_idata_n2729,
         oc8051_ram_top1_oc8051_idata_n2728,
         oc8051_ram_top1_oc8051_idata_n2727,
         oc8051_ram_top1_oc8051_idata_n2726,
         oc8051_ram_top1_oc8051_idata_n2725,
         oc8051_ram_top1_oc8051_idata_n2724,
         oc8051_ram_top1_oc8051_idata_n2723,
         oc8051_ram_top1_oc8051_idata_n2722,
         oc8051_ram_top1_oc8051_idata_n2721,
         oc8051_ram_top1_oc8051_idata_n2720,
         oc8051_ram_top1_oc8051_idata_n2719,
         oc8051_ram_top1_oc8051_idata_n2718,
         oc8051_ram_top1_oc8051_idata_n2717,
         oc8051_ram_top1_oc8051_idata_n2716,
         oc8051_ram_top1_oc8051_idata_n2715,
         oc8051_ram_top1_oc8051_idata_n2714,
         oc8051_ram_top1_oc8051_idata_n2713,
         oc8051_ram_top1_oc8051_idata_n2712,
         oc8051_ram_top1_oc8051_idata_n2711,
         oc8051_ram_top1_oc8051_idata_n2710,
         oc8051_ram_top1_oc8051_idata_n2709,
         oc8051_ram_top1_oc8051_idata_n2708,
         oc8051_ram_top1_oc8051_idata_n2707,
         oc8051_ram_top1_oc8051_idata_n2706,
         oc8051_ram_top1_oc8051_idata_n2705,
         oc8051_ram_top1_oc8051_idata_n2704,
         oc8051_ram_top1_oc8051_idata_n2703,
         oc8051_ram_top1_oc8051_idata_n2702,
         oc8051_ram_top1_oc8051_idata_n2701,
         oc8051_ram_top1_oc8051_idata_n2700,
         oc8051_ram_top1_oc8051_idata_n2699,
         oc8051_ram_top1_oc8051_idata_n2698,
         oc8051_ram_top1_oc8051_idata_n2697,
         oc8051_ram_top1_oc8051_idata_n2696,
         oc8051_ram_top1_oc8051_idata_n2695,
         oc8051_ram_top1_oc8051_idata_n2694,
         oc8051_ram_top1_oc8051_idata_n2693,
         oc8051_ram_top1_oc8051_idata_n2692,
         oc8051_ram_top1_oc8051_idata_n2691,
         oc8051_ram_top1_oc8051_idata_n2690,
         oc8051_ram_top1_oc8051_idata_n2689,
         oc8051_ram_top1_oc8051_idata_n2688,
         oc8051_ram_top1_oc8051_idata_n2687,
         oc8051_ram_top1_oc8051_idata_n2686,
         oc8051_ram_top1_oc8051_idata_n2685,
         oc8051_ram_top1_oc8051_idata_n2684,
         oc8051_ram_top1_oc8051_idata_n2683,
         oc8051_ram_top1_oc8051_idata_n2682,
         oc8051_ram_top1_oc8051_idata_n2681,
         oc8051_ram_top1_oc8051_idata_n2680,
         oc8051_ram_top1_oc8051_idata_n2679,
         oc8051_ram_top1_oc8051_idata_n2678,
         oc8051_ram_top1_oc8051_idata_n2677,
         oc8051_ram_top1_oc8051_idata_n2676,
         oc8051_ram_top1_oc8051_idata_n2675,
         oc8051_ram_top1_oc8051_idata_n2674,
         oc8051_ram_top1_oc8051_idata_n2673,
         oc8051_ram_top1_oc8051_idata_n2672,
         oc8051_ram_top1_oc8051_idata_n2671,
         oc8051_ram_top1_oc8051_idata_n2670,
         oc8051_ram_top1_oc8051_idata_n2669,
         oc8051_ram_top1_oc8051_idata_n2668,
         oc8051_ram_top1_oc8051_idata_n2667,
         oc8051_ram_top1_oc8051_idata_n2666,
         oc8051_ram_top1_oc8051_idata_n2665,
         oc8051_ram_top1_oc8051_idata_n2664,
         oc8051_ram_top1_oc8051_idata_n2663,
         oc8051_ram_top1_oc8051_idata_n2662,
         oc8051_ram_top1_oc8051_idata_n2661,
         oc8051_ram_top1_oc8051_idata_n2660,
         oc8051_ram_top1_oc8051_idata_n2659,
         oc8051_ram_top1_oc8051_idata_n2658,
         oc8051_ram_top1_oc8051_idata_n2657,
         oc8051_ram_top1_oc8051_idata_n2656,
         oc8051_ram_top1_oc8051_idata_n2655,
         oc8051_ram_top1_oc8051_idata_n2654,
         oc8051_ram_top1_oc8051_idata_n2653,
         oc8051_ram_top1_oc8051_idata_n2652,
         oc8051_ram_top1_oc8051_idata_n2651,
         oc8051_ram_top1_oc8051_idata_n2650,
         oc8051_ram_top1_oc8051_idata_n2649,
         oc8051_ram_top1_oc8051_idata_n2648,
         oc8051_ram_top1_oc8051_idata_n2647,
         oc8051_ram_top1_oc8051_idata_n2646,
         oc8051_ram_top1_oc8051_idata_n2645,
         oc8051_ram_top1_oc8051_idata_n2644,
         oc8051_ram_top1_oc8051_idata_n2643,
         oc8051_ram_top1_oc8051_idata_n2642,
         oc8051_ram_top1_oc8051_idata_n2641,
         oc8051_ram_top1_oc8051_idata_n2640,
         oc8051_ram_top1_oc8051_idata_n2639,
         oc8051_ram_top1_oc8051_idata_n2638,
         oc8051_ram_top1_oc8051_idata_n2637,
         oc8051_ram_top1_oc8051_idata_n2636,
         oc8051_ram_top1_oc8051_idata_n2635,
         oc8051_ram_top1_oc8051_idata_n2634,
         oc8051_ram_top1_oc8051_idata_n2633,
         oc8051_ram_top1_oc8051_idata_n2632,
         oc8051_ram_top1_oc8051_idata_n2631,
         oc8051_ram_top1_oc8051_idata_n2630,
         oc8051_ram_top1_oc8051_idata_n2629,
         oc8051_ram_top1_oc8051_idata_n2628,
         oc8051_ram_top1_oc8051_idata_n2627,
         oc8051_ram_top1_oc8051_idata_n2626,
         oc8051_ram_top1_oc8051_idata_n2625,
         oc8051_ram_top1_oc8051_idata_n2624,
         oc8051_ram_top1_oc8051_idata_n2623,
         oc8051_ram_top1_oc8051_idata_n2622,
         oc8051_ram_top1_oc8051_idata_n2621,
         oc8051_ram_top1_oc8051_idata_n2620,
         oc8051_ram_top1_oc8051_idata_n2619,
         oc8051_ram_top1_oc8051_idata_n2618,
         oc8051_ram_top1_oc8051_idata_n2617,
         oc8051_ram_top1_oc8051_idata_n2616,
         oc8051_ram_top1_oc8051_idata_n2615,
         oc8051_ram_top1_oc8051_idata_n2614,
         oc8051_ram_top1_oc8051_idata_n2613,
         oc8051_ram_top1_oc8051_idata_n2612,
         oc8051_ram_top1_oc8051_idata_n2611,
         oc8051_ram_top1_oc8051_idata_n2610,
         oc8051_ram_top1_oc8051_idata_n2609,
         oc8051_ram_top1_oc8051_idata_n2608,
         oc8051_ram_top1_oc8051_idata_n2607,
         oc8051_ram_top1_oc8051_idata_n2606,
         oc8051_ram_top1_oc8051_idata_n2605,
         oc8051_ram_top1_oc8051_idata_n2604,
         oc8051_ram_top1_oc8051_idata_n2603,
         oc8051_ram_top1_oc8051_idata_n2602,
         oc8051_ram_top1_oc8051_idata_n2601,
         oc8051_ram_top1_oc8051_idata_n2600,
         oc8051_ram_top1_oc8051_idata_n2599,
         oc8051_ram_top1_oc8051_idata_n2598,
         oc8051_ram_top1_oc8051_idata_n2597,
         oc8051_ram_top1_oc8051_idata_n2596,
         oc8051_ram_top1_oc8051_idata_n2595,
         oc8051_ram_top1_oc8051_idata_n2594,
         oc8051_ram_top1_oc8051_idata_n2593,
         oc8051_ram_top1_oc8051_idata_n2592,
         oc8051_ram_top1_oc8051_idata_n2591,
         oc8051_ram_top1_oc8051_idata_n2590,
         oc8051_ram_top1_oc8051_idata_n2589,
         oc8051_ram_top1_oc8051_idata_n2588,
         oc8051_ram_top1_oc8051_idata_n2587,
         oc8051_ram_top1_oc8051_idata_n2586,
         oc8051_ram_top1_oc8051_idata_n2585,
         oc8051_ram_top1_oc8051_idata_n2584,
         oc8051_ram_top1_oc8051_idata_n2583,
         oc8051_ram_top1_oc8051_idata_n2582,
         oc8051_ram_top1_oc8051_idata_n2581,
         oc8051_ram_top1_oc8051_idata_n2580,
         oc8051_ram_top1_oc8051_idata_n2579,
         oc8051_ram_top1_oc8051_idata_n2578,
         oc8051_ram_top1_oc8051_idata_n2577,
         oc8051_ram_top1_oc8051_idata_n2576,
         oc8051_ram_top1_oc8051_idata_n2575,
         oc8051_ram_top1_oc8051_idata_n2574,
         oc8051_ram_top1_oc8051_idata_n2573,
         oc8051_ram_top1_oc8051_idata_n2572,
         oc8051_ram_top1_oc8051_idata_n2571,
         oc8051_ram_top1_oc8051_idata_n2570,
         oc8051_ram_top1_oc8051_idata_n2569,
         oc8051_ram_top1_oc8051_idata_n2568,
         oc8051_ram_top1_oc8051_idata_n2567,
         oc8051_ram_top1_oc8051_idata_n2566,
         oc8051_ram_top1_oc8051_idata_n2565,
         oc8051_ram_top1_oc8051_idata_n2564,
         oc8051_ram_top1_oc8051_idata_n2563,
         oc8051_ram_top1_oc8051_idata_n2562,
         oc8051_ram_top1_oc8051_idata_n2561,
         oc8051_ram_top1_oc8051_idata_n2560,
         oc8051_ram_top1_oc8051_idata_n2559,
         oc8051_ram_top1_oc8051_idata_n2558,
         oc8051_ram_top1_oc8051_idata_n2557,
         oc8051_ram_top1_oc8051_idata_n2556,
         oc8051_ram_top1_oc8051_idata_n2555,
         oc8051_ram_top1_oc8051_idata_n2554,
         oc8051_ram_top1_oc8051_idata_n2553,
         oc8051_ram_top1_oc8051_idata_n2552,
         oc8051_ram_top1_oc8051_idata_n2551,
         oc8051_ram_top1_oc8051_idata_n2550,
         oc8051_ram_top1_oc8051_idata_n2549,
         oc8051_ram_top1_oc8051_idata_n2548,
         oc8051_ram_top1_oc8051_idata_n2547,
         oc8051_ram_top1_oc8051_idata_n2546,
         oc8051_ram_top1_oc8051_idata_n2545,
         oc8051_ram_top1_oc8051_idata_n2544,
         oc8051_ram_top1_oc8051_idata_n2543,
         oc8051_ram_top1_oc8051_idata_n2542,
         oc8051_ram_top1_oc8051_idata_n2541,
         oc8051_ram_top1_oc8051_idata_n2540,
         oc8051_ram_top1_oc8051_idata_n2539,
         oc8051_ram_top1_oc8051_idata_n2538,
         oc8051_ram_top1_oc8051_idata_n2537,
         oc8051_ram_top1_oc8051_idata_n2536,
         oc8051_ram_top1_oc8051_idata_n2535,
         oc8051_ram_top1_oc8051_idata_n2534,
         oc8051_ram_top1_oc8051_idata_n2533,
         oc8051_ram_top1_oc8051_idata_n2532,
         oc8051_ram_top1_oc8051_idata_n2531,
         oc8051_ram_top1_oc8051_idata_n2530,
         oc8051_ram_top1_oc8051_idata_n2529,
         oc8051_ram_top1_oc8051_idata_n2528,
         oc8051_ram_top1_oc8051_idata_n2527,
         oc8051_ram_top1_oc8051_idata_n2526,
         oc8051_ram_top1_oc8051_idata_n2525,
         oc8051_ram_top1_oc8051_idata_n2524,
         oc8051_ram_top1_oc8051_idata_n2523,
         oc8051_ram_top1_oc8051_idata_n2522,
         oc8051_ram_top1_oc8051_idata_n2521,
         oc8051_ram_top1_oc8051_idata_n2520,
         oc8051_ram_top1_oc8051_idata_n2519,
         oc8051_ram_top1_oc8051_idata_n2518,
         oc8051_ram_top1_oc8051_idata_n2517,
         oc8051_ram_top1_oc8051_idata_n2516,
         oc8051_ram_top1_oc8051_idata_n2515,
         oc8051_ram_top1_oc8051_idata_n2514,
         oc8051_ram_top1_oc8051_idata_n2513,
         oc8051_ram_top1_oc8051_idata_n2512,
         oc8051_ram_top1_oc8051_idata_n2511,
         oc8051_ram_top1_oc8051_idata_n2510,
         oc8051_ram_top1_oc8051_idata_n2509,
         oc8051_ram_top1_oc8051_idata_n2508,
         oc8051_ram_top1_oc8051_idata_n2507,
         oc8051_ram_top1_oc8051_idata_n2506,
         oc8051_ram_top1_oc8051_idata_n2505,
         oc8051_ram_top1_oc8051_idata_n2504,
         oc8051_ram_top1_oc8051_idata_n2503,
         oc8051_ram_top1_oc8051_idata_n2502,
         oc8051_ram_top1_oc8051_idata_n2501,
         oc8051_ram_top1_oc8051_idata_n2500,
         oc8051_ram_top1_oc8051_idata_n2499,
         oc8051_ram_top1_oc8051_idata_n2498,
         oc8051_ram_top1_oc8051_idata_n2497,
         oc8051_ram_top1_oc8051_idata_n2496,
         oc8051_ram_top1_oc8051_idata_n2495,
         oc8051_ram_top1_oc8051_idata_n2494,
         oc8051_ram_top1_oc8051_idata_n2493,
         oc8051_ram_top1_oc8051_idata_n2492,
         oc8051_ram_top1_oc8051_idata_n2491,
         oc8051_ram_top1_oc8051_idata_n2490,
         oc8051_ram_top1_oc8051_idata_n2489,
         oc8051_ram_top1_oc8051_idata_n2488,
         oc8051_ram_top1_oc8051_idata_n2487,
         oc8051_ram_top1_oc8051_idata_n2486,
         oc8051_ram_top1_oc8051_idata_n2485,
         oc8051_ram_top1_oc8051_idata_n2484,
         oc8051_ram_top1_oc8051_idata_n2483,
         oc8051_ram_top1_oc8051_idata_n2482,
         oc8051_ram_top1_oc8051_idata_n2481,
         oc8051_ram_top1_oc8051_idata_n2480,
         oc8051_ram_top1_oc8051_idata_n2479,
         oc8051_ram_top1_oc8051_idata_n2478,
         oc8051_ram_top1_oc8051_idata_n2477,
         oc8051_ram_top1_oc8051_idata_n2476,
         oc8051_ram_top1_oc8051_idata_n2475, oc8051_ram_top1_oc8051_idata_n515,
         oc8051_ram_top1_oc8051_idata_n514, oc8051_ram_top1_oc8051_idata_n513,
         oc8051_ram_top1_oc8051_idata_n512, oc8051_ram_top1_oc8051_idata_n511,
         oc8051_ram_top1_oc8051_idata_n510, oc8051_ram_top1_oc8051_idata_n509,
         oc8051_ram_top1_oc8051_idata_n508, oc8051_ram_top1_oc8051_idata_n507,
         oc8051_ram_top1_oc8051_idata_n506, oc8051_ram_top1_oc8051_idata_n505,
         oc8051_ram_top1_oc8051_idata_n504, oc8051_ram_top1_oc8051_idata_n503,
         oc8051_ram_top1_oc8051_idata_n502, oc8051_ram_top1_oc8051_idata_n501,
         oc8051_ram_top1_oc8051_idata_n500, oc8051_ram_top1_oc8051_idata_n499,
         oc8051_ram_top1_oc8051_idata_n498, oc8051_ram_top1_oc8051_idata_n497,
         oc8051_ram_top1_oc8051_idata_n496, oc8051_ram_top1_oc8051_idata_n495,
         oc8051_ram_top1_oc8051_idata_n494, oc8051_ram_top1_oc8051_idata_n493,
         oc8051_ram_top1_oc8051_idata_n492, oc8051_ram_top1_oc8051_idata_n491,
         oc8051_ram_top1_oc8051_idata_n490, oc8051_ram_top1_oc8051_idata_n489,
         oc8051_ram_top1_oc8051_idata_n488, oc8051_ram_top1_oc8051_idata_n487,
         oc8051_ram_top1_oc8051_idata_n486, oc8051_ram_top1_oc8051_idata_n485,
         oc8051_ram_top1_oc8051_idata_n484, oc8051_ram_top1_oc8051_idata_n483,
         oc8051_ram_top1_oc8051_idata_n482, oc8051_ram_top1_oc8051_idata_n481,
         oc8051_ram_top1_oc8051_idata_n480, oc8051_ram_top1_oc8051_idata_n479,
         oc8051_ram_top1_oc8051_idata_n478, oc8051_ram_top1_oc8051_idata_n477,
         oc8051_ram_top1_oc8051_idata_n476, oc8051_ram_top1_oc8051_idata_n475,
         oc8051_ram_top1_oc8051_idata_n474, oc8051_ram_top1_oc8051_idata_n473,
         oc8051_ram_top1_oc8051_idata_n472, oc8051_ram_top1_oc8051_idata_n471,
         oc8051_ram_top1_oc8051_idata_n470, oc8051_ram_top1_oc8051_idata_n469,
         oc8051_ram_top1_oc8051_idata_n468, oc8051_ram_top1_oc8051_idata_n467,
         oc8051_ram_top1_oc8051_idata_n466, oc8051_ram_top1_oc8051_idata_n465,
         oc8051_ram_top1_oc8051_idata_n464, oc8051_ram_top1_oc8051_idata_n463,
         oc8051_ram_top1_oc8051_idata_n462, oc8051_ram_top1_oc8051_idata_n461,
         oc8051_ram_top1_oc8051_idata_n460, oc8051_ram_top1_oc8051_idata_n459,
         oc8051_ram_top1_oc8051_idata_n458, oc8051_ram_top1_oc8051_idata_n457,
         oc8051_ram_top1_oc8051_idata_n456, oc8051_ram_top1_oc8051_idata_n455,
         oc8051_ram_top1_oc8051_idata_n454, oc8051_ram_top1_oc8051_idata_n453,
         oc8051_ram_top1_oc8051_idata_n452, oc8051_ram_top1_oc8051_idata_n451,
         oc8051_ram_top1_oc8051_idata_n450, oc8051_ram_top1_oc8051_idata_n449,
         oc8051_ram_top1_oc8051_idata_n448, oc8051_ram_top1_oc8051_idata_n447,
         oc8051_ram_top1_oc8051_idata_n446, oc8051_ram_top1_oc8051_idata_n445,
         oc8051_ram_top1_oc8051_idata_n444, oc8051_ram_top1_oc8051_idata_n443,
         oc8051_ram_top1_oc8051_idata_n442, oc8051_ram_top1_oc8051_idata_n441,
         oc8051_ram_top1_oc8051_idata_n440, oc8051_ram_top1_oc8051_idata_n439,
         oc8051_ram_top1_oc8051_idata_n438, oc8051_ram_top1_oc8051_idata_n437,
         oc8051_ram_top1_oc8051_idata_n436, oc8051_ram_top1_oc8051_idata_n435,
         oc8051_ram_top1_oc8051_idata_n434, oc8051_ram_top1_oc8051_idata_n433,
         oc8051_ram_top1_oc8051_idata_n432, oc8051_ram_top1_oc8051_idata_n431,
         oc8051_ram_top1_oc8051_idata_n430, oc8051_ram_top1_oc8051_idata_n429,
         oc8051_ram_top1_oc8051_idata_n428, oc8051_ram_top1_oc8051_idata_n427,
         oc8051_ram_top1_oc8051_idata_n426, oc8051_ram_top1_oc8051_idata_n425,
         oc8051_ram_top1_oc8051_idata_n424, oc8051_ram_top1_oc8051_idata_n423,
         oc8051_ram_top1_oc8051_idata_n422, oc8051_ram_top1_oc8051_idata_n421,
         oc8051_ram_top1_oc8051_idata_n420, oc8051_ram_top1_oc8051_idata_n419,
         oc8051_ram_top1_oc8051_idata_n418, oc8051_ram_top1_oc8051_idata_n417,
         oc8051_ram_top1_oc8051_idata_n416, oc8051_ram_top1_oc8051_idata_n415,
         oc8051_ram_top1_oc8051_idata_n414, oc8051_ram_top1_oc8051_idata_n413,
         oc8051_ram_top1_oc8051_idata_n412, oc8051_ram_top1_oc8051_idata_n411,
         oc8051_ram_top1_oc8051_idata_n410, oc8051_ram_top1_oc8051_idata_n409,
         oc8051_ram_top1_oc8051_idata_n408, oc8051_ram_top1_oc8051_idata_n407,
         oc8051_ram_top1_oc8051_idata_n406, oc8051_ram_top1_oc8051_idata_n405,
         oc8051_ram_top1_oc8051_idata_n404, oc8051_ram_top1_oc8051_idata_n403,
         oc8051_ram_top1_oc8051_idata_n402, oc8051_ram_top1_oc8051_idata_n401,
         oc8051_ram_top1_oc8051_idata_n400, oc8051_ram_top1_oc8051_idata_n399,
         oc8051_ram_top1_oc8051_idata_n398, oc8051_ram_top1_oc8051_idata_n397,
         oc8051_ram_top1_oc8051_idata_n396, oc8051_ram_top1_oc8051_idata_n395,
         oc8051_ram_top1_oc8051_idata_n394, oc8051_ram_top1_oc8051_idata_n393,
         oc8051_ram_top1_oc8051_idata_n392, oc8051_ram_top1_oc8051_idata_n391,
         oc8051_ram_top1_oc8051_idata_n390, oc8051_ram_top1_oc8051_idata_n389,
         oc8051_ram_top1_oc8051_idata_n388, oc8051_ram_top1_oc8051_idata_n387,
         oc8051_ram_top1_oc8051_idata_n386, oc8051_ram_top1_oc8051_idata_n385,
         oc8051_ram_top1_oc8051_idata_n384, oc8051_ram_top1_oc8051_idata_n383,
         oc8051_ram_top1_oc8051_idata_n382, oc8051_ram_top1_oc8051_idata_n381,
         oc8051_ram_top1_oc8051_idata_n380, oc8051_ram_top1_oc8051_idata_n379,
         oc8051_ram_top1_oc8051_idata_n378, oc8051_ram_top1_oc8051_idata_n377,
         oc8051_ram_top1_oc8051_idata_n376, oc8051_ram_top1_oc8051_idata_n375,
         oc8051_ram_top1_oc8051_idata_n374, oc8051_ram_top1_oc8051_idata_n373,
         oc8051_ram_top1_oc8051_idata_n372, oc8051_ram_top1_oc8051_idata_n371,
         oc8051_ram_top1_oc8051_idata_n370, oc8051_ram_top1_oc8051_idata_n369,
         oc8051_ram_top1_oc8051_idata_n368, oc8051_ram_top1_oc8051_idata_n367,
         oc8051_ram_top1_oc8051_idata_n366, oc8051_ram_top1_oc8051_idata_n365,
         oc8051_ram_top1_oc8051_idata_n364, oc8051_ram_top1_oc8051_idata_n363,
         oc8051_ram_top1_oc8051_idata_n362, oc8051_ram_top1_oc8051_idata_n361,
         oc8051_ram_top1_oc8051_idata_n360, oc8051_ram_top1_oc8051_idata_n359,
         oc8051_ram_top1_oc8051_idata_n358, oc8051_ram_top1_oc8051_idata_n357,
         oc8051_ram_top1_oc8051_idata_n356, oc8051_ram_top1_oc8051_idata_n355,
         oc8051_ram_top1_oc8051_idata_n354, oc8051_ram_top1_oc8051_idata_n353,
         oc8051_ram_top1_oc8051_idata_n352, oc8051_ram_top1_oc8051_idata_n351,
         oc8051_ram_top1_oc8051_idata_n350, oc8051_ram_top1_oc8051_idata_n349,
         oc8051_ram_top1_oc8051_idata_n348, oc8051_ram_top1_oc8051_idata_n347,
         oc8051_ram_top1_oc8051_idata_n346, oc8051_ram_top1_oc8051_idata_n345,
         oc8051_ram_top1_oc8051_idata_n344, oc8051_ram_top1_oc8051_idata_n343,
         oc8051_ram_top1_oc8051_idata_n342, oc8051_ram_top1_oc8051_idata_n341,
         oc8051_ram_top1_oc8051_idata_n340, oc8051_ram_top1_oc8051_idata_n339,
         oc8051_ram_top1_oc8051_idata_n338, oc8051_ram_top1_oc8051_idata_n337,
         oc8051_ram_top1_oc8051_idata_n336, oc8051_ram_top1_oc8051_idata_n335,
         oc8051_ram_top1_oc8051_idata_n334, oc8051_ram_top1_oc8051_idata_n333,
         oc8051_ram_top1_oc8051_idata_n332, oc8051_ram_top1_oc8051_idata_n331,
         oc8051_ram_top1_oc8051_idata_n330, oc8051_ram_top1_oc8051_idata_n329,
         oc8051_ram_top1_oc8051_idata_n328, oc8051_ram_top1_oc8051_idata_n327,
         oc8051_ram_top1_oc8051_idata_n326, oc8051_ram_top1_oc8051_idata_n325,
         oc8051_ram_top1_oc8051_idata_n324, oc8051_ram_top1_oc8051_idata_n323,
         oc8051_ram_top1_oc8051_idata_n322, oc8051_ram_top1_oc8051_idata_n321,
         oc8051_ram_top1_oc8051_idata_n320, oc8051_ram_top1_oc8051_idata_n319,
         oc8051_ram_top1_oc8051_idata_n318, oc8051_ram_top1_oc8051_idata_n317,
         oc8051_ram_top1_oc8051_idata_n316, oc8051_ram_top1_oc8051_idata_n315,
         oc8051_ram_top1_oc8051_idata_n314, oc8051_ram_top1_oc8051_idata_n313,
         oc8051_ram_top1_oc8051_idata_n312, oc8051_ram_top1_oc8051_idata_n311,
         oc8051_ram_top1_oc8051_idata_n310, oc8051_ram_top1_oc8051_idata_n309,
         oc8051_ram_top1_oc8051_idata_n308, oc8051_ram_top1_oc8051_idata_n307,
         oc8051_ram_top1_oc8051_idata_n306, oc8051_ram_top1_oc8051_idata_n305,
         oc8051_ram_top1_oc8051_idata_n304, oc8051_ram_top1_oc8051_idata_n303,
         oc8051_ram_top1_oc8051_idata_n302, oc8051_ram_top1_oc8051_idata_n301,
         oc8051_ram_top1_oc8051_idata_n300, oc8051_ram_top1_oc8051_idata_n299,
         oc8051_ram_top1_oc8051_idata_n298, oc8051_ram_top1_oc8051_idata_n297,
         oc8051_ram_top1_oc8051_idata_n296, oc8051_ram_top1_oc8051_idata_n295,
         oc8051_ram_top1_oc8051_idata_n294, oc8051_ram_top1_oc8051_idata_n293,
         oc8051_ram_top1_oc8051_idata_n292, oc8051_ram_top1_oc8051_idata_n291,
         oc8051_ram_top1_oc8051_idata_n290, oc8051_ram_top1_oc8051_idata_n289,
         oc8051_ram_top1_oc8051_idata_n288, oc8051_ram_top1_oc8051_idata_n287,
         oc8051_ram_top1_oc8051_idata_n286, oc8051_ram_top1_oc8051_idata_n285,
         oc8051_ram_top1_oc8051_idata_n284, oc8051_ram_top1_oc8051_idata_n283,
         oc8051_ram_top1_oc8051_idata_n282, oc8051_ram_top1_oc8051_idata_n281,
         oc8051_ram_top1_oc8051_idata_n280, oc8051_ram_top1_oc8051_idata_n279,
         oc8051_ram_top1_oc8051_idata_n278, oc8051_ram_top1_oc8051_idata_n277,
         oc8051_ram_top1_oc8051_idata_n276, oc8051_ram_top1_oc8051_idata_n275,
         oc8051_ram_top1_oc8051_idata_n274, oc8051_ram_top1_oc8051_idata_n273,
         oc8051_ram_top1_oc8051_idata_n272, oc8051_ram_top1_oc8051_idata_n271,
         oc8051_ram_top1_oc8051_idata_n270, oc8051_ram_top1_oc8051_idata_n269,
         oc8051_ram_top1_oc8051_idata_n268, oc8051_ram_top1_oc8051_idata_n267,
         oc8051_ram_top1_oc8051_idata_n266, oc8051_ram_top1_oc8051_idata_n265,
         oc8051_ram_top1_oc8051_idata_n264, oc8051_ram_top1_oc8051_idata_n263,
         oc8051_ram_top1_oc8051_idata_n262, oc8051_ram_top1_oc8051_idata_n261,
         oc8051_ram_top1_oc8051_idata_n260, oc8051_ram_top1_oc8051_idata_n259,
         oc8051_ram_top1_oc8051_idata_n258, oc8051_ram_top1_oc8051_idata_n257,
         oc8051_ram_top1_oc8051_idata_n256, oc8051_ram_top1_oc8051_idata_n255,
         oc8051_ram_top1_oc8051_idata_n254, oc8051_ram_top1_oc8051_idata_n253,
         oc8051_ram_top1_oc8051_idata_n252, oc8051_ram_top1_oc8051_idata_n251,
         oc8051_ram_top1_oc8051_idata_n250, oc8051_ram_top1_oc8051_idata_n249,
         oc8051_ram_top1_oc8051_idata_n248, oc8051_ram_top1_oc8051_idata_n247,
         oc8051_ram_top1_oc8051_idata_n246, oc8051_ram_top1_oc8051_idata_n245,
         oc8051_ram_top1_oc8051_idata_n244, oc8051_ram_top1_oc8051_idata_n243,
         oc8051_ram_top1_oc8051_idata_n242, oc8051_ram_top1_oc8051_idata_n241,
         oc8051_ram_top1_oc8051_idata_n240, oc8051_ram_top1_oc8051_idata_n239,
         oc8051_ram_top1_oc8051_idata_n238, oc8051_ram_top1_oc8051_idata_n237,
         oc8051_ram_top1_oc8051_idata_n236, oc8051_ram_top1_oc8051_idata_n235,
         oc8051_ram_top1_oc8051_idata_n234, oc8051_ram_top1_oc8051_idata_n233,
         oc8051_ram_top1_oc8051_idata_n232, oc8051_ram_top1_oc8051_idata_n231,
         oc8051_ram_top1_oc8051_idata_n230, oc8051_ram_top1_oc8051_idata_n229,
         oc8051_ram_top1_oc8051_idata_n228, oc8051_ram_top1_oc8051_idata_n227,
         oc8051_ram_top1_oc8051_idata_n226, oc8051_ram_top1_oc8051_idata_n225,
         oc8051_ram_top1_oc8051_idata_n224, oc8051_ram_top1_oc8051_idata_n223,
         oc8051_ram_top1_oc8051_idata_n222, oc8051_ram_top1_oc8051_idata_n221,
         oc8051_ram_top1_oc8051_idata_n220, oc8051_ram_top1_oc8051_idata_n219,
         oc8051_ram_top1_oc8051_idata_n218, oc8051_ram_top1_oc8051_idata_n217,
         oc8051_ram_top1_oc8051_idata_n216, oc8051_ram_top1_oc8051_idata_n215,
         oc8051_ram_top1_oc8051_idata_n214, oc8051_ram_top1_oc8051_idata_n213,
         oc8051_ram_top1_oc8051_idata_n212, oc8051_ram_top1_oc8051_idata_n211,
         oc8051_ram_top1_oc8051_idata_n210, oc8051_ram_top1_oc8051_idata_n209,
         oc8051_ram_top1_oc8051_idata_n208, oc8051_ram_top1_oc8051_idata_n207,
         oc8051_ram_top1_oc8051_idata_n206, oc8051_ram_top1_oc8051_idata_n205,
         oc8051_ram_top1_oc8051_idata_n204, oc8051_ram_top1_oc8051_idata_n203,
         oc8051_ram_top1_oc8051_idata_n202, oc8051_ram_top1_oc8051_idata_n201,
         oc8051_ram_top1_oc8051_idata_n200, oc8051_ram_top1_oc8051_idata_n199,
         oc8051_ram_top1_oc8051_idata_n198, oc8051_ram_top1_oc8051_idata_n197,
         oc8051_ram_top1_oc8051_idata_n196, oc8051_ram_top1_oc8051_idata_n195,
         oc8051_ram_top1_oc8051_idata_n194, oc8051_ram_top1_oc8051_idata_n193,
         oc8051_ram_top1_oc8051_idata_n192, oc8051_ram_top1_oc8051_idata_n191,
         oc8051_ram_top1_oc8051_idata_n190, oc8051_ram_top1_oc8051_idata_n189,
         oc8051_ram_top1_oc8051_idata_n188, oc8051_ram_top1_oc8051_idata_n187,
         oc8051_ram_top1_oc8051_idata_n186, oc8051_ram_top1_oc8051_idata_n185,
         oc8051_ram_top1_oc8051_idata_n184, oc8051_ram_top1_oc8051_idata_n183,
         oc8051_ram_top1_oc8051_idata_n182, oc8051_ram_top1_oc8051_idata_n181,
         oc8051_ram_top1_oc8051_idata_n180, oc8051_ram_top1_oc8051_idata_n179,
         oc8051_ram_top1_oc8051_idata_n178, oc8051_ram_top1_oc8051_idata_n177,
         oc8051_ram_top1_oc8051_idata_n176, oc8051_ram_top1_oc8051_idata_n175,
         oc8051_ram_top1_oc8051_idata_n174, oc8051_ram_top1_oc8051_idata_n173,
         oc8051_ram_top1_oc8051_idata_n172, oc8051_ram_top1_oc8051_idata_n171,
         oc8051_ram_top1_oc8051_idata_n170, oc8051_ram_top1_oc8051_idata_n169,
         oc8051_ram_top1_oc8051_idata_n168, oc8051_ram_top1_oc8051_idata_n167,
         oc8051_ram_top1_oc8051_idata_n166, oc8051_ram_top1_oc8051_idata_n165,
         oc8051_ram_top1_oc8051_idata_n164, oc8051_ram_top1_oc8051_idata_n163,
         oc8051_ram_top1_oc8051_idata_n162, oc8051_ram_top1_oc8051_idata_n161,
         oc8051_ram_top1_oc8051_idata_n160, oc8051_ram_top1_oc8051_idata_n159,
         oc8051_ram_top1_oc8051_idata_n158, oc8051_ram_top1_oc8051_idata_n157,
         oc8051_ram_top1_oc8051_idata_n156, oc8051_ram_top1_oc8051_idata_n155,
         oc8051_ram_top1_oc8051_idata_n154, oc8051_ram_top1_oc8051_idata_n153,
         oc8051_ram_top1_oc8051_idata_n152, oc8051_ram_top1_oc8051_idata_n151,
         oc8051_ram_top1_oc8051_idata_n150, oc8051_ram_top1_oc8051_idata_n149,
         oc8051_ram_top1_oc8051_idata_n148, oc8051_ram_top1_oc8051_idata_n147,
         oc8051_ram_top1_oc8051_idata_n146, oc8051_ram_top1_oc8051_idata_n145,
         oc8051_ram_top1_oc8051_idata_n144, oc8051_ram_top1_oc8051_idata_n143,
         oc8051_ram_top1_oc8051_idata_n142, oc8051_ram_top1_oc8051_idata_n141,
         oc8051_ram_top1_oc8051_idata_n140, oc8051_ram_top1_oc8051_idata_n139,
         oc8051_ram_top1_oc8051_idata_n138, oc8051_ram_top1_oc8051_idata_n137,
         oc8051_ram_top1_oc8051_idata_n136, oc8051_ram_top1_oc8051_idata_n135,
         oc8051_ram_top1_oc8051_idata_n134, oc8051_ram_top1_oc8051_idata_n133,
         oc8051_ram_top1_oc8051_idata_n132, oc8051_ram_top1_oc8051_idata_n131,
         oc8051_ram_top1_oc8051_idata_n130, oc8051_ram_top1_oc8051_idata_n129,
         oc8051_ram_top1_oc8051_idata_n128, oc8051_ram_top1_oc8051_idata_n127,
         oc8051_ram_top1_oc8051_idata_n126, oc8051_ram_top1_oc8051_idata_n125,
         oc8051_ram_top1_oc8051_idata_n124, oc8051_ram_top1_oc8051_idata_n123,
         oc8051_ram_top1_oc8051_idata_n122, oc8051_ram_top1_oc8051_idata_n121,
         oc8051_ram_top1_oc8051_idata_n120, oc8051_ram_top1_oc8051_idata_n119,
         oc8051_ram_top1_oc8051_idata_n118, oc8051_ram_top1_oc8051_idata_n117,
         oc8051_ram_top1_oc8051_idata_n116, oc8051_ram_top1_oc8051_idata_n115,
         oc8051_ram_top1_oc8051_idata_n114, oc8051_ram_top1_oc8051_idata_n113,
         oc8051_ram_top1_oc8051_idata_n112, oc8051_ram_top1_oc8051_idata_n111,
         oc8051_ram_top1_oc8051_idata_n110, oc8051_ram_top1_oc8051_idata_n109,
         oc8051_ram_top1_oc8051_idata_n108, oc8051_ram_top1_oc8051_idata_n107,
         oc8051_ram_top1_oc8051_idata_n106, oc8051_ram_top1_oc8051_idata_n105,
         oc8051_ram_top1_oc8051_idata_n104, oc8051_ram_top1_oc8051_idata_n103,
         oc8051_ram_top1_oc8051_idata_n102, oc8051_ram_top1_oc8051_idata_n101,
         oc8051_ram_top1_oc8051_idata_n100, oc8051_ram_top1_oc8051_idata_n99,
         oc8051_ram_top1_oc8051_idata_n98, oc8051_ram_top1_oc8051_idata_n97,
         oc8051_ram_top1_oc8051_idata_n96, oc8051_ram_top1_oc8051_idata_n95,
         oc8051_ram_top1_oc8051_idata_n94, oc8051_ram_top1_oc8051_idata_n93,
         oc8051_ram_top1_oc8051_idata_n92, oc8051_ram_top1_oc8051_idata_n91,
         oc8051_ram_top1_oc8051_idata_n90, oc8051_ram_top1_oc8051_idata_n89,
         oc8051_ram_top1_oc8051_idata_n88, oc8051_ram_top1_oc8051_idata_n87,
         oc8051_ram_top1_oc8051_idata_n86, oc8051_ram_top1_oc8051_idata_n85,
         oc8051_ram_top1_oc8051_idata_n84, oc8051_ram_top1_oc8051_idata_n83,
         oc8051_ram_top1_oc8051_idata_n82, oc8051_ram_top1_oc8051_idata_n81,
         oc8051_ram_top1_oc8051_idata_n80, oc8051_ram_top1_oc8051_idata_n79,
         oc8051_ram_top1_oc8051_idata_n78, oc8051_ram_top1_oc8051_idata_n77,
         oc8051_ram_top1_oc8051_idata_n76, oc8051_ram_top1_oc8051_idata_n75,
         oc8051_ram_top1_oc8051_idata_n74, oc8051_ram_top1_oc8051_idata_n73,
         oc8051_ram_top1_oc8051_idata_n72, oc8051_ram_top1_oc8051_idata_n71,
         oc8051_ram_top1_oc8051_idata_n70, oc8051_ram_top1_oc8051_idata_n69,
         oc8051_ram_top1_oc8051_idata_n68, oc8051_ram_top1_oc8051_idata_n67,
         oc8051_ram_top1_oc8051_idata_n66, oc8051_ram_top1_oc8051_idata_n65,
         oc8051_ram_top1_oc8051_idata_n64, oc8051_ram_top1_oc8051_idata_n63,
         oc8051_ram_top1_oc8051_idata_n62, oc8051_ram_top1_oc8051_idata_n61,
         oc8051_ram_top1_oc8051_idata_n60, oc8051_ram_top1_oc8051_idata_n59,
         oc8051_ram_top1_oc8051_idata_n58, oc8051_ram_top1_oc8051_idata_n57,
         oc8051_ram_top1_oc8051_idata_n56, oc8051_ram_top1_oc8051_idata_n55,
         oc8051_ram_top1_oc8051_idata_n54, oc8051_ram_top1_oc8051_idata_n53,
         oc8051_ram_top1_oc8051_idata_n52, oc8051_ram_top1_oc8051_idata_n51,
         oc8051_ram_top1_oc8051_idata_n50, oc8051_ram_top1_oc8051_idata_n49,
         oc8051_ram_top1_oc8051_idata_n48, oc8051_ram_top1_oc8051_idata_n47,
         oc8051_ram_top1_oc8051_idata_n46, oc8051_ram_top1_oc8051_idata_n45,
         oc8051_ram_top1_oc8051_idata_n44, oc8051_ram_top1_oc8051_idata_n43,
         oc8051_ram_top1_oc8051_idata_n42, oc8051_ram_top1_oc8051_idata_n41,
         oc8051_ram_top1_oc8051_idata_n40, oc8051_ram_top1_oc8051_idata_n39,
         oc8051_ram_top1_oc8051_idata_n38, oc8051_ram_top1_oc8051_idata_n37,
         oc8051_ram_top1_oc8051_idata_n36, oc8051_ram_top1_oc8051_idata_n35,
         oc8051_ram_top1_oc8051_idata_n34, oc8051_ram_top1_oc8051_idata_n33,
         oc8051_ram_top1_oc8051_idata_n32, oc8051_ram_top1_oc8051_idata_n31,
         oc8051_ram_top1_oc8051_idata_n30, oc8051_ram_top1_oc8051_idata_n29,
         oc8051_ram_top1_oc8051_idata_n28, oc8051_ram_top1_oc8051_idata_n27,
         oc8051_ram_top1_oc8051_idata_n26, oc8051_ram_top1_oc8051_idata_n25,
         oc8051_ram_top1_oc8051_idata_n24, oc8051_ram_top1_oc8051_idata_n23,
         oc8051_ram_top1_oc8051_idata_n22, oc8051_ram_top1_oc8051_idata_n21,
         oc8051_ram_top1_oc8051_idata_n20, oc8051_ram_top1_oc8051_idata_n19,
         oc8051_ram_top1_oc8051_idata_n18, oc8051_ram_top1_oc8051_idata_n17,
         oc8051_ram_top1_oc8051_idata_n16, oc8051_ram_top1_oc8051_idata_n15,
         oc8051_ram_top1_oc8051_idata_n14, oc8051_ram_top1_oc8051_idata_n13,
         oc8051_ram_top1_oc8051_idata_n12, oc8051_ram_top1_oc8051_idata_n11,
         oc8051_ram_top1_oc8051_idata_n10, oc8051_ram_top1_oc8051_idata_n9,
         oc8051_ram_top1_oc8051_idata_n8, oc8051_ram_top1_oc8051_idata_n7,
         oc8051_ram_top1_oc8051_idata_n6, oc8051_ram_top1_oc8051_idata_n5,
         oc8051_ram_top1_oc8051_idata_n4,
         oc8051_ram_top1_oc8051_idata_buff_127__0_,
         oc8051_ram_top1_oc8051_idata_buff_127__1_,
         oc8051_ram_top1_oc8051_idata_buff_127__2_,
         oc8051_ram_top1_oc8051_idata_buff_127__3_,
         oc8051_ram_top1_oc8051_idata_buff_127__4_,
         oc8051_ram_top1_oc8051_idata_buff_127__5_,
         oc8051_ram_top1_oc8051_idata_buff_127__6_,
         oc8051_ram_top1_oc8051_idata_buff_127__7_,
         oc8051_ram_top1_oc8051_idata_buff_126__0_,
         oc8051_ram_top1_oc8051_idata_buff_126__1_,
         oc8051_ram_top1_oc8051_idata_buff_126__2_,
         oc8051_ram_top1_oc8051_idata_buff_126__3_,
         oc8051_ram_top1_oc8051_idata_buff_126__4_,
         oc8051_ram_top1_oc8051_idata_buff_126__5_,
         oc8051_ram_top1_oc8051_idata_buff_126__6_,
         oc8051_ram_top1_oc8051_idata_buff_126__7_,
         oc8051_ram_top1_oc8051_idata_buff_125__0_,
         oc8051_ram_top1_oc8051_idata_buff_125__1_,
         oc8051_ram_top1_oc8051_idata_buff_125__2_,
         oc8051_ram_top1_oc8051_idata_buff_125__3_,
         oc8051_ram_top1_oc8051_idata_buff_125__4_,
         oc8051_ram_top1_oc8051_idata_buff_125__5_,
         oc8051_ram_top1_oc8051_idata_buff_125__6_,
         oc8051_ram_top1_oc8051_idata_buff_125__7_,
         oc8051_ram_top1_oc8051_idata_buff_124__0_,
         oc8051_ram_top1_oc8051_idata_buff_124__1_,
         oc8051_ram_top1_oc8051_idata_buff_124__2_,
         oc8051_ram_top1_oc8051_idata_buff_124__3_,
         oc8051_ram_top1_oc8051_idata_buff_124__4_,
         oc8051_ram_top1_oc8051_idata_buff_124__5_,
         oc8051_ram_top1_oc8051_idata_buff_124__6_,
         oc8051_ram_top1_oc8051_idata_buff_124__7_,
         oc8051_ram_top1_oc8051_idata_buff_123__0_,
         oc8051_ram_top1_oc8051_idata_buff_123__1_,
         oc8051_ram_top1_oc8051_idata_buff_123__2_,
         oc8051_ram_top1_oc8051_idata_buff_123__3_,
         oc8051_ram_top1_oc8051_idata_buff_123__4_,
         oc8051_ram_top1_oc8051_idata_buff_123__5_,
         oc8051_ram_top1_oc8051_idata_buff_123__6_,
         oc8051_ram_top1_oc8051_idata_buff_123__7_,
         oc8051_ram_top1_oc8051_idata_buff_122__0_,
         oc8051_ram_top1_oc8051_idata_buff_122__1_,
         oc8051_ram_top1_oc8051_idata_buff_122__2_,
         oc8051_ram_top1_oc8051_idata_buff_122__3_,
         oc8051_ram_top1_oc8051_idata_buff_122__4_,
         oc8051_ram_top1_oc8051_idata_buff_122__5_,
         oc8051_ram_top1_oc8051_idata_buff_122__6_,
         oc8051_ram_top1_oc8051_idata_buff_122__7_,
         oc8051_ram_top1_oc8051_idata_buff_121__0_,
         oc8051_ram_top1_oc8051_idata_buff_121__1_,
         oc8051_ram_top1_oc8051_idata_buff_121__2_,
         oc8051_ram_top1_oc8051_idata_buff_121__3_,
         oc8051_ram_top1_oc8051_idata_buff_121__4_,
         oc8051_ram_top1_oc8051_idata_buff_121__5_,
         oc8051_ram_top1_oc8051_idata_buff_121__6_,
         oc8051_ram_top1_oc8051_idata_buff_121__7_,
         oc8051_ram_top1_oc8051_idata_buff_120__0_,
         oc8051_ram_top1_oc8051_idata_buff_120__1_,
         oc8051_ram_top1_oc8051_idata_buff_120__2_,
         oc8051_ram_top1_oc8051_idata_buff_120__3_,
         oc8051_ram_top1_oc8051_idata_buff_120__4_,
         oc8051_ram_top1_oc8051_idata_buff_120__5_,
         oc8051_ram_top1_oc8051_idata_buff_120__6_,
         oc8051_ram_top1_oc8051_idata_buff_120__7_,
         oc8051_ram_top1_oc8051_idata_buff_117__0_,
         oc8051_ram_top1_oc8051_idata_buff_117__1_,
         oc8051_ram_top1_oc8051_idata_buff_117__2_,
         oc8051_ram_top1_oc8051_idata_buff_117__3_,
         oc8051_ram_top1_oc8051_idata_buff_117__4_,
         oc8051_ram_top1_oc8051_idata_buff_117__5_,
         oc8051_ram_top1_oc8051_idata_buff_117__6_,
         oc8051_ram_top1_oc8051_idata_buff_117__7_,
         oc8051_ram_top1_oc8051_idata_buff_116__0_,
         oc8051_ram_top1_oc8051_idata_buff_116__1_,
         oc8051_ram_top1_oc8051_idata_buff_116__2_,
         oc8051_ram_top1_oc8051_idata_buff_116__3_,
         oc8051_ram_top1_oc8051_idata_buff_116__4_,
         oc8051_ram_top1_oc8051_idata_buff_116__5_,
         oc8051_ram_top1_oc8051_idata_buff_116__6_,
         oc8051_ram_top1_oc8051_idata_buff_116__7_,
         oc8051_ram_top1_oc8051_idata_buff_113__0_,
         oc8051_ram_top1_oc8051_idata_buff_113__1_,
         oc8051_ram_top1_oc8051_idata_buff_113__2_,
         oc8051_ram_top1_oc8051_idata_buff_113__3_,
         oc8051_ram_top1_oc8051_idata_buff_113__4_,
         oc8051_ram_top1_oc8051_idata_buff_113__5_,
         oc8051_ram_top1_oc8051_idata_buff_113__6_,
         oc8051_ram_top1_oc8051_idata_buff_113__7_,
         oc8051_ram_top1_oc8051_idata_buff_112__0_,
         oc8051_ram_top1_oc8051_idata_buff_112__1_,
         oc8051_ram_top1_oc8051_idata_buff_112__2_,
         oc8051_ram_top1_oc8051_idata_buff_112__3_,
         oc8051_ram_top1_oc8051_idata_buff_112__4_,
         oc8051_ram_top1_oc8051_idata_buff_112__5_,
         oc8051_ram_top1_oc8051_idata_buff_112__6_,
         oc8051_ram_top1_oc8051_idata_buff_112__7_,
         oc8051_ram_top1_oc8051_idata_buff_111__0_,
         oc8051_ram_top1_oc8051_idata_buff_111__1_,
         oc8051_ram_top1_oc8051_idata_buff_111__2_,
         oc8051_ram_top1_oc8051_idata_buff_111__3_,
         oc8051_ram_top1_oc8051_idata_buff_111__4_,
         oc8051_ram_top1_oc8051_idata_buff_111__5_,
         oc8051_ram_top1_oc8051_idata_buff_111__6_,
         oc8051_ram_top1_oc8051_idata_buff_111__7_,
         oc8051_ram_top1_oc8051_idata_buff_110__0_,
         oc8051_ram_top1_oc8051_idata_buff_110__1_,
         oc8051_ram_top1_oc8051_idata_buff_110__2_,
         oc8051_ram_top1_oc8051_idata_buff_110__3_,
         oc8051_ram_top1_oc8051_idata_buff_110__4_,
         oc8051_ram_top1_oc8051_idata_buff_110__5_,
         oc8051_ram_top1_oc8051_idata_buff_110__6_,
         oc8051_ram_top1_oc8051_idata_buff_110__7_,
         oc8051_ram_top1_oc8051_idata_buff_109__0_,
         oc8051_ram_top1_oc8051_idata_buff_109__1_,
         oc8051_ram_top1_oc8051_idata_buff_109__2_,
         oc8051_ram_top1_oc8051_idata_buff_109__3_,
         oc8051_ram_top1_oc8051_idata_buff_109__4_,
         oc8051_ram_top1_oc8051_idata_buff_109__5_,
         oc8051_ram_top1_oc8051_idata_buff_109__6_,
         oc8051_ram_top1_oc8051_idata_buff_109__7_,
         oc8051_ram_top1_oc8051_idata_buff_108__0_,
         oc8051_ram_top1_oc8051_idata_buff_108__1_,
         oc8051_ram_top1_oc8051_idata_buff_108__2_,
         oc8051_ram_top1_oc8051_idata_buff_108__3_,
         oc8051_ram_top1_oc8051_idata_buff_108__4_,
         oc8051_ram_top1_oc8051_idata_buff_108__5_,
         oc8051_ram_top1_oc8051_idata_buff_108__6_,
         oc8051_ram_top1_oc8051_idata_buff_108__7_,
         oc8051_ram_top1_oc8051_idata_buff_107__0_,
         oc8051_ram_top1_oc8051_idata_buff_107__1_,
         oc8051_ram_top1_oc8051_idata_buff_107__2_,
         oc8051_ram_top1_oc8051_idata_buff_107__3_,
         oc8051_ram_top1_oc8051_idata_buff_107__4_,
         oc8051_ram_top1_oc8051_idata_buff_107__5_,
         oc8051_ram_top1_oc8051_idata_buff_107__6_,
         oc8051_ram_top1_oc8051_idata_buff_107__7_,
         oc8051_ram_top1_oc8051_idata_buff_106__0_,
         oc8051_ram_top1_oc8051_idata_buff_106__1_,
         oc8051_ram_top1_oc8051_idata_buff_106__2_,
         oc8051_ram_top1_oc8051_idata_buff_106__3_,
         oc8051_ram_top1_oc8051_idata_buff_106__4_,
         oc8051_ram_top1_oc8051_idata_buff_106__5_,
         oc8051_ram_top1_oc8051_idata_buff_106__6_,
         oc8051_ram_top1_oc8051_idata_buff_106__7_,
         oc8051_ram_top1_oc8051_idata_buff_105__0_,
         oc8051_ram_top1_oc8051_idata_buff_105__1_,
         oc8051_ram_top1_oc8051_idata_buff_105__2_,
         oc8051_ram_top1_oc8051_idata_buff_105__3_,
         oc8051_ram_top1_oc8051_idata_buff_105__4_,
         oc8051_ram_top1_oc8051_idata_buff_105__5_,
         oc8051_ram_top1_oc8051_idata_buff_105__6_,
         oc8051_ram_top1_oc8051_idata_buff_105__7_,
         oc8051_ram_top1_oc8051_idata_buff_104__0_,
         oc8051_ram_top1_oc8051_idata_buff_104__1_,
         oc8051_ram_top1_oc8051_idata_buff_104__2_,
         oc8051_ram_top1_oc8051_idata_buff_104__3_,
         oc8051_ram_top1_oc8051_idata_buff_104__4_,
         oc8051_ram_top1_oc8051_idata_buff_104__5_,
         oc8051_ram_top1_oc8051_idata_buff_104__6_,
         oc8051_ram_top1_oc8051_idata_buff_104__7_,
         oc8051_ram_top1_oc8051_idata_buff_103__0_,
         oc8051_ram_top1_oc8051_idata_buff_103__1_,
         oc8051_ram_top1_oc8051_idata_buff_103__2_,
         oc8051_ram_top1_oc8051_idata_buff_103__3_,
         oc8051_ram_top1_oc8051_idata_buff_103__4_,
         oc8051_ram_top1_oc8051_idata_buff_103__5_,
         oc8051_ram_top1_oc8051_idata_buff_103__6_,
         oc8051_ram_top1_oc8051_idata_buff_103__7_,
         oc8051_ram_top1_oc8051_idata_buff_102__0_,
         oc8051_ram_top1_oc8051_idata_buff_102__1_,
         oc8051_ram_top1_oc8051_idata_buff_102__2_,
         oc8051_ram_top1_oc8051_idata_buff_102__3_,
         oc8051_ram_top1_oc8051_idata_buff_102__4_,
         oc8051_ram_top1_oc8051_idata_buff_102__5_,
         oc8051_ram_top1_oc8051_idata_buff_102__6_,
         oc8051_ram_top1_oc8051_idata_buff_102__7_,
         oc8051_ram_top1_oc8051_idata_buff_99__0_,
         oc8051_ram_top1_oc8051_idata_buff_99__1_,
         oc8051_ram_top1_oc8051_idata_buff_99__2_,
         oc8051_ram_top1_oc8051_idata_buff_99__3_,
         oc8051_ram_top1_oc8051_idata_buff_99__4_,
         oc8051_ram_top1_oc8051_idata_buff_99__5_,
         oc8051_ram_top1_oc8051_idata_buff_99__6_,
         oc8051_ram_top1_oc8051_idata_buff_99__7_,
         oc8051_ram_top1_oc8051_idata_buff_98__0_,
         oc8051_ram_top1_oc8051_idata_buff_98__1_,
         oc8051_ram_top1_oc8051_idata_buff_98__2_,
         oc8051_ram_top1_oc8051_idata_buff_98__3_,
         oc8051_ram_top1_oc8051_idata_buff_98__4_,
         oc8051_ram_top1_oc8051_idata_buff_98__5_,
         oc8051_ram_top1_oc8051_idata_buff_98__6_,
         oc8051_ram_top1_oc8051_idata_buff_98__7_,
         oc8051_ram_top1_oc8051_idata_buff_95__0_,
         oc8051_ram_top1_oc8051_idata_buff_95__1_,
         oc8051_ram_top1_oc8051_idata_buff_95__2_,
         oc8051_ram_top1_oc8051_idata_buff_95__3_,
         oc8051_ram_top1_oc8051_idata_buff_95__4_,
         oc8051_ram_top1_oc8051_idata_buff_95__5_,
         oc8051_ram_top1_oc8051_idata_buff_95__6_,
         oc8051_ram_top1_oc8051_idata_buff_95__7_,
         oc8051_ram_top1_oc8051_idata_buff_94__0_,
         oc8051_ram_top1_oc8051_idata_buff_94__1_,
         oc8051_ram_top1_oc8051_idata_buff_94__2_,
         oc8051_ram_top1_oc8051_idata_buff_94__3_,
         oc8051_ram_top1_oc8051_idata_buff_94__4_,
         oc8051_ram_top1_oc8051_idata_buff_94__5_,
         oc8051_ram_top1_oc8051_idata_buff_94__6_,
         oc8051_ram_top1_oc8051_idata_buff_94__7_,
         oc8051_ram_top1_oc8051_idata_buff_93__0_,
         oc8051_ram_top1_oc8051_idata_buff_93__1_,
         oc8051_ram_top1_oc8051_idata_buff_93__2_,
         oc8051_ram_top1_oc8051_idata_buff_93__3_,
         oc8051_ram_top1_oc8051_idata_buff_93__4_,
         oc8051_ram_top1_oc8051_idata_buff_93__5_,
         oc8051_ram_top1_oc8051_idata_buff_93__6_,
         oc8051_ram_top1_oc8051_idata_buff_93__7_,
         oc8051_ram_top1_oc8051_idata_buff_92__0_,
         oc8051_ram_top1_oc8051_idata_buff_92__1_,
         oc8051_ram_top1_oc8051_idata_buff_92__2_,
         oc8051_ram_top1_oc8051_idata_buff_92__3_,
         oc8051_ram_top1_oc8051_idata_buff_92__4_,
         oc8051_ram_top1_oc8051_idata_buff_92__5_,
         oc8051_ram_top1_oc8051_idata_buff_92__6_,
         oc8051_ram_top1_oc8051_idata_buff_92__7_,
         oc8051_ram_top1_oc8051_idata_buff_91__0_,
         oc8051_ram_top1_oc8051_idata_buff_91__1_,
         oc8051_ram_top1_oc8051_idata_buff_91__2_,
         oc8051_ram_top1_oc8051_idata_buff_91__3_,
         oc8051_ram_top1_oc8051_idata_buff_91__4_,
         oc8051_ram_top1_oc8051_idata_buff_91__5_,
         oc8051_ram_top1_oc8051_idata_buff_91__6_,
         oc8051_ram_top1_oc8051_idata_buff_91__7_,
         oc8051_ram_top1_oc8051_idata_buff_90__0_,
         oc8051_ram_top1_oc8051_idata_buff_90__1_,
         oc8051_ram_top1_oc8051_idata_buff_90__2_,
         oc8051_ram_top1_oc8051_idata_buff_90__3_,
         oc8051_ram_top1_oc8051_idata_buff_90__4_,
         oc8051_ram_top1_oc8051_idata_buff_90__5_,
         oc8051_ram_top1_oc8051_idata_buff_90__6_,
         oc8051_ram_top1_oc8051_idata_buff_90__7_,
         oc8051_ram_top1_oc8051_idata_buff_89__0_,
         oc8051_ram_top1_oc8051_idata_buff_89__1_,
         oc8051_ram_top1_oc8051_idata_buff_89__2_,
         oc8051_ram_top1_oc8051_idata_buff_89__3_,
         oc8051_ram_top1_oc8051_idata_buff_89__4_,
         oc8051_ram_top1_oc8051_idata_buff_89__5_,
         oc8051_ram_top1_oc8051_idata_buff_89__6_,
         oc8051_ram_top1_oc8051_idata_buff_89__7_,
         oc8051_ram_top1_oc8051_idata_buff_88__0_,
         oc8051_ram_top1_oc8051_idata_buff_88__1_,
         oc8051_ram_top1_oc8051_idata_buff_88__2_,
         oc8051_ram_top1_oc8051_idata_buff_88__3_,
         oc8051_ram_top1_oc8051_idata_buff_88__4_,
         oc8051_ram_top1_oc8051_idata_buff_88__5_,
         oc8051_ram_top1_oc8051_idata_buff_88__6_,
         oc8051_ram_top1_oc8051_idata_buff_88__7_,
         oc8051_ram_top1_oc8051_idata_buff_87__0_,
         oc8051_ram_top1_oc8051_idata_buff_87__1_,
         oc8051_ram_top1_oc8051_idata_buff_87__2_,
         oc8051_ram_top1_oc8051_idata_buff_87__3_,
         oc8051_ram_top1_oc8051_idata_buff_87__4_,
         oc8051_ram_top1_oc8051_idata_buff_87__5_,
         oc8051_ram_top1_oc8051_idata_buff_87__6_,
         oc8051_ram_top1_oc8051_idata_buff_87__7_,
         oc8051_ram_top1_oc8051_idata_buff_86__0_,
         oc8051_ram_top1_oc8051_idata_buff_86__1_,
         oc8051_ram_top1_oc8051_idata_buff_86__2_,
         oc8051_ram_top1_oc8051_idata_buff_86__3_,
         oc8051_ram_top1_oc8051_idata_buff_86__4_,
         oc8051_ram_top1_oc8051_idata_buff_86__5_,
         oc8051_ram_top1_oc8051_idata_buff_86__6_,
         oc8051_ram_top1_oc8051_idata_buff_86__7_,
         oc8051_ram_top1_oc8051_idata_buff_85__0_,
         oc8051_ram_top1_oc8051_idata_buff_85__1_,
         oc8051_ram_top1_oc8051_idata_buff_85__2_,
         oc8051_ram_top1_oc8051_idata_buff_85__3_,
         oc8051_ram_top1_oc8051_idata_buff_85__4_,
         oc8051_ram_top1_oc8051_idata_buff_85__5_,
         oc8051_ram_top1_oc8051_idata_buff_85__6_,
         oc8051_ram_top1_oc8051_idata_buff_85__7_,
         oc8051_ram_top1_oc8051_idata_buff_84__0_,
         oc8051_ram_top1_oc8051_idata_buff_84__1_,
         oc8051_ram_top1_oc8051_idata_buff_84__2_,
         oc8051_ram_top1_oc8051_idata_buff_84__3_,
         oc8051_ram_top1_oc8051_idata_buff_84__4_,
         oc8051_ram_top1_oc8051_idata_buff_84__5_,
         oc8051_ram_top1_oc8051_idata_buff_84__6_,
         oc8051_ram_top1_oc8051_idata_buff_84__7_,
         oc8051_ram_top1_oc8051_idata_buff_83__0_,
         oc8051_ram_top1_oc8051_idata_buff_83__1_,
         oc8051_ram_top1_oc8051_idata_buff_83__2_,
         oc8051_ram_top1_oc8051_idata_buff_83__3_,
         oc8051_ram_top1_oc8051_idata_buff_83__4_,
         oc8051_ram_top1_oc8051_idata_buff_83__5_,
         oc8051_ram_top1_oc8051_idata_buff_83__6_,
         oc8051_ram_top1_oc8051_idata_buff_83__7_,
         oc8051_ram_top1_oc8051_idata_buff_82__0_,
         oc8051_ram_top1_oc8051_idata_buff_82__1_,
         oc8051_ram_top1_oc8051_idata_buff_82__2_,
         oc8051_ram_top1_oc8051_idata_buff_82__3_,
         oc8051_ram_top1_oc8051_idata_buff_82__4_,
         oc8051_ram_top1_oc8051_idata_buff_82__5_,
         oc8051_ram_top1_oc8051_idata_buff_82__6_,
         oc8051_ram_top1_oc8051_idata_buff_82__7_,
         oc8051_ram_top1_oc8051_idata_buff_81__0_,
         oc8051_ram_top1_oc8051_idata_buff_81__1_,
         oc8051_ram_top1_oc8051_idata_buff_81__2_,
         oc8051_ram_top1_oc8051_idata_buff_81__3_,
         oc8051_ram_top1_oc8051_idata_buff_81__4_,
         oc8051_ram_top1_oc8051_idata_buff_81__5_,
         oc8051_ram_top1_oc8051_idata_buff_81__6_,
         oc8051_ram_top1_oc8051_idata_buff_81__7_,
         oc8051_ram_top1_oc8051_idata_buff_80__0_,
         oc8051_ram_top1_oc8051_idata_buff_80__1_,
         oc8051_ram_top1_oc8051_idata_buff_80__2_,
         oc8051_ram_top1_oc8051_idata_buff_80__3_,
         oc8051_ram_top1_oc8051_idata_buff_80__4_,
         oc8051_ram_top1_oc8051_idata_buff_80__5_,
         oc8051_ram_top1_oc8051_idata_buff_80__6_,
         oc8051_ram_top1_oc8051_idata_buff_80__7_,
         oc8051_ram_top1_oc8051_idata_buff_77__0_,
         oc8051_ram_top1_oc8051_idata_buff_77__1_,
         oc8051_ram_top1_oc8051_idata_buff_77__2_,
         oc8051_ram_top1_oc8051_idata_buff_77__3_,
         oc8051_ram_top1_oc8051_idata_buff_77__4_,
         oc8051_ram_top1_oc8051_idata_buff_77__5_,
         oc8051_ram_top1_oc8051_idata_buff_77__6_,
         oc8051_ram_top1_oc8051_idata_buff_77__7_,
         oc8051_ram_top1_oc8051_idata_buff_76__0_,
         oc8051_ram_top1_oc8051_idata_buff_76__1_,
         oc8051_ram_top1_oc8051_idata_buff_76__2_,
         oc8051_ram_top1_oc8051_idata_buff_76__3_,
         oc8051_ram_top1_oc8051_idata_buff_76__4_,
         oc8051_ram_top1_oc8051_idata_buff_76__5_,
         oc8051_ram_top1_oc8051_idata_buff_76__6_,
         oc8051_ram_top1_oc8051_idata_buff_76__7_,
         oc8051_ram_top1_oc8051_idata_buff_75__0_,
         oc8051_ram_top1_oc8051_idata_buff_75__1_,
         oc8051_ram_top1_oc8051_idata_buff_75__2_,
         oc8051_ram_top1_oc8051_idata_buff_75__3_,
         oc8051_ram_top1_oc8051_idata_buff_75__4_,
         oc8051_ram_top1_oc8051_idata_buff_75__5_,
         oc8051_ram_top1_oc8051_idata_buff_75__6_,
         oc8051_ram_top1_oc8051_idata_buff_75__7_,
         oc8051_ram_top1_oc8051_idata_buff_74__0_,
         oc8051_ram_top1_oc8051_idata_buff_74__1_,
         oc8051_ram_top1_oc8051_idata_buff_74__2_,
         oc8051_ram_top1_oc8051_idata_buff_74__3_,
         oc8051_ram_top1_oc8051_idata_buff_74__4_,
         oc8051_ram_top1_oc8051_idata_buff_74__5_,
         oc8051_ram_top1_oc8051_idata_buff_74__6_,
         oc8051_ram_top1_oc8051_idata_buff_74__7_,
         oc8051_ram_top1_oc8051_idata_buff_71__0_,
         oc8051_ram_top1_oc8051_idata_buff_71__1_,
         oc8051_ram_top1_oc8051_idata_buff_71__2_,
         oc8051_ram_top1_oc8051_idata_buff_71__3_,
         oc8051_ram_top1_oc8051_idata_buff_71__4_,
         oc8051_ram_top1_oc8051_idata_buff_71__5_,
         oc8051_ram_top1_oc8051_idata_buff_71__6_,
         oc8051_ram_top1_oc8051_idata_buff_71__7_,
         oc8051_ram_top1_oc8051_idata_buff_70__0_,
         oc8051_ram_top1_oc8051_idata_buff_70__1_,
         oc8051_ram_top1_oc8051_idata_buff_70__2_,
         oc8051_ram_top1_oc8051_idata_buff_70__3_,
         oc8051_ram_top1_oc8051_idata_buff_70__4_,
         oc8051_ram_top1_oc8051_idata_buff_70__5_,
         oc8051_ram_top1_oc8051_idata_buff_70__6_,
         oc8051_ram_top1_oc8051_idata_buff_70__7_,
         oc8051_ram_top1_oc8051_idata_buff_67__0_,
         oc8051_ram_top1_oc8051_idata_buff_67__1_,
         oc8051_ram_top1_oc8051_idata_buff_67__2_,
         oc8051_ram_top1_oc8051_idata_buff_67__3_,
         oc8051_ram_top1_oc8051_idata_buff_67__4_,
         oc8051_ram_top1_oc8051_idata_buff_67__5_,
         oc8051_ram_top1_oc8051_idata_buff_67__6_,
         oc8051_ram_top1_oc8051_idata_buff_67__7_,
         oc8051_ram_top1_oc8051_idata_buff_66__0_,
         oc8051_ram_top1_oc8051_idata_buff_66__1_,
         oc8051_ram_top1_oc8051_idata_buff_66__2_,
         oc8051_ram_top1_oc8051_idata_buff_66__3_,
         oc8051_ram_top1_oc8051_idata_buff_66__4_,
         oc8051_ram_top1_oc8051_idata_buff_66__5_,
         oc8051_ram_top1_oc8051_idata_buff_66__6_,
         oc8051_ram_top1_oc8051_idata_buff_66__7_,
         oc8051_ram_top1_oc8051_idata_buff_191__0_,
         oc8051_ram_top1_oc8051_idata_buff_191__1_,
         oc8051_ram_top1_oc8051_idata_buff_191__2_,
         oc8051_ram_top1_oc8051_idata_buff_191__3_,
         oc8051_ram_top1_oc8051_idata_buff_191__4_,
         oc8051_ram_top1_oc8051_idata_buff_191__5_,
         oc8051_ram_top1_oc8051_idata_buff_191__6_,
         oc8051_ram_top1_oc8051_idata_buff_191__7_,
         oc8051_ram_top1_oc8051_idata_buff_190__0_,
         oc8051_ram_top1_oc8051_idata_buff_190__1_,
         oc8051_ram_top1_oc8051_idata_buff_190__2_,
         oc8051_ram_top1_oc8051_idata_buff_190__3_,
         oc8051_ram_top1_oc8051_idata_buff_190__4_,
         oc8051_ram_top1_oc8051_idata_buff_190__5_,
         oc8051_ram_top1_oc8051_idata_buff_190__6_,
         oc8051_ram_top1_oc8051_idata_buff_190__7_,
         oc8051_ram_top1_oc8051_idata_buff_189__0_,
         oc8051_ram_top1_oc8051_idata_buff_189__1_,
         oc8051_ram_top1_oc8051_idata_buff_189__2_,
         oc8051_ram_top1_oc8051_idata_buff_189__3_,
         oc8051_ram_top1_oc8051_idata_buff_189__4_,
         oc8051_ram_top1_oc8051_idata_buff_189__5_,
         oc8051_ram_top1_oc8051_idata_buff_189__6_,
         oc8051_ram_top1_oc8051_idata_buff_189__7_,
         oc8051_ram_top1_oc8051_idata_buff_188__0_,
         oc8051_ram_top1_oc8051_idata_buff_188__1_,
         oc8051_ram_top1_oc8051_idata_buff_188__2_,
         oc8051_ram_top1_oc8051_idata_buff_188__3_,
         oc8051_ram_top1_oc8051_idata_buff_188__4_,
         oc8051_ram_top1_oc8051_idata_buff_188__5_,
         oc8051_ram_top1_oc8051_idata_buff_188__6_,
         oc8051_ram_top1_oc8051_idata_buff_188__7_,
         oc8051_ram_top1_oc8051_idata_buff_187__0_,
         oc8051_ram_top1_oc8051_idata_buff_187__1_,
         oc8051_ram_top1_oc8051_idata_buff_187__2_,
         oc8051_ram_top1_oc8051_idata_buff_187__3_,
         oc8051_ram_top1_oc8051_idata_buff_187__4_,
         oc8051_ram_top1_oc8051_idata_buff_187__5_,
         oc8051_ram_top1_oc8051_idata_buff_187__6_,
         oc8051_ram_top1_oc8051_idata_buff_187__7_,
         oc8051_ram_top1_oc8051_idata_buff_186__0_,
         oc8051_ram_top1_oc8051_idata_buff_186__1_,
         oc8051_ram_top1_oc8051_idata_buff_186__2_,
         oc8051_ram_top1_oc8051_idata_buff_186__3_,
         oc8051_ram_top1_oc8051_idata_buff_186__4_,
         oc8051_ram_top1_oc8051_idata_buff_186__5_,
         oc8051_ram_top1_oc8051_idata_buff_186__6_,
         oc8051_ram_top1_oc8051_idata_buff_186__7_,
         oc8051_ram_top1_oc8051_idata_buff_185__0_,
         oc8051_ram_top1_oc8051_idata_buff_185__1_,
         oc8051_ram_top1_oc8051_idata_buff_185__2_,
         oc8051_ram_top1_oc8051_idata_buff_185__3_,
         oc8051_ram_top1_oc8051_idata_buff_185__4_,
         oc8051_ram_top1_oc8051_idata_buff_185__5_,
         oc8051_ram_top1_oc8051_idata_buff_185__6_,
         oc8051_ram_top1_oc8051_idata_buff_185__7_,
         oc8051_ram_top1_oc8051_idata_buff_184__0_,
         oc8051_ram_top1_oc8051_idata_buff_184__1_,
         oc8051_ram_top1_oc8051_idata_buff_184__2_,
         oc8051_ram_top1_oc8051_idata_buff_184__3_,
         oc8051_ram_top1_oc8051_idata_buff_184__4_,
         oc8051_ram_top1_oc8051_idata_buff_184__5_,
         oc8051_ram_top1_oc8051_idata_buff_184__6_,
         oc8051_ram_top1_oc8051_idata_buff_184__7_,
         oc8051_ram_top1_oc8051_idata_buff_181__0_,
         oc8051_ram_top1_oc8051_idata_buff_181__1_,
         oc8051_ram_top1_oc8051_idata_buff_181__2_,
         oc8051_ram_top1_oc8051_idata_buff_181__3_,
         oc8051_ram_top1_oc8051_idata_buff_181__4_,
         oc8051_ram_top1_oc8051_idata_buff_181__5_,
         oc8051_ram_top1_oc8051_idata_buff_181__6_,
         oc8051_ram_top1_oc8051_idata_buff_181__7_,
         oc8051_ram_top1_oc8051_idata_buff_180__0_,
         oc8051_ram_top1_oc8051_idata_buff_180__1_,
         oc8051_ram_top1_oc8051_idata_buff_180__2_,
         oc8051_ram_top1_oc8051_idata_buff_180__3_,
         oc8051_ram_top1_oc8051_idata_buff_180__4_,
         oc8051_ram_top1_oc8051_idata_buff_180__5_,
         oc8051_ram_top1_oc8051_idata_buff_180__6_,
         oc8051_ram_top1_oc8051_idata_buff_180__7_,
         oc8051_ram_top1_oc8051_idata_buff_177__0_,
         oc8051_ram_top1_oc8051_idata_buff_177__1_,
         oc8051_ram_top1_oc8051_idata_buff_177__2_,
         oc8051_ram_top1_oc8051_idata_buff_177__3_,
         oc8051_ram_top1_oc8051_idata_buff_177__4_,
         oc8051_ram_top1_oc8051_idata_buff_177__5_,
         oc8051_ram_top1_oc8051_idata_buff_177__6_,
         oc8051_ram_top1_oc8051_idata_buff_177__7_,
         oc8051_ram_top1_oc8051_idata_buff_176__0_,
         oc8051_ram_top1_oc8051_idata_buff_176__1_,
         oc8051_ram_top1_oc8051_idata_buff_176__2_,
         oc8051_ram_top1_oc8051_idata_buff_176__3_,
         oc8051_ram_top1_oc8051_idata_buff_176__4_,
         oc8051_ram_top1_oc8051_idata_buff_176__5_,
         oc8051_ram_top1_oc8051_idata_buff_176__6_,
         oc8051_ram_top1_oc8051_idata_buff_176__7_,
         oc8051_ram_top1_oc8051_idata_buff_175__0_,
         oc8051_ram_top1_oc8051_idata_buff_175__1_,
         oc8051_ram_top1_oc8051_idata_buff_175__2_,
         oc8051_ram_top1_oc8051_idata_buff_175__3_,
         oc8051_ram_top1_oc8051_idata_buff_175__4_,
         oc8051_ram_top1_oc8051_idata_buff_175__5_,
         oc8051_ram_top1_oc8051_idata_buff_175__6_,
         oc8051_ram_top1_oc8051_idata_buff_175__7_,
         oc8051_ram_top1_oc8051_idata_buff_174__0_,
         oc8051_ram_top1_oc8051_idata_buff_174__1_,
         oc8051_ram_top1_oc8051_idata_buff_174__2_,
         oc8051_ram_top1_oc8051_idata_buff_174__3_,
         oc8051_ram_top1_oc8051_idata_buff_174__4_,
         oc8051_ram_top1_oc8051_idata_buff_174__5_,
         oc8051_ram_top1_oc8051_idata_buff_174__6_,
         oc8051_ram_top1_oc8051_idata_buff_174__7_,
         oc8051_ram_top1_oc8051_idata_buff_173__0_,
         oc8051_ram_top1_oc8051_idata_buff_173__1_,
         oc8051_ram_top1_oc8051_idata_buff_173__2_,
         oc8051_ram_top1_oc8051_idata_buff_173__3_,
         oc8051_ram_top1_oc8051_idata_buff_173__4_,
         oc8051_ram_top1_oc8051_idata_buff_173__5_,
         oc8051_ram_top1_oc8051_idata_buff_173__6_,
         oc8051_ram_top1_oc8051_idata_buff_173__7_,
         oc8051_ram_top1_oc8051_idata_buff_172__0_,
         oc8051_ram_top1_oc8051_idata_buff_172__1_,
         oc8051_ram_top1_oc8051_idata_buff_172__2_,
         oc8051_ram_top1_oc8051_idata_buff_172__3_,
         oc8051_ram_top1_oc8051_idata_buff_172__4_,
         oc8051_ram_top1_oc8051_idata_buff_172__5_,
         oc8051_ram_top1_oc8051_idata_buff_172__6_,
         oc8051_ram_top1_oc8051_idata_buff_172__7_,
         oc8051_ram_top1_oc8051_idata_buff_171__0_,
         oc8051_ram_top1_oc8051_idata_buff_171__1_,
         oc8051_ram_top1_oc8051_idata_buff_171__2_,
         oc8051_ram_top1_oc8051_idata_buff_171__3_,
         oc8051_ram_top1_oc8051_idata_buff_171__4_,
         oc8051_ram_top1_oc8051_idata_buff_171__5_,
         oc8051_ram_top1_oc8051_idata_buff_171__6_,
         oc8051_ram_top1_oc8051_idata_buff_171__7_,
         oc8051_ram_top1_oc8051_idata_buff_170__0_,
         oc8051_ram_top1_oc8051_idata_buff_170__1_,
         oc8051_ram_top1_oc8051_idata_buff_170__2_,
         oc8051_ram_top1_oc8051_idata_buff_170__3_,
         oc8051_ram_top1_oc8051_idata_buff_170__4_,
         oc8051_ram_top1_oc8051_idata_buff_170__5_,
         oc8051_ram_top1_oc8051_idata_buff_170__6_,
         oc8051_ram_top1_oc8051_idata_buff_170__7_,
         oc8051_ram_top1_oc8051_idata_buff_169__0_,
         oc8051_ram_top1_oc8051_idata_buff_169__1_,
         oc8051_ram_top1_oc8051_idata_buff_169__2_,
         oc8051_ram_top1_oc8051_idata_buff_169__3_,
         oc8051_ram_top1_oc8051_idata_buff_169__4_,
         oc8051_ram_top1_oc8051_idata_buff_169__5_,
         oc8051_ram_top1_oc8051_idata_buff_169__6_,
         oc8051_ram_top1_oc8051_idata_buff_169__7_,
         oc8051_ram_top1_oc8051_idata_buff_168__0_,
         oc8051_ram_top1_oc8051_idata_buff_168__1_,
         oc8051_ram_top1_oc8051_idata_buff_168__2_,
         oc8051_ram_top1_oc8051_idata_buff_168__3_,
         oc8051_ram_top1_oc8051_idata_buff_168__4_,
         oc8051_ram_top1_oc8051_idata_buff_168__5_,
         oc8051_ram_top1_oc8051_idata_buff_168__6_,
         oc8051_ram_top1_oc8051_idata_buff_168__7_,
         oc8051_ram_top1_oc8051_idata_buff_167__0_,
         oc8051_ram_top1_oc8051_idata_buff_167__1_,
         oc8051_ram_top1_oc8051_idata_buff_167__2_,
         oc8051_ram_top1_oc8051_idata_buff_167__3_,
         oc8051_ram_top1_oc8051_idata_buff_167__4_,
         oc8051_ram_top1_oc8051_idata_buff_167__5_,
         oc8051_ram_top1_oc8051_idata_buff_167__6_,
         oc8051_ram_top1_oc8051_idata_buff_167__7_,
         oc8051_ram_top1_oc8051_idata_buff_166__0_,
         oc8051_ram_top1_oc8051_idata_buff_166__1_,
         oc8051_ram_top1_oc8051_idata_buff_166__2_,
         oc8051_ram_top1_oc8051_idata_buff_166__3_,
         oc8051_ram_top1_oc8051_idata_buff_166__4_,
         oc8051_ram_top1_oc8051_idata_buff_166__5_,
         oc8051_ram_top1_oc8051_idata_buff_166__6_,
         oc8051_ram_top1_oc8051_idata_buff_166__7_,
         oc8051_ram_top1_oc8051_idata_buff_163__0_,
         oc8051_ram_top1_oc8051_idata_buff_163__1_,
         oc8051_ram_top1_oc8051_idata_buff_163__2_,
         oc8051_ram_top1_oc8051_idata_buff_163__3_,
         oc8051_ram_top1_oc8051_idata_buff_163__4_,
         oc8051_ram_top1_oc8051_idata_buff_163__5_,
         oc8051_ram_top1_oc8051_idata_buff_163__6_,
         oc8051_ram_top1_oc8051_idata_buff_163__7_,
         oc8051_ram_top1_oc8051_idata_buff_162__0_,
         oc8051_ram_top1_oc8051_idata_buff_162__1_,
         oc8051_ram_top1_oc8051_idata_buff_162__2_,
         oc8051_ram_top1_oc8051_idata_buff_162__3_,
         oc8051_ram_top1_oc8051_idata_buff_162__4_,
         oc8051_ram_top1_oc8051_idata_buff_162__5_,
         oc8051_ram_top1_oc8051_idata_buff_162__6_,
         oc8051_ram_top1_oc8051_idata_buff_162__7_,
         oc8051_ram_top1_oc8051_idata_buff_159__0_,
         oc8051_ram_top1_oc8051_idata_buff_159__1_,
         oc8051_ram_top1_oc8051_idata_buff_159__2_,
         oc8051_ram_top1_oc8051_idata_buff_159__3_,
         oc8051_ram_top1_oc8051_idata_buff_159__4_,
         oc8051_ram_top1_oc8051_idata_buff_159__5_,
         oc8051_ram_top1_oc8051_idata_buff_159__6_,
         oc8051_ram_top1_oc8051_idata_buff_159__7_,
         oc8051_ram_top1_oc8051_idata_buff_158__0_,
         oc8051_ram_top1_oc8051_idata_buff_158__1_,
         oc8051_ram_top1_oc8051_idata_buff_158__2_,
         oc8051_ram_top1_oc8051_idata_buff_158__3_,
         oc8051_ram_top1_oc8051_idata_buff_158__4_,
         oc8051_ram_top1_oc8051_idata_buff_158__5_,
         oc8051_ram_top1_oc8051_idata_buff_158__6_,
         oc8051_ram_top1_oc8051_idata_buff_158__7_,
         oc8051_ram_top1_oc8051_idata_buff_157__0_,
         oc8051_ram_top1_oc8051_idata_buff_157__1_,
         oc8051_ram_top1_oc8051_idata_buff_157__2_,
         oc8051_ram_top1_oc8051_idata_buff_157__3_,
         oc8051_ram_top1_oc8051_idata_buff_157__4_,
         oc8051_ram_top1_oc8051_idata_buff_157__5_,
         oc8051_ram_top1_oc8051_idata_buff_157__6_,
         oc8051_ram_top1_oc8051_idata_buff_157__7_,
         oc8051_ram_top1_oc8051_idata_buff_156__0_,
         oc8051_ram_top1_oc8051_idata_buff_156__1_,
         oc8051_ram_top1_oc8051_idata_buff_156__2_,
         oc8051_ram_top1_oc8051_idata_buff_156__3_,
         oc8051_ram_top1_oc8051_idata_buff_156__4_,
         oc8051_ram_top1_oc8051_idata_buff_156__5_,
         oc8051_ram_top1_oc8051_idata_buff_156__6_,
         oc8051_ram_top1_oc8051_idata_buff_156__7_,
         oc8051_ram_top1_oc8051_idata_buff_155__0_,
         oc8051_ram_top1_oc8051_idata_buff_155__1_,
         oc8051_ram_top1_oc8051_idata_buff_155__2_,
         oc8051_ram_top1_oc8051_idata_buff_155__3_,
         oc8051_ram_top1_oc8051_idata_buff_155__4_,
         oc8051_ram_top1_oc8051_idata_buff_155__5_,
         oc8051_ram_top1_oc8051_idata_buff_155__6_,
         oc8051_ram_top1_oc8051_idata_buff_155__7_,
         oc8051_ram_top1_oc8051_idata_buff_154__0_,
         oc8051_ram_top1_oc8051_idata_buff_154__1_,
         oc8051_ram_top1_oc8051_idata_buff_154__2_,
         oc8051_ram_top1_oc8051_idata_buff_154__3_,
         oc8051_ram_top1_oc8051_idata_buff_154__4_,
         oc8051_ram_top1_oc8051_idata_buff_154__5_,
         oc8051_ram_top1_oc8051_idata_buff_154__6_,
         oc8051_ram_top1_oc8051_idata_buff_154__7_,
         oc8051_ram_top1_oc8051_idata_buff_153__0_,
         oc8051_ram_top1_oc8051_idata_buff_153__1_,
         oc8051_ram_top1_oc8051_idata_buff_153__2_,
         oc8051_ram_top1_oc8051_idata_buff_153__3_,
         oc8051_ram_top1_oc8051_idata_buff_153__4_,
         oc8051_ram_top1_oc8051_idata_buff_153__5_,
         oc8051_ram_top1_oc8051_idata_buff_153__6_,
         oc8051_ram_top1_oc8051_idata_buff_153__7_,
         oc8051_ram_top1_oc8051_idata_buff_152__0_,
         oc8051_ram_top1_oc8051_idata_buff_152__1_,
         oc8051_ram_top1_oc8051_idata_buff_152__2_,
         oc8051_ram_top1_oc8051_idata_buff_152__3_,
         oc8051_ram_top1_oc8051_idata_buff_152__4_,
         oc8051_ram_top1_oc8051_idata_buff_152__5_,
         oc8051_ram_top1_oc8051_idata_buff_152__6_,
         oc8051_ram_top1_oc8051_idata_buff_152__7_,
         oc8051_ram_top1_oc8051_idata_buff_151__0_,
         oc8051_ram_top1_oc8051_idata_buff_151__1_,
         oc8051_ram_top1_oc8051_idata_buff_151__2_,
         oc8051_ram_top1_oc8051_idata_buff_151__3_,
         oc8051_ram_top1_oc8051_idata_buff_151__4_,
         oc8051_ram_top1_oc8051_idata_buff_151__5_,
         oc8051_ram_top1_oc8051_idata_buff_151__6_,
         oc8051_ram_top1_oc8051_idata_buff_151__7_,
         oc8051_ram_top1_oc8051_idata_buff_150__0_,
         oc8051_ram_top1_oc8051_idata_buff_150__1_,
         oc8051_ram_top1_oc8051_idata_buff_150__2_,
         oc8051_ram_top1_oc8051_idata_buff_150__3_,
         oc8051_ram_top1_oc8051_idata_buff_150__4_,
         oc8051_ram_top1_oc8051_idata_buff_150__5_,
         oc8051_ram_top1_oc8051_idata_buff_150__6_,
         oc8051_ram_top1_oc8051_idata_buff_150__7_,
         oc8051_ram_top1_oc8051_idata_buff_149__0_,
         oc8051_ram_top1_oc8051_idata_buff_149__1_,
         oc8051_ram_top1_oc8051_idata_buff_149__2_,
         oc8051_ram_top1_oc8051_idata_buff_149__3_,
         oc8051_ram_top1_oc8051_idata_buff_149__4_,
         oc8051_ram_top1_oc8051_idata_buff_149__5_,
         oc8051_ram_top1_oc8051_idata_buff_149__6_,
         oc8051_ram_top1_oc8051_idata_buff_149__7_,
         oc8051_ram_top1_oc8051_idata_buff_148__0_,
         oc8051_ram_top1_oc8051_idata_buff_148__1_,
         oc8051_ram_top1_oc8051_idata_buff_148__2_,
         oc8051_ram_top1_oc8051_idata_buff_148__3_,
         oc8051_ram_top1_oc8051_idata_buff_148__4_,
         oc8051_ram_top1_oc8051_idata_buff_148__5_,
         oc8051_ram_top1_oc8051_idata_buff_148__6_,
         oc8051_ram_top1_oc8051_idata_buff_148__7_,
         oc8051_ram_top1_oc8051_idata_buff_147__0_,
         oc8051_ram_top1_oc8051_idata_buff_147__1_,
         oc8051_ram_top1_oc8051_idata_buff_147__2_,
         oc8051_ram_top1_oc8051_idata_buff_147__3_,
         oc8051_ram_top1_oc8051_idata_buff_147__4_,
         oc8051_ram_top1_oc8051_idata_buff_147__5_,
         oc8051_ram_top1_oc8051_idata_buff_147__6_,
         oc8051_ram_top1_oc8051_idata_buff_147__7_,
         oc8051_ram_top1_oc8051_idata_buff_146__0_,
         oc8051_ram_top1_oc8051_idata_buff_146__1_,
         oc8051_ram_top1_oc8051_idata_buff_146__2_,
         oc8051_ram_top1_oc8051_idata_buff_146__3_,
         oc8051_ram_top1_oc8051_idata_buff_146__4_,
         oc8051_ram_top1_oc8051_idata_buff_146__5_,
         oc8051_ram_top1_oc8051_idata_buff_146__6_,
         oc8051_ram_top1_oc8051_idata_buff_146__7_,
         oc8051_ram_top1_oc8051_idata_buff_145__0_,
         oc8051_ram_top1_oc8051_idata_buff_145__1_,
         oc8051_ram_top1_oc8051_idata_buff_145__2_,
         oc8051_ram_top1_oc8051_idata_buff_145__3_,
         oc8051_ram_top1_oc8051_idata_buff_145__4_,
         oc8051_ram_top1_oc8051_idata_buff_145__5_,
         oc8051_ram_top1_oc8051_idata_buff_145__6_,
         oc8051_ram_top1_oc8051_idata_buff_145__7_,
         oc8051_ram_top1_oc8051_idata_buff_144__0_,
         oc8051_ram_top1_oc8051_idata_buff_144__1_,
         oc8051_ram_top1_oc8051_idata_buff_144__2_,
         oc8051_ram_top1_oc8051_idata_buff_144__3_,
         oc8051_ram_top1_oc8051_idata_buff_144__4_,
         oc8051_ram_top1_oc8051_idata_buff_144__5_,
         oc8051_ram_top1_oc8051_idata_buff_144__6_,
         oc8051_ram_top1_oc8051_idata_buff_144__7_,
         oc8051_ram_top1_oc8051_idata_buff_141__0_,
         oc8051_ram_top1_oc8051_idata_buff_141__1_,
         oc8051_ram_top1_oc8051_idata_buff_141__2_,
         oc8051_ram_top1_oc8051_idata_buff_141__3_,
         oc8051_ram_top1_oc8051_idata_buff_141__4_,
         oc8051_ram_top1_oc8051_idata_buff_141__5_,
         oc8051_ram_top1_oc8051_idata_buff_141__6_,
         oc8051_ram_top1_oc8051_idata_buff_141__7_,
         oc8051_ram_top1_oc8051_idata_buff_140__0_,
         oc8051_ram_top1_oc8051_idata_buff_140__1_,
         oc8051_ram_top1_oc8051_idata_buff_140__2_,
         oc8051_ram_top1_oc8051_idata_buff_140__3_,
         oc8051_ram_top1_oc8051_idata_buff_140__4_,
         oc8051_ram_top1_oc8051_idata_buff_140__5_,
         oc8051_ram_top1_oc8051_idata_buff_140__6_,
         oc8051_ram_top1_oc8051_idata_buff_140__7_,
         oc8051_ram_top1_oc8051_idata_buff_139__0_,
         oc8051_ram_top1_oc8051_idata_buff_139__1_,
         oc8051_ram_top1_oc8051_idata_buff_139__2_,
         oc8051_ram_top1_oc8051_idata_buff_139__3_,
         oc8051_ram_top1_oc8051_idata_buff_139__4_,
         oc8051_ram_top1_oc8051_idata_buff_139__5_,
         oc8051_ram_top1_oc8051_idata_buff_139__6_,
         oc8051_ram_top1_oc8051_idata_buff_139__7_,
         oc8051_ram_top1_oc8051_idata_buff_138__0_,
         oc8051_ram_top1_oc8051_idata_buff_138__1_,
         oc8051_ram_top1_oc8051_idata_buff_138__2_,
         oc8051_ram_top1_oc8051_idata_buff_138__3_,
         oc8051_ram_top1_oc8051_idata_buff_138__4_,
         oc8051_ram_top1_oc8051_idata_buff_138__5_,
         oc8051_ram_top1_oc8051_idata_buff_138__6_,
         oc8051_ram_top1_oc8051_idata_buff_138__7_,
         oc8051_ram_top1_oc8051_idata_buff_135__0_,
         oc8051_ram_top1_oc8051_idata_buff_135__1_,
         oc8051_ram_top1_oc8051_idata_buff_135__2_,
         oc8051_ram_top1_oc8051_idata_buff_135__3_,
         oc8051_ram_top1_oc8051_idata_buff_135__4_,
         oc8051_ram_top1_oc8051_idata_buff_135__5_,
         oc8051_ram_top1_oc8051_idata_buff_135__6_,
         oc8051_ram_top1_oc8051_idata_buff_135__7_,
         oc8051_ram_top1_oc8051_idata_buff_134__0_,
         oc8051_ram_top1_oc8051_idata_buff_134__1_,
         oc8051_ram_top1_oc8051_idata_buff_134__2_,
         oc8051_ram_top1_oc8051_idata_buff_134__3_,
         oc8051_ram_top1_oc8051_idata_buff_134__4_,
         oc8051_ram_top1_oc8051_idata_buff_134__5_,
         oc8051_ram_top1_oc8051_idata_buff_134__6_,
         oc8051_ram_top1_oc8051_idata_buff_134__7_,
         oc8051_ram_top1_oc8051_idata_buff_131__0_,
         oc8051_ram_top1_oc8051_idata_buff_131__1_,
         oc8051_ram_top1_oc8051_idata_buff_131__2_,
         oc8051_ram_top1_oc8051_idata_buff_131__3_,
         oc8051_ram_top1_oc8051_idata_buff_131__4_,
         oc8051_ram_top1_oc8051_idata_buff_131__5_,
         oc8051_ram_top1_oc8051_idata_buff_131__6_,
         oc8051_ram_top1_oc8051_idata_buff_131__7_,
         oc8051_ram_top1_oc8051_idata_buff_130__0_,
         oc8051_ram_top1_oc8051_idata_buff_130__1_,
         oc8051_ram_top1_oc8051_idata_buff_130__2_,
         oc8051_ram_top1_oc8051_idata_buff_130__3_,
         oc8051_ram_top1_oc8051_idata_buff_130__4_,
         oc8051_ram_top1_oc8051_idata_buff_130__5_,
         oc8051_ram_top1_oc8051_idata_buff_130__6_,
         oc8051_ram_top1_oc8051_idata_buff_130__7_,
         oc8051_ram_top1_oc8051_idata_buff_255__0_,
         oc8051_ram_top1_oc8051_idata_buff_255__1_,
         oc8051_ram_top1_oc8051_idata_buff_255__2_,
         oc8051_ram_top1_oc8051_idata_buff_255__3_,
         oc8051_ram_top1_oc8051_idata_buff_255__4_,
         oc8051_ram_top1_oc8051_idata_buff_255__5_,
         oc8051_ram_top1_oc8051_idata_buff_255__6_,
         oc8051_ram_top1_oc8051_idata_buff_255__7_,
         oc8051_ram_top1_oc8051_idata_buff_254__0_,
         oc8051_ram_top1_oc8051_idata_buff_254__1_,
         oc8051_ram_top1_oc8051_idata_buff_254__2_,
         oc8051_ram_top1_oc8051_idata_buff_254__3_,
         oc8051_ram_top1_oc8051_idata_buff_254__4_,
         oc8051_ram_top1_oc8051_idata_buff_254__5_,
         oc8051_ram_top1_oc8051_idata_buff_254__6_,
         oc8051_ram_top1_oc8051_idata_buff_254__7_,
         oc8051_ram_top1_oc8051_idata_buff_253__0_,
         oc8051_ram_top1_oc8051_idata_buff_253__1_,
         oc8051_ram_top1_oc8051_idata_buff_253__2_,
         oc8051_ram_top1_oc8051_idata_buff_253__3_,
         oc8051_ram_top1_oc8051_idata_buff_253__4_,
         oc8051_ram_top1_oc8051_idata_buff_253__5_,
         oc8051_ram_top1_oc8051_idata_buff_253__6_,
         oc8051_ram_top1_oc8051_idata_buff_253__7_,
         oc8051_ram_top1_oc8051_idata_buff_252__0_,
         oc8051_ram_top1_oc8051_idata_buff_252__1_,
         oc8051_ram_top1_oc8051_idata_buff_252__2_,
         oc8051_ram_top1_oc8051_idata_buff_252__3_,
         oc8051_ram_top1_oc8051_idata_buff_252__4_,
         oc8051_ram_top1_oc8051_idata_buff_252__5_,
         oc8051_ram_top1_oc8051_idata_buff_252__6_,
         oc8051_ram_top1_oc8051_idata_buff_252__7_,
         oc8051_ram_top1_oc8051_idata_buff_251__0_,
         oc8051_ram_top1_oc8051_idata_buff_251__1_,
         oc8051_ram_top1_oc8051_idata_buff_251__2_,
         oc8051_ram_top1_oc8051_idata_buff_251__3_,
         oc8051_ram_top1_oc8051_idata_buff_251__4_,
         oc8051_ram_top1_oc8051_idata_buff_251__5_,
         oc8051_ram_top1_oc8051_idata_buff_251__6_,
         oc8051_ram_top1_oc8051_idata_buff_251__7_,
         oc8051_ram_top1_oc8051_idata_buff_250__0_,
         oc8051_ram_top1_oc8051_idata_buff_250__1_,
         oc8051_ram_top1_oc8051_idata_buff_250__2_,
         oc8051_ram_top1_oc8051_idata_buff_250__3_,
         oc8051_ram_top1_oc8051_idata_buff_250__4_,
         oc8051_ram_top1_oc8051_idata_buff_250__5_,
         oc8051_ram_top1_oc8051_idata_buff_250__6_,
         oc8051_ram_top1_oc8051_idata_buff_250__7_,
         oc8051_ram_top1_oc8051_idata_buff_249__0_,
         oc8051_ram_top1_oc8051_idata_buff_249__1_,
         oc8051_ram_top1_oc8051_idata_buff_249__2_,
         oc8051_ram_top1_oc8051_idata_buff_249__3_,
         oc8051_ram_top1_oc8051_idata_buff_249__4_,
         oc8051_ram_top1_oc8051_idata_buff_249__5_,
         oc8051_ram_top1_oc8051_idata_buff_249__6_,
         oc8051_ram_top1_oc8051_idata_buff_249__7_,
         oc8051_ram_top1_oc8051_idata_buff_248__0_,
         oc8051_ram_top1_oc8051_idata_buff_248__1_,
         oc8051_ram_top1_oc8051_idata_buff_248__2_,
         oc8051_ram_top1_oc8051_idata_buff_248__3_,
         oc8051_ram_top1_oc8051_idata_buff_248__4_,
         oc8051_ram_top1_oc8051_idata_buff_248__5_,
         oc8051_ram_top1_oc8051_idata_buff_248__6_,
         oc8051_ram_top1_oc8051_idata_buff_248__7_,
         oc8051_ram_top1_oc8051_idata_buff_245__0_,
         oc8051_ram_top1_oc8051_idata_buff_245__1_,
         oc8051_ram_top1_oc8051_idata_buff_245__2_,
         oc8051_ram_top1_oc8051_idata_buff_245__3_,
         oc8051_ram_top1_oc8051_idata_buff_245__4_,
         oc8051_ram_top1_oc8051_idata_buff_245__5_,
         oc8051_ram_top1_oc8051_idata_buff_245__6_,
         oc8051_ram_top1_oc8051_idata_buff_245__7_,
         oc8051_ram_top1_oc8051_idata_buff_244__0_,
         oc8051_ram_top1_oc8051_idata_buff_244__1_,
         oc8051_ram_top1_oc8051_idata_buff_244__2_,
         oc8051_ram_top1_oc8051_idata_buff_244__3_,
         oc8051_ram_top1_oc8051_idata_buff_244__4_,
         oc8051_ram_top1_oc8051_idata_buff_244__5_,
         oc8051_ram_top1_oc8051_idata_buff_244__6_,
         oc8051_ram_top1_oc8051_idata_buff_244__7_,
         oc8051_ram_top1_oc8051_idata_buff_241__0_,
         oc8051_ram_top1_oc8051_idata_buff_241__1_,
         oc8051_ram_top1_oc8051_idata_buff_241__2_,
         oc8051_ram_top1_oc8051_idata_buff_241__3_,
         oc8051_ram_top1_oc8051_idata_buff_241__4_,
         oc8051_ram_top1_oc8051_idata_buff_241__5_,
         oc8051_ram_top1_oc8051_idata_buff_241__6_,
         oc8051_ram_top1_oc8051_idata_buff_241__7_,
         oc8051_ram_top1_oc8051_idata_buff_240__0_,
         oc8051_ram_top1_oc8051_idata_buff_240__1_,
         oc8051_ram_top1_oc8051_idata_buff_240__2_,
         oc8051_ram_top1_oc8051_idata_buff_240__3_,
         oc8051_ram_top1_oc8051_idata_buff_240__4_,
         oc8051_ram_top1_oc8051_idata_buff_240__5_,
         oc8051_ram_top1_oc8051_idata_buff_240__6_,
         oc8051_ram_top1_oc8051_idata_buff_240__7_,
         oc8051_ram_top1_oc8051_idata_buff_239__0_,
         oc8051_ram_top1_oc8051_idata_buff_239__1_,
         oc8051_ram_top1_oc8051_idata_buff_239__2_,
         oc8051_ram_top1_oc8051_idata_buff_239__3_,
         oc8051_ram_top1_oc8051_idata_buff_239__4_,
         oc8051_ram_top1_oc8051_idata_buff_239__5_,
         oc8051_ram_top1_oc8051_idata_buff_239__6_,
         oc8051_ram_top1_oc8051_idata_buff_239__7_,
         oc8051_ram_top1_oc8051_idata_buff_238__0_,
         oc8051_ram_top1_oc8051_idata_buff_238__1_,
         oc8051_ram_top1_oc8051_idata_buff_238__2_,
         oc8051_ram_top1_oc8051_idata_buff_238__3_,
         oc8051_ram_top1_oc8051_idata_buff_238__4_,
         oc8051_ram_top1_oc8051_idata_buff_238__5_,
         oc8051_ram_top1_oc8051_idata_buff_238__6_,
         oc8051_ram_top1_oc8051_idata_buff_238__7_,
         oc8051_ram_top1_oc8051_idata_buff_237__0_,
         oc8051_ram_top1_oc8051_idata_buff_237__1_,
         oc8051_ram_top1_oc8051_idata_buff_237__2_,
         oc8051_ram_top1_oc8051_idata_buff_237__3_,
         oc8051_ram_top1_oc8051_idata_buff_237__4_,
         oc8051_ram_top1_oc8051_idata_buff_237__5_,
         oc8051_ram_top1_oc8051_idata_buff_237__6_,
         oc8051_ram_top1_oc8051_idata_buff_237__7_,
         oc8051_ram_top1_oc8051_idata_buff_236__0_,
         oc8051_ram_top1_oc8051_idata_buff_236__1_,
         oc8051_ram_top1_oc8051_idata_buff_236__2_,
         oc8051_ram_top1_oc8051_idata_buff_236__3_,
         oc8051_ram_top1_oc8051_idata_buff_236__4_,
         oc8051_ram_top1_oc8051_idata_buff_236__5_,
         oc8051_ram_top1_oc8051_idata_buff_236__6_,
         oc8051_ram_top1_oc8051_idata_buff_236__7_,
         oc8051_ram_top1_oc8051_idata_buff_235__0_,
         oc8051_ram_top1_oc8051_idata_buff_235__1_,
         oc8051_ram_top1_oc8051_idata_buff_235__2_,
         oc8051_ram_top1_oc8051_idata_buff_235__3_,
         oc8051_ram_top1_oc8051_idata_buff_235__4_,
         oc8051_ram_top1_oc8051_idata_buff_235__5_,
         oc8051_ram_top1_oc8051_idata_buff_235__6_,
         oc8051_ram_top1_oc8051_idata_buff_235__7_,
         oc8051_ram_top1_oc8051_idata_buff_234__0_,
         oc8051_ram_top1_oc8051_idata_buff_234__1_,
         oc8051_ram_top1_oc8051_idata_buff_234__2_,
         oc8051_ram_top1_oc8051_idata_buff_234__3_,
         oc8051_ram_top1_oc8051_idata_buff_234__4_,
         oc8051_ram_top1_oc8051_idata_buff_234__5_,
         oc8051_ram_top1_oc8051_idata_buff_234__6_,
         oc8051_ram_top1_oc8051_idata_buff_234__7_,
         oc8051_ram_top1_oc8051_idata_buff_233__0_,
         oc8051_ram_top1_oc8051_idata_buff_233__1_,
         oc8051_ram_top1_oc8051_idata_buff_233__2_,
         oc8051_ram_top1_oc8051_idata_buff_233__3_,
         oc8051_ram_top1_oc8051_idata_buff_233__4_,
         oc8051_ram_top1_oc8051_idata_buff_233__5_,
         oc8051_ram_top1_oc8051_idata_buff_233__6_,
         oc8051_ram_top1_oc8051_idata_buff_233__7_,
         oc8051_ram_top1_oc8051_idata_buff_232__0_,
         oc8051_ram_top1_oc8051_idata_buff_232__1_,
         oc8051_ram_top1_oc8051_idata_buff_232__2_,
         oc8051_ram_top1_oc8051_idata_buff_232__3_,
         oc8051_ram_top1_oc8051_idata_buff_232__4_,
         oc8051_ram_top1_oc8051_idata_buff_232__5_,
         oc8051_ram_top1_oc8051_idata_buff_232__6_,
         oc8051_ram_top1_oc8051_idata_buff_232__7_,
         oc8051_ram_top1_oc8051_idata_buff_231__0_,
         oc8051_ram_top1_oc8051_idata_buff_231__1_,
         oc8051_ram_top1_oc8051_idata_buff_231__2_,
         oc8051_ram_top1_oc8051_idata_buff_231__3_,
         oc8051_ram_top1_oc8051_idata_buff_231__4_,
         oc8051_ram_top1_oc8051_idata_buff_231__5_,
         oc8051_ram_top1_oc8051_idata_buff_231__6_,
         oc8051_ram_top1_oc8051_idata_buff_231__7_,
         oc8051_ram_top1_oc8051_idata_buff_230__0_,
         oc8051_ram_top1_oc8051_idata_buff_230__1_,
         oc8051_ram_top1_oc8051_idata_buff_230__2_,
         oc8051_ram_top1_oc8051_idata_buff_230__3_,
         oc8051_ram_top1_oc8051_idata_buff_230__4_,
         oc8051_ram_top1_oc8051_idata_buff_230__5_,
         oc8051_ram_top1_oc8051_idata_buff_230__6_,
         oc8051_ram_top1_oc8051_idata_buff_230__7_,
         oc8051_ram_top1_oc8051_idata_buff_227__0_,
         oc8051_ram_top1_oc8051_idata_buff_227__1_,
         oc8051_ram_top1_oc8051_idata_buff_227__2_,
         oc8051_ram_top1_oc8051_idata_buff_227__3_,
         oc8051_ram_top1_oc8051_idata_buff_227__4_,
         oc8051_ram_top1_oc8051_idata_buff_227__5_,
         oc8051_ram_top1_oc8051_idata_buff_227__6_,
         oc8051_ram_top1_oc8051_idata_buff_227__7_,
         oc8051_ram_top1_oc8051_idata_buff_226__0_,
         oc8051_ram_top1_oc8051_idata_buff_226__1_,
         oc8051_ram_top1_oc8051_idata_buff_226__2_,
         oc8051_ram_top1_oc8051_idata_buff_226__3_,
         oc8051_ram_top1_oc8051_idata_buff_226__4_,
         oc8051_ram_top1_oc8051_idata_buff_226__5_,
         oc8051_ram_top1_oc8051_idata_buff_226__6_,
         oc8051_ram_top1_oc8051_idata_buff_226__7_,
         oc8051_ram_top1_oc8051_idata_buff_223__0_,
         oc8051_ram_top1_oc8051_idata_buff_223__1_,
         oc8051_ram_top1_oc8051_idata_buff_223__2_,
         oc8051_ram_top1_oc8051_idata_buff_223__3_,
         oc8051_ram_top1_oc8051_idata_buff_223__4_,
         oc8051_ram_top1_oc8051_idata_buff_223__5_,
         oc8051_ram_top1_oc8051_idata_buff_223__6_,
         oc8051_ram_top1_oc8051_idata_buff_223__7_,
         oc8051_ram_top1_oc8051_idata_buff_222__0_,
         oc8051_ram_top1_oc8051_idata_buff_222__1_,
         oc8051_ram_top1_oc8051_idata_buff_222__2_,
         oc8051_ram_top1_oc8051_idata_buff_222__3_,
         oc8051_ram_top1_oc8051_idata_buff_222__4_,
         oc8051_ram_top1_oc8051_idata_buff_222__5_,
         oc8051_ram_top1_oc8051_idata_buff_222__6_,
         oc8051_ram_top1_oc8051_idata_buff_222__7_,
         oc8051_ram_top1_oc8051_idata_buff_221__0_,
         oc8051_ram_top1_oc8051_idata_buff_221__1_,
         oc8051_ram_top1_oc8051_idata_buff_221__2_,
         oc8051_ram_top1_oc8051_idata_buff_221__3_,
         oc8051_ram_top1_oc8051_idata_buff_221__4_,
         oc8051_ram_top1_oc8051_idata_buff_221__5_,
         oc8051_ram_top1_oc8051_idata_buff_221__6_,
         oc8051_ram_top1_oc8051_idata_buff_221__7_,
         oc8051_ram_top1_oc8051_idata_buff_220__0_,
         oc8051_ram_top1_oc8051_idata_buff_220__1_,
         oc8051_ram_top1_oc8051_idata_buff_220__2_,
         oc8051_ram_top1_oc8051_idata_buff_220__3_,
         oc8051_ram_top1_oc8051_idata_buff_220__4_,
         oc8051_ram_top1_oc8051_idata_buff_220__5_,
         oc8051_ram_top1_oc8051_idata_buff_220__6_,
         oc8051_ram_top1_oc8051_idata_buff_220__7_,
         oc8051_ram_top1_oc8051_idata_buff_219__0_,
         oc8051_ram_top1_oc8051_idata_buff_219__1_,
         oc8051_ram_top1_oc8051_idata_buff_219__2_,
         oc8051_ram_top1_oc8051_idata_buff_219__3_,
         oc8051_ram_top1_oc8051_idata_buff_219__4_,
         oc8051_ram_top1_oc8051_idata_buff_219__5_,
         oc8051_ram_top1_oc8051_idata_buff_219__6_,
         oc8051_ram_top1_oc8051_idata_buff_219__7_,
         oc8051_ram_top1_oc8051_idata_buff_218__0_,
         oc8051_ram_top1_oc8051_idata_buff_218__1_,
         oc8051_ram_top1_oc8051_idata_buff_218__2_,
         oc8051_ram_top1_oc8051_idata_buff_218__3_,
         oc8051_ram_top1_oc8051_idata_buff_218__4_,
         oc8051_ram_top1_oc8051_idata_buff_218__5_,
         oc8051_ram_top1_oc8051_idata_buff_218__6_,
         oc8051_ram_top1_oc8051_idata_buff_218__7_,
         oc8051_ram_top1_oc8051_idata_buff_217__0_,
         oc8051_ram_top1_oc8051_idata_buff_217__1_,
         oc8051_ram_top1_oc8051_idata_buff_217__2_,
         oc8051_ram_top1_oc8051_idata_buff_217__3_,
         oc8051_ram_top1_oc8051_idata_buff_217__4_,
         oc8051_ram_top1_oc8051_idata_buff_217__5_,
         oc8051_ram_top1_oc8051_idata_buff_217__6_,
         oc8051_ram_top1_oc8051_idata_buff_217__7_,
         oc8051_ram_top1_oc8051_idata_buff_216__0_,
         oc8051_ram_top1_oc8051_idata_buff_216__1_,
         oc8051_ram_top1_oc8051_idata_buff_216__2_,
         oc8051_ram_top1_oc8051_idata_buff_216__3_,
         oc8051_ram_top1_oc8051_idata_buff_216__4_,
         oc8051_ram_top1_oc8051_idata_buff_216__5_,
         oc8051_ram_top1_oc8051_idata_buff_216__6_,
         oc8051_ram_top1_oc8051_idata_buff_216__7_,
         oc8051_ram_top1_oc8051_idata_buff_215__0_,
         oc8051_ram_top1_oc8051_idata_buff_215__1_,
         oc8051_ram_top1_oc8051_idata_buff_215__2_,
         oc8051_ram_top1_oc8051_idata_buff_215__3_,
         oc8051_ram_top1_oc8051_idata_buff_215__4_,
         oc8051_ram_top1_oc8051_idata_buff_215__5_,
         oc8051_ram_top1_oc8051_idata_buff_215__6_,
         oc8051_ram_top1_oc8051_idata_buff_215__7_,
         oc8051_ram_top1_oc8051_idata_buff_214__0_,
         oc8051_ram_top1_oc8051_idata_buff_214__1_,
         oc8051_ram_top1_oc8051_idata_buff_214__2_,
         oc8051_ram_top1_oc8051_idata_buff_214__3_,
         oc8051_ram_top1_oc8051_idata_buff_214__4_,
         oc8051_ram_top1_oc8051_idata_buff_214__5_,
         oc8051_ram_top1_oc8051_idata_buff_214__6_,
         oc8051_ram_top1_oc8051_idata_buff_214__7_,
         oc8051_ram_top1_oc8051_idata_buff_213__0_,
         oc8051_ram_top1_oc8051_idata_buff_213__1_,
         oc8051_ram_top1_oc8051_idata_buff_213__2_,
         oc8051_ram_top1_oc8051_idata_buff_213__3_,
         oc8051_ram_top1_oc8051_idata_buff_213__4_,
         oc8051_ram_top1_oc8051_idata_buff_213__5_,
         oc8051_ram_top1_oc8051_idata_buff_213__6_,
         oc8051_ram_top1_oc8051_idata_buff_213__7_,
         oc8051_ram_top1_oc8051_idata_buff_212__0_,
         oc8051_ram_top1_oc8051_idata_buff_212__1_,
         oc8051_ram_top1_oc8051_idata_buff_212__2_,
         oc8051_ram_top1_oc8051_idata_buff_212__3_,
         oc8051_ram_top1_oc8051_idata_buff_212__4_,
         oc8051_ram_top1_oc8051_idata_buff_212__5_,
         oc8051_ram_top1_oc8051_idata_buff_212__6_,
         oc8051_ram_top1_oc8051_idata_buff_212__7_,
         oc8051_ram_top1_oc8051_idata_buff_211__0_,
         oc8051_ram_top1_oc8051_idata_buff_211__1_,
         oc8051_ram_top1_oc8051_idata_buff_211__2_,
         oc8051_ram_top1_oc8051_idata_buff_211__3_,
         oc8051_ram_top1_oc8051_idata_buff_211__4_,
         oc8051_ram_top1_oc8051_idata_buff_211__5_,
         oc8051_ram_top1_oc8051_idata_buff_211__6_,
         oc8051_ram_top1_oc8051_idata_buff_211__7_,
         oc8051_ram_top1_oc8051_idata_buff_210__0_,
         oc8051_ram_top1_oc8051_idata_buff_210__1_,
         oc8051_ram_top1_oc8051_idata_buff_210__2_,
         oc8051_ram_top1_oc8051_idata_buff_210__3_,
         oc8051_ram_top1_oc8051_idata_buff_210__4_,
         oc8051_ram_top1_oc8051_idata_buff_210__5_,
         oc8051_ram_top1_oc8051_idata_buff_210__6_,
         oc8051_ram_top1_oc8051_idata_buff_210__7_,
         oc8051_ram_top1_oc8051_idata_buff_209__0_,
         oc8051_ram_top1_oc8051_idata_buff_209__1_,
         oc8051_ram_top1_oc8051_idata_buff_209__2_,
         oc8051_ram_top1_oc8051_idata_buff_209__3_,
         oc8051_ram_top1_oc8051_idata_buff_209__4_,
         oc8051_ram_top1_oc8051_idata_buff_209__5_,
         oc8051_ram_top1_oc8051_idata_buff_209__6_,
         oc8051_ram_top1_oc8051_idata_buff_209__7_,
         oc8051_ram_top1_oc8051_idata_buff_208__0_,
         oc8051_ram_top1_oc8051_idata_buff_208__1_,
         oc8051_ram_top1_oc8051_idata_buff_208__2_,
         oc8051_ram_top1_oc8051_idata_buff_208__3_,
         oc8051_ram_top1_oc8051_idata_buff_208__4_,
         oc8051_ram_top1_oc8051_idata_buff_208__5_,
         oc8051_ram_top1_oc8051_idata_buff_208__6_,
         oc8051_ram_top1_oc8051_idata_buff_208__7_,
         oc8051_ram_top1_oc8051_idata_buff_205__0_,
         oc8051_ram_top1_oc8051_idata_buff_205__1_,
         oc8051_ram_top1_oc8051_idata_buff_205__2_,
         oc8051_ram_top1_oc8051_idata_buff_205__3_,
         oc8051_ram_top1_oc8051_idata_buff_205__4_,
         oc8051_ram_top1_oc8051_idata_buff_205__5_,
         oc8051_ram_top1_oc8051_idata_buff_205__6_,
         oc8051_ram_top1_oc8051_idata_buff_205__7_,
         oc8051_ram_top1_oc8051_idata_buff_204__0_,
         oc8051_ram_top1_oc8051_idata_buff_204__1_,
         oc8051_ram_top1_oc8051_idata_buff_204__2_,
         oc8051_ram_top1_oc8051_idata_buff_204__3_,
         oc8051_ram_top1_oc8051_idata_buff_204__4_,
         oc8051_ram_top1_oc8051_idata_buff_204__5_,
         oc8051_ram_top1_oc8051_idata_buff_204__6_,
         oc8051_ram_top1_oc8051_idata_buff_204__7_,
         oc8051_ram_top1_oc8051_idata_buff_203__0_,
         oc8051_ram_top1_oc8051_idata_buff_203__1_,
         oc8051_ram_top1_oc8051_idata_buff_203__2_,
         oc8051_ram_top1_oc8051_idata_buff_203__3_,
         oc8051_ram_top1_oc8051_idata_buff_203__4_,
         oc8051_ram_top1_oc8051_idata_buff_203__5_,
         oc8051_ram_top1_oc8051_idata_buff_203__6_,
         oc8051_ram_top1_oc8051_idata_buff_203__7_,
         oc8051_ram_top1_oc8051_idata_buff_202__0_,
         oc8051_ram_top1_oc8051_idata_buff_202__1_,
         oc8051_ram_top1_oc8051_idata_buff_202__2_,
         oc8051_ram_top1_oc8051_idata_buff_202__3_,
         oc8051_ram_top1_oc8051_idata_buff_202__4_,
         oc8051_ram_top1_oc8051_idata_buff_202__5_,
         oc8051_ram_top1_oc8051_idata_buff_202__6_,
         oc8051_ram_top1_oc8051_idata_buff_202__7_,
         oc8051_ram_top1_oc8051_idata_buff_199__0_,
         oc8051_ram_top1_oc8051_idata_buff_199__1_,
         oc8051_ram_top1_oc8051_idata_buff_199__2_,
         oc8051_ram_top1_oc8051_idata_buff_199__3_,
         oc8051_ram_top1_oc8051_idata_buff_199__4_,
         oc8051_ram_top1_oc8051_idata_buff_199__5_,
         oc8051_ram_top1_oc8051_idata_buff_199__6_,
         oc8051_ram_top1_oc8051_idata_buff_199__7_,
         oc8051_ram_top1_oc8051_idata_buff_198__0_,
         oc8051_ram_top1_oc8051_idata_buff_198__1_,
         oc8051_ram_top1_oc8051_idata_buff_198__2_,
         oc8051_ram_top1_oc8051_idata_buff_198__3_,
         oc8051_ram_top1_oc8051_idata_buff_198__4_,
         oc8051_ram_top1_oc8051_idata_buff_198__5_,
         oc8051_ram_top1_oc8051_idata_buff_198__6_,
         oc8051_ram_top1_oc8051_idata_buff_198__7_,
         oc8051_ram_top1_oc8051_idata_buff_195__0_,
         oc8051_ram_top1_oc8051_idata_buff_195__1_,
         oc8051_ram_top1_oc8051_idata_buff_195__2_,
         oc8051_ram_top1_oc8051_idata_buff_195__3_,
         oc8051_ram_top1_oc8051_idata_buff_195__4_,
         oc8051_ram_top1_oc8051_idata_buff_195__5_,
         oc8051_ram_top1_oc8051_idata_buff_195__6_,
         oc8051_ram_top1_oc8051_idata_buff_195__7_,
         oc8051_ram_top1_oc8051_idata_buff_194__0_,
         oc8051_ram_top1_oc8051_idata_buff_194__1_,
         oc8051_ram_top1_oc8051_idata_buff_194__2_,
         oc8051_ram_top1_oc8051_idata_buff_194__3_,
         oc8051_ram_top1_oc8051_idata_buff_194__4_,
         oc8051_ram_top1_oc8051_idata_buff_194__5_,
         oc8051_ram_top1_oc8051_idata_buff_194__6_,
         oc8051_ram_top1_oc8051_idata_buff_194__7_,
         oc8051_ram_top1_oc8051_idata_buff_63__0_,
         oc8051_ram_top1_oc8051_idata_buff_63__1_,
         oc8051_ram_top1_oc8051_idata_buff_63__2_,
         oc8051_ram_top1_oc8051_idata_buff_63__3_,
         oc8051_ram_top1_oc8051_idata_buff_63__4_,
         oc8051_ram_top1_oc8051_idata_buff_63__5_,
         oc8051_ram_top1_oc8051_idata_buff_63__6_,
         oc8051_ram_top1_oc8051_idata_buff_63__7_,
         oc8051_ram_top1_oc8051_idata_buff_62__0_,
         oc8051_ram_top1_oc8051_idata_buff_62__1_,
         oc8051_ram_top1_oc8051_idata_buff_62__2_,
         oc8051_ram_top1_oc8051_idata_buff_62__3_,
         oc8051_ram_top1_oc8051_idata_buff_62__4_,
         oc8051_ram_top1_oc8051_idata_buff_62__5_,
         oc8051_ram_top1_oc8051_idata_buff_62__6_,
         oc8051_ram_top1_oc8051_idata_buff_62__7_,
         oc8051_ram_top1_oc8051_idata_buff_61__0_,
         oc8051_ram_top1_oc8051_idata_buff_61__1_,
         oc8051_ram_top1_oc8051_idata_buff_61__2_,
         oc8051_ram_top1_oc8051_idata_buff_61__3_,
         oc8051_ram_top1_oc8051_idata_buff_61__4_,
         oc8051_ram_top1_oc8051_idata_buff_61__5_,
         oc8051_ram_top1_oc8051_idata_buff_61__6_,
         oc8051_ram_top1_oc8051_idata_buff_61__7_,
         oc8051_ram_top1_oc8051_idata_buff_60__0_,
         oc8051_ram_top1_oc8051_idata_buff_60__1_,
         oc8051_ram_top1_oc8051_idata_buff_60__2_,
         oc8051_ram_top1_oc8051_idata_buff_60__3_,
         oc8051_ram_top1_oc8051_idata_buff_60__4_,
         oc8051_ram_top1_oc8051_idata_buff_60__5_,
         oc8051_ram_top1_oc8051_idata_buff_60__6_,
         oc8051_ram_top1_oc8051_idata_buff_60__7_,
         oc8051_ram_top1_oc8051_idata_buff_59__0_,
         oc8051_ram_top1_oc8051_idata_buff_59__1_,
         oc8051_ram_top1_oc8051_idata_buff_59__2_,
         oc8051_ram_top1_oc8051_idata_buff_59__3_,
         oc8051_ram_top1_oc8051_idata_buff_59__4_,
         oc8051_ram_top1_oc8051_idata_buff_59__5_,
         oc8051_ram_top1_oc8051_idata_buff_59__6_,
         oc8051_ram_top1_oc8051_idata_buff_59__7_,
         oc8051_ram_top1_oc8051_idata_buff_58__0_,
         oc8051_ram_top1_oc8051_idata_buff_58__1_,
         oc8051_ram_top1_oc8051_idata_buff_58__2_,
         oc8051_ram_top1_oc8051_idata_buff_58__3_,
         oc8051_ram_top1_oc8051_idata_buff_58__4_,
         oc8051_ram_top1_oc8051_idata_buff_58__5_,
         oc8051_ram_top1_oc8051_idata_buff_58__6_,
         oc8051_ram_top1_oc8051_idata_buff_58__7_,
         oc8051_ram_top1_oc8051_idata_buff_57__0_,
         oc8051_ram_top1_oc8051_idata_buff_57__1_,
         oc8051_ram_top1_oc8051_idata_buff_57__2_,
         oc8051_ram_top1_oc8051_idata_buff_57__3_,
         oc8051_ram_top1_oc8051_idata_buff_57__4_,
         oc8051_ram_top1_oc8051_idata_buff_57__5_,
         oc8051_ram_top1_oc8051_idata_buff_57__6_,
         oc8051_ram_top1_oc8051_idata_buff_57__7_,
         oc8051_ram_top1_oc8051_idata_buff_56__0_,
         oc8051_ram_top1_oc8051_idata_buff_56__1_,
         oc8051_ram_top1_oc8051_idata_buff_56__2_,
         oc8051_ram_top1_oc8051_idata_buff_56__3_,
         oc8051_ram_top1_oc8051_idata_buff_56__4_,
         oc8051_ram_top1_oc8051_idata_buff_56__5_,
         oc8051_ram_top1_oc8051_idata_buff_56__6_,
         oc8051_ram_top1_oc8051_idata_buff_56__7_,
         oc8051_ram_top1_oc8051_idata_buff_53__0_,
         oc8051_ram_top1_oc8051_idata_buff_53__1_,
         oc8051_ram_top1_oc8051_idata_buff_53__2_,
         oc8051_ram_top1_oc8051_idata_buff_53__3_,
         oc8051_ram_top1_oc8051_idata_buff_53__4_,
         oc8051_ram_top1_oc8051_idata_buff_53__5_,
         oc8051_ram_top1_oc8051_idata_buff_53__6_,
         oc8051_ram_top1_oc8051_idata_buff_53__7_,
         oc8051_ram_top1_oc8051_idata_buff_52__0_,
         oc8051_ram_top1_oc8051_idata_buff_52__1_,
         oc8051_ram_top1_oc8051_idata_buff_52__2_,
         oc8051_ram_top1_oc8051_idata_buff_52__3_,
         oc8051_ram_top1_oc8051_idata_buff_52__4_,
         oc8051_ram_top1_oc8051_idata_buff_52__5_,
         oc8051_ram_top1_oc8051_idata_buff_52__6_,
         oc8051_ram_top1_oc8051_idata_buff_52__7_,
         oc8051_ram_top1_oc8051_idata_buff_49__0_,
         oc8051_ram_top1_oc8051_idata_buff_49__1_,
         oc8051_ram_top1_oc8051_idata_buff_49__2_,
         oc8051_ram_top1_oc8051_idata_buff_49__3_,
         oc8051_ram_top1_oc8051_idata_buff_49__4_,
         oc8051_ram_top1_oc8051_idata_buff_49__5_,
         oc8051_ram_top1_oc8051_idata_buff_49__6_,
         oc8051_ram_top1_oc8051_idata_buff_49__7_,
         oc8051_ram_top1_oc8051_idata_buff_48__0_,
         oc8051_ram_top1_oc8051_idata_buff_48__1_,
         oc8051_ram_top1_oc8051_idata_buff_48__2_,
         oc8051_ram_top1_oc8051_idata_buff_48__3_,
         oc8051_ram_top1_oc8051_idata_buff_48__4_,
         oc8051_ram_top1_oc8051_idata_buff_48__5_,
         oc8051_ram_top1_oc8051_idata_buff_48__6_,
         oc8051_ram_top1_oc8051_idata_buff_48__7_,
         oc8051_ram_top1_oc8051_idata_buff_47__0_,
         oc8051_ram_top1_oc8051_idata_buff_47__1_,
         oc8051_ram_top1_oc8051_idata_buff_47__2_,
         oc8051_ram_top1_oc8051_idata_buff_47__3_,
         oc8051_ram_top1_oc8051_idata_buff_47__4_,
         oc8051_ram_top1_oc8051_idata_buff_47__5_,
         oc8051_ram_top1_oc8051_idata_buff_47__6_,
         oc8051_ram_top1_oc8051_idata_buff_47__7_,
         oc8051_ram_top1_oc8051_idata_buff_46__0_,
         oc8051_ram_top1_oc8051_idata_buff_46__1_,
         oc8051_ram_top1_oc8051_idata_buff_46__2_,
         oc8051_ram_top1_oc8051_idata_buff_46__3_,
         oc8051_ram_top1_oc8051_idata_buff_46__4_,
         oc8051_ram_top1_oc8051_idata_buff_46__5_,
         oc8051_ram_top1_oc8051_idata_buff_46__6_,
         oc8051_ram_top1_oc8051_idata_buff_46__7_,
         oc8051_ram_top1_oc8051_idata_buff_45__0_,
         oc8051_ram_top1_oc8051_idata_buff_45__1_,
         oc8051_ram_top1_oc8051_idata_buff_45__2_,
         oc8051_ram_top1_oc8051_idata_buff_45__3_,
         oc8051_ram_top1_oc8051_idata_buff_45__4_,
         oc8051_ram_top1_oc8051_idata_buff_45__5_,
         oc8051_ram_top1_oc8051_idata_buff_45__6_,
         oc8051_ram_top1_oc8051_idata_buff_45__7_,
         oc8051_ram_top1_oc8051_idata_buff_44__0_,
         oc8051_ram_top1_oc8051_idata_buff_44__1_,
         oc8051_ram_top1_oc8051_idata_buff_44__2_,
         oc8051_ram_top1_oc8051_idata_buff_44__3_,
         oc8051_ram_top1_oc8051_idata_buff_44__4_,
         oc8051_ram_top1_oc8051_idata_buff_44__5_,
         oc8051_ram_top1_oc8051_idata_buff_44__6_,
         oc8051_ram_top1_oc8051_idata_buff_44__7_,
         oc8051_ram_top1_oc8051_idata_buff_43__0_,
         oc8051_ram_top1_oc8051_idata_buff_43__1_,
         oc8051_ram_top1_oc8051_idata_buff_43__2_,
         oc8051_ram_top1_oc8051_idata_buff_43__3_,
         oc8051_ram_top1_oc8051_idata_buff_43__4_,
         oc8051_ram_top1_oc8051_idata_buff_43__5_,
         oc8051_ram_top1_oc8051_idata_buff_43__6_,
         oc8051_ram_top1_oc8051_idata_buff_43__7_,
         oc8051_ram_top1_oc8051_idata_buff_42__0_,
         oc8051_ram_top1_oc8051_idata_buff_42__1_,
         oc8051_ram_top1_oc8051_idata_buff_42__2_,
         oc8051_ram_top1_oc8051_idata_buff_42__3_,
         oc8051_ram_top1_oc8051_idata_buff_42__4_,
         oc8051_ram_top1_oc8051_idata_buff_42__5_,
         oc8051_ram_top1_oc8051_idata_buff_42__6_,
         oc8051_ram_top1_oc8051_idata_buff_42__7_,
         oc8051_ram_top1_oc8051_idata_buff_41__0_,
         oc8051_ram_top1_oc8051_idata_buff_41__1_,
         oc8051_ram_top1_oc8051_idata_buff_41__2_,
         oc8051_ram_top1_oc8051_idata_buff_41__3_,
         oc8051_ram_top1_oc8051_idata_buff_41__4_,
         oc8051_ram_top1_oc8051_idata_buff_41__5_,
         oc8051_ram_top1_oc8051_idata_buff_41__6_,
         oc8051_ram_top1_oc8051_idata_buff_41__7_,
         oc8051_ram_top1_oc8051_idata_buff_40__0_,
         oc8051_ram_top1_oc8051_idata_buff_40__1_,
         oc8051_ram_top1_oc8051_idata_buff_40__2_,
         oc8051_ram_top1_oc8051_idata_buff_40__3_,
         oc8051_ram_top1_oc8051_idata_buff_40__4_,
         oc8051_ram_top1_oc8051_idata_buff_40__5_,
         oc8051_ram_top1_oc8051_idata_buff_40__6_,
         oc8051_ram_top1_oc8051_idata_buff_40__7_,
         oc8051_ram_top1_oc8051_idata_buff_39__0_,
         oc8051_ram_top1_oc8051_idata_buff_39__1_,
         oc8051_ram_top1_oc8051_idata_buff_39__2_,
         oc8051_ram_top1_oc8051_idata_buff_39__3_,
         oc8051_ram_top1_oc8051_idata_buff_39__4_,
         oc8051_ram_top1_oc8051_idata_buff_39__5_,
         oc8051_ram_top1_oc8051_idata_buff_39__6_,
         oc8051_ram_top1_oc8051_idata_buff_39__7_,
         oc8051_ram_top1_oc8051_idata_buff_38__0_,
         oc8051_ram_top1_oc8051_idata_buff_38__1_,
         oc8051_ram_top1_oc8051_idata_buff_38__2_,
         oc8051_ram_top1_oc8051_idata_buff_38__3_,
         oc8051_ram_top1_oc8051_idata_buff_38__4_,
         oc8051_ram_top1_oc8051_idata_buff_38__5_,
         oc8051_ram_top1_oc8051_idata_buff_38__6_,
         oc8051_ram_top1_oc8051_idata_buff_38__7_,
         oc8051_ram_top1_oc8051_idata_buff_35__0_,
         oc8051_ram_top1_oc8051_idata_buff_35__1_,
         oc8051_ram_top1_oc8051_idata_buff_35__2_,
         oc8051_ram_top1_oc8051_idata_buff_35__3_,
         oc8051_ram_top1_oc8051_idata_buff_35__4_,
         oc8051_ram_top1_oc8051_idata_buff_35__5_,
         oc8051_ram_top1_oc8051_idata_buff_35__6_,
         oc8051_ram_top1_oc8051_idata_buff_35__7_,
         oc8051_ram_top1_oc8051_idata_buff_34__0_,
         oc8051_ram_top1_oc8051_idata_buff_34__1_,
         oc8051_ram_top1_oc8051_idata_buff_34__2_,
         oc8051_ram_top1_oc8051_idata_buff_34__3_,
         oc8051_ram_top1_oc8051_idata_buff_34__4_,
         oc8051_ram_top1_oc8051_idata_buff_34__5_,
         oc8051_ram_top1_oc8051_idata_buff_34__6_,
         oc8051_ram_top1_oc8051_idata_buff_34__7_,
         oc8051_ram_top1_oc8051_idata_buff_31__0_,
         oc8051_ram_top1_oc8051_idata_buff_31__1_,
         oc8051_ram_top1_oc8051_idata_buff_31__2_,
         oc8051_ram_top1_oc8051_idata_buff_31__3_,
         oc8051_ram_top1_oc8051_idata_buff_31__4_,
         oc8051_ram_top1_oc8051_idata_buff_31__5_,
         oc8051_ram_top1_oc8051_idata_buff_31__6_,
         oc8051_ram_top1_oc8051_idata_buff_31__7_,
         oc8051_ram_top1_oc8051_idata_buff_30__0_,
         oc8051_ram_top1_oc8051_idata_buff_30__1_,
         oc8051_ram_top1_oc8051_idata_buff_30__2_,
         oc8051_ram_top1_oc8051_idata_buff_30__3_,
         oc8051_ram_top1_oc8051_idata_buff_30__4_,
         oc8051_ram_top1_oc8051_idata_buff_30__5_,
         oc8051_ram_top1_oc8051_idata_buff_30__6_,
         oc8051_ram_top1_oc8051_idata_buff_30__7_,
         oc8051_ram_top1_oc8051_idata_buff_29__0_,
         oc8051_ram_top1_oc8051_idata_buff_29__1_,
         oc8051_ram_top1_oc8051_idata_buff_29__2_,
         oc8051_ram_top1_oc8051_idata_buff_29__3_,
         oc8051_ram_top1_oc8051_idata_buff_29__4_,
         oc8051_ram_top1_oc8051_idata_buff_29__5_,
         oc8051_ram_top1_oc8051_idata_buff_29__6_,
         oc8051_ram_top1_oc8051_idata_buff_29__7_,
         oc8051_ram_top1_oc8051_idata_buff_28__0_,
         oc8051_ram_top1_oc8051_idata_buff_28__1_,
         oc8051_ram_top1_oc8051_idata_buff_28__2_,
         oc8051_ram_top1_oc8051_idata_buff_28__3_,
         oc8051_ram_top1_oc8051_idata_buff_28__4_,
         oc8051_ram_top1_oc8051_idata_buff_28__5_,
         oc8051_ram_top1_oc8051_idata_buff_28__6_,
         oc8051_ram_top1_oc8051_idata_buff_28__7_,
         oc8051_ram_top1_oc8051_idata_buff_27__0_,
         oc8051_ram_top1_oc8051_idata_buff_27__1_,
         oc8051_ram_top1_oc8051_idata_buff_27__2_,
         oc8051_ram_top1_oc8051_idata_buff_27__3_,
         oc8051_ram_top1_oc8051_idata_buff_27__4_,
         oc8051_ram_top1_oc8051_idata_buff_27__5_,
         oc8051_ram_top1_oc8051_idata_buff_27__6_,
         oc8051_ram_top1_oc8051_idata_buff_27__7_,
         oc8051_ram_top1_oc8051_idata_buff_26__0_,
         oc8051_ram_top1_oc8051_idata_buff_26__1_,
         oc8051_ram_top1_oc8051_idata_buff_26__2_,
         oc8051_ram_top1_oc8051_idata_buff_26__3_,
         oc8051_ram_top1_oc8051_idata_buff_26__4_,
         oc8051_ram_top1_oc8051_idata_buff_26__5_,
         oc8051_ram_top1_oc8051_idata_buff_26__6_,
         oc8051_ram_top1_oc8051_idata_buff_26__7_,
         oc8051_ram_top1_oc8051_idata_buff_25__0_,
         oc8051_ram_top1_oc8051_idata_buff_25__1_,
         oc8051_ram_top1_oc8051_idata_buff_25__2_,
         oc8051_ram_top1_oc8051_idata_buff_25__3_,
         oc8051_ram_top1_oc8051_idata_buff_25__4_,
         oc8051_ram_top1_oc8051_idata_buff_25__5_,
         oc8051_ram_top1_oc8051_idata_buff_25__6_,
         oc8051_ram_top1_oc8051_idata_buff_25__7_,
         oc8051_ram_top1_oc8051_idata_buff_24__0_,
         oc8051_ram_top1_oc8051_idata_buff_24__1_,
         oc8051_ram_top1_oc8051_idata_buff_24__2_,
         oc8051_ram_top1_oc8051_idata_buff_24__3_,
         oc8051_ram_top1_oc8051_idata_buff_24__4_,
         oc8051_ram_top1_oc8051_idata_buff_24__5_,
         oc8051_ram_top1_oc8051_idata_buff_24__6_,
         oc8051_ram_top1_oc8051_idata_buff_24__7_,
         oc8051_ram_top1_oc8051_idata_buff_23__0_,
         oc8051_ram_top1_oc8051_idata_buff_23__1_,
         oc8051_ram_top1_oc8051_idata_buff_23__2_,
         oc8051_ram_top1_oc8051_idata_buff_23__3_,
         oc8051_ram_top1_oc8051_idata_buff_23__4_,
         oc8051_ram_top1_oc8051_idata_buff_23__5_,
         oc8051_ram_top1_oc8051_idata_buff_23__6_,
         oc8051_ram_top1_oc8051_idata_buff_23__7_,
         oc8051_ram_top1_oc8051_idata_buff_22__0_,
         oc8051_ram_top1_oc8051_idata_buff_22__1_,
         oc8051_ram_top1_oc8051_idata_buff_22__2_,
         oc8051_ram_top1_oc8051_idata_buff_22__3_,
         oc8051_ram_top1_oc8051_idata_buff_22__4_,
         oc8051_ram_top1_oc8051_idata_buff_22__5_,
         oc8051_ram_top1_oc8051_idata_buff_22__6_,
         oc8051_ram_top1_oc8051_idata_buff_22__7_,
         oc8051_ram_top1_oc8051_idata_buff_21__0_,
         oc8051_ram_top1_oc8051_idata_buff_21__1_,
         oc8051_ram_top1_oc8051_idata_buff_21__2_,
         oc8051_ram_top1_oc8051_idata_buff_21__3_,
         oc8051_ram_top1_oc8051_idata_buff_21__4_,
         oc8051_ram_top1_oc8051_idata_buff_21__5_,
         oc8051_ram_top1_oc8051_idata_buff_21__6_,
         oc8051_ram_top1_oc8051_idata_buff_21__7_,
         oc8051_ram_top1_oc8051_idata_buff_20__0_,
         oc8051_ram_top1_oc8051_idata_buff_20__1_,
         oc8051_ram_top1_oc8051_idata_buff_20__2_,
         oc8051_ram_top1_oc8051_idata_buff_20__3_,
         oc8051_ram_top1_oc8051_idata_buff_20__4_,
         oc8051_ram_top1_oc8051_idata_buff_20__5_,
         oc8051_ram_top1_oc8051_idata_buff_20__6_,
         oc8051_ram_top1_oc8051_idata_buff_20__7_,
         oc8051_ram_top1_oc8051_idata_buff_19__0_,
         oc8051_ram_top1_oc8051_idata_buff_19__1_,
         oc8051_ram_top1_oc8051_idata_buff_19__2_,
         oc8051_ram_top1_oc8051_idata_buff_19__3_,
         oc8051_ram_top1_oc8051_idata_buff_19__4_,
         oc8051_ram_top1_oc8051_idata_buff_19__5_,
         oc8051_ram_top1_oc8051_idata_buff_19__6_,
         oc8051_ram_top1_oc8051_idata_buff_19__7_,
         oc8051_ram_top1_oc8051_idata_buff_18__0_,
         oc8051_ram_top1_oc8051_idata_buff_18__1_,
         oc8051_ram_top1_oc8051_idata_buff_18__2_,
         oc8051_ram_top1_oc8051_idata_buff_18__3_,
         oc8051_ram_top1_oc8051_idata_buff_18__4_,
         oc8051_ram_top1_oc8051_idata_buff_18__5_,
         oc8051_ram_top1_oc8051_idata_buff_18__6_,
         oc8051_ram_top1_oc8051_idata_buff_18__7_,
         oc8051_ram_top1_oc8051_idata_buff_17__0_,
         oc8051_ram_top1_oc8051_idata_buff_17__1_,
         oc8051_ram_top1_oc8051_idata_buff_17__2_,
         oc8051_ram_top1_oc8051_idata_buff_17__3_,
         oc8051_ram_top1_oc8051_idata_buff_17__4_,
         oc8051_ram_top1_oc8051_idata_buff_17__5_,
         oc8051_ram_top1_oc8051_idata_buff_17__6_,
         oc8051_ram_top1_oc8051_idata_buff_17__7_,
         oc8051_ram_top1_oc8051_idata_buff_16__0_,
         oc8051_ram_top1_oc8051_idata_buff_16__1_,
         oc8051_ram_top1_oc8051_idata_buff_16__2_,
         oc8051_ram_top1_oc8051_idata_buff_16__3_,
         oc8051_ram_top1_oc8051_idata_buff_16__4_,
         oc8051_ram_top1_oc8051_idata_buff_16__5_,
         oc8051_ram_top1_oc8051_idata_buff_16__6_,
         oc8051_ram_top1_oc8051_idata_buff_16__7_,
         oc8051_ram_top1_oc8051_idata_buff_13__0_,
         oc8051_ram_top1_oc8051_idata_buff_13__1_,
         oc8051_ram_top1_oc8051_idata_buff_13__2_,
         oc8051_ram_top1_oc8051_idata_buff_13__3_,
         oc8051_ram_top1_oc8051_idata_buff_13__4_,
         oc8051_ram_top1_oc8051_idata_buff_13__5_,
         oc8051_ram_top1_oc8051_idata_buff_13__6_,
         oc8051_ram_top1_oc8051_idata_buff_13__7_,
         oc8051_ram_top1_oc8051_idata_buff_12__0_,
         oc8051_ram_top1_oc8051_idata_buff_12__1_,
         oc8051_ram_top1_oc8051_idata_buff_12__2_,
         oc8051_ram_top1_oc8051_idata_buff_12__3_,
         oc8051_ram_top1_oc8051_idata_buff_12__4_,
         oc8051_ram_top1_oc8051_idata_buff_12__5_,
         oc8051_ram_top1_oc8051_idata_buff_12__6_,
         oc8051_ram_top1_oc8051_idata_buff_12__7_,
         oc8051_ram_top1_oc8051_idata_buff_11__0_,
         oc8051_ram_top1_oc8051_idata_buff_11__1_,
         oc8051_ram_top1_oc8051_idata_buff_11__2_,
         oc8051_ram_top1_oc8051_idata_buff_11__3_,
         oc8051_ram_top1_oc8051_idata_buff_11__4_,
         oc8051_ram_top1_oc8051_idata_buff_11__5_,
         oc8051_ram_top1_oc8051_idata_buff_11__6_,
         oc8051_ram_top1_oc8051_idata_buff_11__7_,
         oc8051_ram_top1_oc8051_idata_buff_10__0_,
         oc8051_ram_top1_oc8051_idata_buff_10__1_,
         oc8051_ram_top1_oc8051_idata_buff_10__2_,
         oc8051_ram_top1_oc8051_idata_buff_10__3_,
         oc8051_ram_top1_oc8051_idata_buff_10__4_,
         oc8051_ram_top1_oc8051_idata_buff_10__5_,
         oc8051_ram_top1_oc8051_idata_buff_10__6_,
         oc8051_ram_top1_oc8051_idata_buff_10__7_,
         oc8051_ram_top1_oc8051_idata_buff_7__0_,
         oc8051_ram_top1_oc8051_idata_buff_7__1_,
         oc8051_ram_top1_oc8051_idata_buff_7__2_,
         oc8051_ram_top1_oc8051_idata_buff_7__3_,
         oc8051_ram_top1_oc8051_idata_buff_7__4_,
         oc8051_ram_top1_oc8051_idata_buff_7__5_,
         oc8051_ram_top1_oc8051_idata_buff_7__6_,
         oc8051_ram_top1_oc8051_idata_buff_7__7_,
         oc8051_ram_top1_oc8051_idata_buff_6__0_,
         oc8051_ram_top1_oc8051_idata_buff_6__1_,
         oc8051_ram_top1_oc8051_idata_buff_6__2_,
         oc8051_ram_top1_oc8051_idata_buff_6__3_,
         oc8051_ram_top1_oc8051_idata_buff_6__4_,
         oc8051_ram_top1_oc8051_idata_buff_6__5_,
         oc8051_ram_top1_oc8051_idata_buff_6__6_,
         oc8051_ram_top1_oc8051_idata_buff_6__7_,
         oc8051_ram_top1_oc8051_idata_buff_3__0_,
         oc8051_ram_top1_oc8051_idata_buff_3__1_,
         oc8051_ram_top1_oc8051_idata_buff_3__2_,
         oc8051_ram_top1_oc8051_idata_buff_3__3_,
         oc8051_ram_top1_oc8051_idata_buff_3__4_,
         oc8051_ram_top1_oc8051_idata_buff_3__5_,
         oc8051_ram_top1_oc8051_idata_buff_3__6_,
         oc8051_ram_top1_oc8051_idata_buff_3__7_,
         oc8051_ram_top1_oc8051_idata_buff_2__0_,
         oc8051_ram_top1_oc8051_idata_buff_2__1_,
         oc8051_ram_top1_oc8051_idata_buff_2__2_,
         oc8051_ram_top1_oc8051_idata_buff_2__3_,
         oc8051_ram_top1_oc8051_idata_buff_2__4_,
         oc8051_ram_top1_oc8051_idata_buff_2__5_,
         oc8051_ram_top1_oc8051_idata_buff_2__6_,
         oc8051_ram_top1_oc8051_idata_buff_2__7_, oc8051_alu_src_sel1_n61,
         oc8051_alu_src_sel1_n60, oc8051_alu_src_sel1_n59,
         oc8051_alu_src_sel1_n58, oc8051_alu_src_sel1_n57,
         oc8051_alu_src_sel1_n56, oc8051_alu_src_sel1_n55,
         oc8051_alu_src_sel1_n54, oc8051_alu_src_sel1_n53,
         oc8051_alu_src_sel1_n52, oc8051_alu_src_sel1_n51,
         oc8051_alu_src_sel1_n50, oc8051_alu_src_sel1_n49,
         oc8051_alu_src_sel1_n48, oc8051_alu_src_sel1_n47,
         oc8051_alu_src_sel1_n46, oc8051_alu_src_sel1_n45,
         oc8051_alu_src_sel1_n44, oc8051_alu_src_sel1_n43,
         oc8051_alu_src_sel1_n42, oc8051_alu_src_sel1_n41,
         oc8051_alu_src_sel1_n40, oc8051_alu_src_sel1_n39,
         oc8051_alu_src_sel1_n38, oc8051_alu_src_sel1_n37,
         oc8051_alu_src_sel1_n36, oc8051_alu_src_sel1_n35,
         oc8051_alu_src_sel1_n34, oc8051_alu_src_sel1_n33,
         oc8051_alu_src_sel1_n32, oc8051_alu_src_sel1_n31,
         oc8051_alu_src_sel1_n30, oc8051_alu_src_sel1_n29,
         oc8051_alu_src_sel1_n28, oc8051_alu_src_sel1_n27,
         oc8051_alu_src_sel1_n26, oc8051_alu_src_sel1_n25,
         oc8051_alu_src_sel1_n24, oc8051_alu_src_sel1_n23,
         oc8051_alu_src_sel1_n22, oc8051_alu_src_sel1_n21,
         oc8051_alu_src_sel1_n20, oc8051_alu_src_sel1_n19,
         oc8051_alu_src_sel1_n18, oc8051_alu_src_sel1_n17,
         oc8051_alu_src_sel1_n16, oc8051_alu_src_sel1_n15,
         oc8051_alu_src_sel1_n14, oc8051_alu_src_sel1_n13,
         oc8051_alu_src_sel1_n12, oc8051_alu_src_sel1_n11,
         oc8051_alu_src_sel1_n10, oc8051_alu_src_sel1_n9,
         oc8051_alu_src_sel1_n8, oc8051_alu_src_sel1_n7,
         oc8051_alu_src_sel1_n6, oc8051_alu_src_sel1_n5,
         oc8051_alu_src_sel1_n4, oc8051_alu_src_sel1_n3,
         oc8051_alu_src_sel1_n2, oc8051_alu_src_sel1_n1,
         oc8051_alu_src_sel1_op2_r_0_, oc8051_alu_src_sel1_op2_r_1_,
         oc8051_alu_src_sel1_op2_r_2_, oc8051_alu_src_sel1_op2_r_3_,
         oc8051_alu_src_sel1_op2_r_4_, oc8051_alu_src_sel1_op2_r_5_,
         oc8051_alu_src_sel1_op2_r_6_, oc8051_alu_src_sel1_op2_r_7_,
         oc8051_comp1_n10, oc8051_comp1_n9, oc8051_comp1_n8, oc8051_comp1_n7,
         oc8051_comp1_n6, oc8051_comp1_n5, oc8051_comp1_n4, oc8051_comp1_n3,
         oc8051_comp1_n2, oc8051_comp1_n1, oc8051_rom1_data_o_0_,
         oc8051_rom1_ea_int, oc8051_cy_select1_n1, oc8051_indi_addr1_n98,
         oc8051_indi_addr1_n97, oc8051_indi_addr1_n96, oc8051_indi_addr1_n95,
         oc8051_indi_addr1_n94, oc8051_indi_addr1_n93, oc8051_indi_addr1_n92,
         oc8051_indi_addr1_n27, oc8051_indi_addr1_n26, oc8051_indi_addr1_n25,
         oc8051_indi_addr1_n24, oc8051_indi_addr1_n23, oc8051_indi_addr1_n22,
         oc8051_indi_addr1_n21, oc8051_indi_addr1_n20, oc8051_indi_addr1_n19,
         oc8051_indi_addr1_n18, oc8051_indi_addr1_n17, oc8051_indi_addr1_n16,
         oc8051_indi_addr1_n15, oc8051_indi_addr1_n14, oc8051_indi_addr1_n13,
         oc8051_indi_addr1_n12, oc8051_indi_addr1_n11, oc8051_indi_addr1_n10,
         oc8051_indi_addr1_n9, oc8051_indi_addr1_n8, oc8051_indi_addr1_n7,
         oc8051_indi_addr1_n6, oc8051_indi_addr1_n5, oc8051_indi_addr1_n4,
         oc8051_indi_addr1_n3, oc8051_indi_addr1_n2, oc8051_indi_addr1_n1,
         oc8051_indi_addr1_n91, oc8051_indi_addr1_n90, oc8051_indi_addr1_n89,
         oc8051_indi_addr1_n88, oc8051_indi_addr1_n87, oc8051_indi_addr1_n86,
         oc8051_indi_addr1_n85, oc8051_indi_addr1_n84, oc8051_indi_addr1_n83,
         oc8051_indi_addr1_n82, oc8051_indi_addr1_n81, oc8051_indi_addr1_n80,
         oc8051_indi_addr1_n79, oc8051_indi_addr1_n78, oc8051_indi_addr1_n77,
         oc8051_indi_addr1_n76, oc8051_indi_addr1_n75, oc8051_indi_addr1_n74,
         oc8051_indi_addr1_n73, oc8051_indi_addr1_n72, oc8051_indi_addr1_n71,
         oc8051_indi_addr1_n70, oc8051_indi_addr1_n69, oc8051_indi_addr1_n68,
         oc8051_indi_addr1_n67, oc8051_indi_addr1_n66, oc8051_indi_addr1_n65,
         oc8051_indi_addr1_n64, oc8051_indi_addr1_n63, oc8051_indi_addr1_n62,
         oc8051_indi_addr1_n61, oc8051_indi_addr1_n60, oc8051_indi_addr1_n59,
         oc8051_indi_addr1_n58, oc8051_indi_addr1_n57, oc8051_indi_addr1_n56,
         oc8051_indi_addr1_n55, oc8051_indi_addr1_n54, oc8051_indi_addr1_n53,
         oc8051_indi_addr1_n52, oc8051_indi_addr1_n51, oc8051_indi_addr1_n50,
         oc8051_indi_addr1_n49, oc8051_indi_addr1_n48, oc8051_indi_addr1_n47,
         oc8051_indi_addr1_n46, oc8051_indi_addr1_n45, oc8051_indi_addr1_n44,
         oc8051_indi_addr1_n43, oc8051_indi_addr1_n42, oc8051_indi_addr1_n41,
         oc8051_indi_addr1_n40, oc8051_indi_addr1_n39, oc8051_indi_addr1_n38,
         oc8051_indi_addr1_n37, oc8051_indi_addr1_n36, oc8051_indi_addr1_n35,
         oc8051_indi_addr1_n34, oc8051_indi_addr1_n33, oc8051_indi_addr1_n32,
         oc8051_indi_addr1_n31, oc8051_indi_addr1_n30, oc8051_indi_addr1_n29,
         oc8051_indi_addr1_n28, oc8051_indi_addr1_n106, oc8051_indi_addr1_n105,
         oc8051_indi_addr1_n104, oc8051_indi_addr1_n103,
         oc8051_indi_addr1_n102, oc8051_indi_addr1_n101,
         oc8051_indi_addr1_n100, oc8051_indi_addr1_n99,
         oc8051_indi_addr1_wr_bit_r, oc8051_indi_addr1_buff_7__0_,
         oc8051_indi_addr1_buff_7__1_, oc8051_indi_addr1_buff_7__2_,
         oc8051_indi_addr1_buff_7__3_, oc8051_indi_addr1_buff_7__4_,
         oc8051_indi_addr1_buff_7__5_, oc8051_indi_addr1_buff_7__6_,
         oc8051_indi_addr1_buff_7__7_, oc8051_indi_addr1_buff_6__0_,
         oc8051_indi_addr1_buff_6__1_, oc8051_indi_addr1_buff_6__2_,
         oc8051_indi_addr1_buff_6__3_, oc8051_indi_addr1_buff_6__4_,
         oc8051_indi_addr1_buff_6__5_, oc8051_indi_addr1_buff_6__6_,
         oc8051_indi_addr1_buff_6__7_, oc8051_indi_addr1_buff_5__0_,
         oc8051_indi_addr1_buff_5__1_, oc8051_indi_addr1_buff_5__2_,
         oc8051_indi_addr1_buff_5__3_, oc8051_indi_addr1_buff_5__4_,
         oc8051_indi_addr1_buff_5__5_, oc8051_indi_addr1_buff_5__6_,
         oc8051_indi_addr1_buff_5__7_, oc8051_indi_addr1_buff_4__0_,
         oc8051_indi_addr1_buff_4__1_, oc8051_indi_addr1_buff_4__2_,
         oc8051_indi_addr1_buff_4__3_, oc8051_indi_addr1_buff_4__4_,
         oc8051_indi_addr1_buff_4__5_, oc8051_indi_addr1_buff_4__6_,
         oc8051_indi_addr1_buff_4__7_, oc8051_indi_addr1_buff_3__0_,
         oc8051_indi_addr1_buff_3__1_, oc8051_indi_addr1_buff_3__2_,
         oc8051_indi_addr1_buff_3__3_, oc8051_indi_addr1_buff_3__4_,
         oc8051_indi_addr1_buff_3__5_, oc8051_indi_addr1_buff_3__6_,
         oc8051_indi_addr1_buff_3__7_, oc8051_indi_addr1_buff_2__0_,
         oc8051_indi_addr1_buff_2__1_, oc8051_indi_addr1_buff_2__2_,
         oc8051_indi_addr1_buff_2__3_, oc8051_indi_addr1_buff_2__4_,
         oc8051_indi_addr1_buff_2__5_, oc8051_indi_addr1_buff_2__6_,
         oc8051_indi_addr1_buff_2__7_, oc8051_indi_addr1_buff_1__0_,
         oc8051_indi_addr1_buff_1__1_, oc8051_indi_addr1_buff_1__2_,
         oc8051_indi_addr1_buff_1__3_, oc8051_indi_addr1_buff_1__4_,
         oc8051_indi_addr1_buff_1__5_, oc8051_indi_addr1_buff_1__6_,
         oc8051_indi_addr1_buff_1__7_, oc8051_indi_addr1_buff_0__0_,
         oc8051_indi_addr1_buff_0__1_, oc8051_indi_addr1_buff_0__2_,
         oc8051_indi_addr1_buff_0__3_, oc8051_indi_addr1_buff_0__4_,
         oc8051_indi_addr1_buff_0__5_, oc8051_indi_addr1_buff_0__6_,
         oc8051_indi_addr1_buff_0__7_, oc8051_memory_interface1_n813,
         oc8051_memory_interface1_n804, oc8051_memory_interface1_n803,
         oc8051_memory_interface1_n802, oc8051_memory_interface1_n801,
         oc8051_memory_interface1_n800, oc8051_memory_interface1_n799,
         oc8051_memory_interface1_n798, oc8051_memory_interface1_n797,
         oc8051_memory_interface1_n796, oc8051_memory_interface1_n795,
         oc8051_memory_interface1_n794, oc8051_memory_interface1_n793,
         oc8051_memory_interface1_n792, oc8051_memory_interface1_n791,
         oc8051_memory_interface1_n790, oc8051_memory_interface1_n789,
         oc8051_memory_interface1_n772, oc8051_memory_interface1_n771,
         oc8051_memory_interface1_n770, oc8051_memory_interface1_n769,
         oc8051_memory_interface1_n768, oc8051_memory_interface1_n767,
         oc8051_memory_interface1_n766, oc8051_memory_interface1_n765,
         oc8051_memory_interface1_n764, oc8051_memory_interface1_n763,
         oc8051_memory_interface1_n762, oc8051_memory_interface1_n761,
         oc8051_memory_interface1_n760, oc8051_memory_interface1_n759,
         oc8051_memory_interface1_n758, oc8051_memory_interface1_n757,
         oc8051_memory_interface1_n756, oc8051_memory_interface1_n755,
         oc8051_memory_interface1_n754, oc8051_memory_interface1_n753,
         oc8051_memory_interface1_n752, oc8051_memory_interface1_n751,
         oc8051_memory_interface1_n750, oc8051_memory_interface1_n749,
         oc8051_memory_interface1_n748, oc8051_memory_interface1_n747,
         oc8051_memory_interface1_n746, oc8051_memory_interface1_n745,
         oc8051_memory_interface1_n744, oc8051_memory_interface1_n743,
         oc8051_memory_interface1_n742, oc8051_memory_interface1_n741,
         oc8051_memory_interface1_n740, oc8051_memory_interface1_n739,
         oc8051_memory_interface1_n738, oc8051_memory_interface1_n737,
         oc8051_memory_interface1_n736, oc8051_memory_interface1_n735,
         oc8051_memory_interface1_n734, oc8051_memory_interface1_n733,
         oc8051_memory_interface1_n732, oc8051_memory_interface1_n731,
         oc8051_memory_interface1_n730, oc8051_memory_interface1_n729,
         oc8051_memory_interface1_n728, oc8051_memory_interface1_n727,
         oc8051_memory_interface1_n726, oc8051_memory_interface1_n725,
         oc8051_memory_interface1_n724, oc8051_memory_interface1_n723,
         oc8051_memory_interface1_n722, oc8051_memory_interface1_n721,
         oc8051_memory_interface1_n720, oc8051_memory_interface1_n719,
         oc8051_memory_interface1_n718, oc8051_memory_interface1_n717,
         oc8051_memory_interface1_n716, oc8051_memory_interface1_n715,
         oc8051_memory_interface1_n714, oc8051_memory_interface1_n713,
         oc8051_memory_interface1_n712, oc8051_memory_interface1_n711,
         oc8051_memory_interface1_n710, oc8051_memory_interface1_n709,
         oc8051_memory_interface1_n708, oc8051_memory_interface1_n707,
         oc8051_memory_interface1_n706, oc8051_memory_interface1_n705,
         oc8051_memory_interface1_n704, oc8051_memory_interface1_n703,
         oc8051_memory_interface1_n702, oc8051_memory_interface1_n701,
         oc8051_memory_interface1_n700, oc8051_memory_interface1_n699,
         oc8051_memory_interface1_n698, oc8051_memory_interface1_n697,
         oc8051_memory_interface1_n696, oc8051_memory_interface1_n695,
         oc8051_memory_interface1_n694, oc8051_memory_interface1_n693,
         oc8051_memory_interface1_n692, oc8051_memory_interface1_n691,
         oc8051_memory_interface1_n690, oc8051_memory_interface1_n689,
         oc8051_memory_interface1_n688, oc8051_memory_interface1_n687,
         oc8051_memory_interface1_n686, oc8051_memory_interface1_n685,
         oc8051_memory_interface1_n684, oc8051_memory_interface1_n683,
         oc8051_memory_interface1_n682, oc8051_memory_interface1_n681,
         oc8051_memory_interface1_n680, oc8051_memory_interface1_n679,
         oc8051_memory_interface1_n678, oc8051_memory_interface1_n677,
         oc8051_memory_interface1_n676, oc8051_memory_interface1_n675,
         oc8051_memory_interface1_n674, oc8051_memory_interface1_n673,
         oc8051_memory_interface1_n672, oc8051_memory_interface1_n671,
         oc8051_memory_interface1_n670, oc8051_memory_interface1_n669,
         oc8051_memory_interface1_n668, oc8051_memory_interface1_n667,
         oc8051_memory_interface1_n666, oc8051_memory_interface1_n665,
         oc8051_memory_interface1_n664, oc8051_memory_interface1_n663,
         oc8051_memory_interface1_n662, oc8051_memory_interface1_n661,
         oc8051_memory_interface1_n660, oc8051_memory_interface1_n659,
         oc8051_memory_interface1_n658, oc8051_memory_interface1_n657,
         oc8051_memory_interface1_n656, oc8051_memory_interface1_n655,
         oc8051_memory_interface1_n654, oc8051_memory_interface1_n653,
         oc8051_memory_interface1_n652, oc8051_memory_interface1_n651,
         oc8051_memory_interface1_n650, oc8051_memory_interface1_n649,
         oc8051_memory_interface1_n648, oc8051_memory_interface1_n647,
         oc8051_memory_interface1_n646, oc8051_memory_interface1_n645,
         oc8051_memory_interface1_n644, oc8051_memory_interface1_n643,
         oc8051_memory_interface1_n642, oc8051_memory_interface1_n641,
         oc8051_memory_interface1_n640, oc8051_memory_interface1_n639,
         oc8051_memory_interface1_n638, oc8051_memory_interface1_n637,
         oc8051_memory_interface1_n636, oc8051_memory_interface1_n635,
         oc8051_memory_interface1_n634, oc8051_memory_interface1_n633,
         oc8051_memory_interface1_n632, oc8051_memory_interface1_n631,
         oc8051_memory_interface1_n630, oc8051_memory_interface1_n629,
         oc8051_memory_interface1_n628, oc8051_memory_interface1_n627,
         oc8051_memory_interface1_n626, oc8051_memory_interface1_n625,
         oc8051_memory_interface1_n624, oc8051_memory_interface1_n623,
         oc8051_memory_interface1_n622, oc8051_memory_interface1_n621,
         oc8051_memory_interface1_n620, oc8051_memory_interface1_n619,
         oc8051_memory_interface1_n618, oc8051_memory_interface1_n617,
         oc8051_memory_interface1_n616, oc8051_memory_interface1_n615,
         oc8051_memory_interface1_n614, oc8051_memory_interface1_n613,
         oc8051_memory_interface1_n612, oc8051_memory_interface1_n611,
         oc8051_memory_interface1_n610, oc8051_memory_interface1_n609,
         oc8051_memory_interface1_n608, oc8051_memory_interface1_n607,
         oc8051_memory_interface1_n606, oc8051_memory_interface1_n605,
         oc8051_memory_interface1_n604, oc8051_memory_interface1_n603,
         oc8051_memory_interface1_n602, oc8051_memory_interface1_n601,
         oc8051_memory_interface1_n600, oc8051_memory_interface1_n599,
         oc8051_memory_interface1_n598, oc8051_memory_interface1_n597,
         oc8051_memory_interface1_n596, oc8051_memory_interface1_n595,
         oc8051_memory_interface1_n594, oc8051_memory_interface1_n593,
         oc8051_memory_interface1_n592, oc8051_memory_interface1_n591,
         oc8051_memory_interface1_n590, oc8051_memory_interface1_n589,
         oc8051_memory_interface1_n588, oc8051_memory_interface1_n587,
         oc8051_memory_interface1_n586, oc8051_memory_interface1_n585,
         oc8051_memory_interface1_n556, oc8051_memory_interface1_n554,
         oc8051_memory_interface1_n552, oc8051_memory_interface1_n550,
         oc8051_memory_interface1_n548, oc8051_memory_interface1_n546,
         oc8051_memory_interface1_n544, oc8051_memory_interface1_n542,
         oc8051_memory_interface1_n458, oc8051_memory_interface1_n457,
         oc8051_memory_interface1_n456, oc8051_memory_interface1_n439,
         oc8051_memory_interface1_n438, oc8051_memory_interface1_n437,
         oc8051_memory_interface1_n436, oc8051_memory_interface1_n435,
         oc8051_memory_interface1_n434, oc8051_memory_interface1_n433,
         oc8051_memory_interface1_n432, oc8051_memory_interface1_n415,
         oc8051_memory_interface1_n414, oc8051_memory_interface1_n413,
         oc8051_memory_interface1_n412, oc8051_memory_interface1_n411,
         oc8051_memory_interface1_n410, oc8051_memory_interface1_n409,
         oc8051_memory_interface1_n408, oc8051_memory_interface1_n407,
         oc8051_memory_interface1_n406, oc8051_memory_interface1_n405,
         oc8051_memory_interface1_n404, oc8051_memory_interface1_n403,
         oc8051_memory_interface1_n402, oc8051_memory_interface1_n401,
         oc8051_memory_interface1_n400, oc8051_memory_interface1_n391,
         oc8051_memory_interface1_n390, oc8051_memory_interface1_n389,
         oc8051_memory_interface1_n388, oc8051_memory_interface1_n387,
         oc8051_memory_interface1_n386, oc8051_memory_interface1_n385,
         oc8051_memory_interface1_n384, oc8051_memory_interface1_n383,
         oc8051_memory_interface1_n382, oc8051_memory_interface1_n381,
         oc8051_memory_interface1_n380, oc8051_memory_interface1_n379,
         oc8051_memory_interface1_n378, oc8051_memory_interface1_n377,
         oc8051_memory_interface1_n376, oc8051_memory_interface1_n375,
         oc8051_memory_interface1_n374, oc8051_memory_interface1_n373,
         oc8051_memory_interface1_n372, oc8051_memory_interface1_n371,
         oc8051_memory_interface1_n370, oc8051_memory_interface1_n369,
         oc8051_memory_interface1_n368, oc8051_memory_interface1_n367,
         oc8051_memory_interface1_n366, oc8051_memory_interface1_n365,
         oc8051_memory_interface1_n364, oc8051_memory_interface1_n363,
         oc8051_memory_interface1_n362, oc8051_memory_interface1_n361,
         oc8051_memory_interface1_n360, oc8051_memory_interface1_n359,
         oc8051_memory_interface1_n358, oc8051_memory_interface1_n357,
         oc8051_memory_interface1_n356, oc8051_memory_interface1_n355,
         oc8051_memory_interface1_n354, oc8051_memory_interface1_n353,
         oc8051_memory_interface1_n352, oc8051_memory_interface1_n351,
         oc8051_memory_interface1_n350, oc8051_memory_interface1_n349,
         oc8051_memory_interface1_n348, oc8051_memory_interface1_n347,
         oc8051_memory_interface1_n346, oc8051_memory_interface1_n345,
         oc8051_memory_interface1_n344, oc8051_memory_interface1_n343,
         oc8051_memory_interface1_n342, oc8051_memory_interface1_n341,
         oc8051_memory_interface1_n340, oc8051_memory_interface1_n339,
         oc8051_memory_interface1_n338, oc8051_memory_interface1_n337,
         oc8051_memory_interface1_n336, oc8051_memory_interface1_n335,
         oc8051_memory_interface1_n334, oc8051_memory_interface1_n333,
         oc8051_memory_interface1_n332, oc8051_memory_interface1_n331,
         oc8051_memory_interface1_n330, oc8051_memory_interface1_n329,
         oc8051_memory_interface1_n328, oc8051_memory_interface1_n327,
         oc8051_memory_interface1_n326, oc8051_memory_interface1_n325,
         oc8051_memory_interface1_n324, oc8051_memory_interface1_n323,
         oc8051_memory_interface1_n322, oc8051_memory_interface1_n321,
         oc8051_memory_interface1_n320, oc8051_memory_interface1_n319,
         oc8051_memory_interface1_n318, oc8051_memory_interface1_n317,
         oc8051_memory_interface1_n316, oc8051_memory_interface1_n315,
         oc8051_memory_interface1_n314, oc8051_memory_interface1_n313,
         oc8051_memory_interface1_n312, oc8051_memory_interface1_n311,
         oc8051_memory_interface1_n310, oc8051_memory_interface1_n309,
         oc8051_memory_interface1_n308, oc8051_memory_interface1_n307,
         oc8051_memory_interface1_n306, oc8051_memory_interface1_n305,
         oc8051_memory_interface1_n304, oc8051_memory_interface1_n303,
         oc8051_memory_interface1_n302, oc8051_memory_interface1_n301,
         oc8051_memory_interface1_n300, oc8051_memory_interface1_n299,
         oc8051_memory_interface1_n298, oc8051_memory_interface1_n297,
         oc8051_memory_interface1_n296, oc8051_memory_interface1_n295,
         oc8051_memory_interface1_n294, oc8051_memory_interface1_n293,
         oc8051_memory_interface1_n292, oc8051_memory_interface1_n291,
         oc8051_memory_interface1_n290, oc8051_memory_interface1_n289,
         oc8051_memory_interface1_n288, oc8051_memory_interface1_n287,
         oc8051_memory_interface1_n286, oc8051_memory_interface1_n285,
         oc8051_memory_interface1_n284, oc8051_memory_interface1_n283,
         oc8051_memory_interface1_n282, oc8051_memory_interface1_n281,
         oc8051_memory_interface1_n280, oc8051_memory_interface1_n279,
         oc8051_memory_interface1_n278, oc8051_memory_interface1_n277,
         oc8051_memory_interface1_n276, oc8051_memory_interface1_n275,
         oc8051_memory_interface1_n274, oc8051_memory_interface1_n273,
         oc8051_memory_interface1_n272, oc8051_memory_interface1_n271,
         oc8051_memory_interface1_n270, oc8051_memory_interface1_n269,
         oc8051_memory_interface1_n268, oc8051_memory_interface1_n267,
         oc8051_memory_interface1_n266, oc8051_memory_interface1_n265,
         oc8051_memory_interface1_n264, oc8051_memory_interface1_n263,
         oc8051_memory_interface1_n262, oc8051_memory_interface1_n261,
         oc8051_memory_interface1_n260, oc8051_memory_interface1_n259,
         oc8051_memory_interface1_n258, oc8051_memory_interface1_n257,
         oc8051_memory_interface1_n256, oc8051_memory_interface1_n255,
         oc8051_memory_interface1_n254, oc8051_memory_interface1_n253,
         oc8051_memory_interface1_n252, oc8051_memory_interface1_n251,
         oc8051_memory_interface1_n250, oc8051_memory_interface1_n249,
         oc8051_memory_interface1_n248, oc8051_memory_interface1_n247,
         oc8051_memory_interface1_n246, oc8051_memory_interface1_n245,
         oc8051_memory_interface1_n244, oc8051_memory_interface1_n243,
         oc8051_memory_interface1_n242, oc8051_memory_interface1_n241,
         oc8051_memory_interface1_n240, oc8051_memory_interface1_n239,
         oc8051_memory_interface1_n238, oc8051_memory_interface1_n237,
         oc8051_memory_interface1_n236, oc8051_memory_interface1_n235,
         oc8051_memory_interface1_n234, oc8051_memory_interface1_n233,
         oc8051_memory_interface1_n232, oc8051_memory_interface1_n231,
         oc8051_memory_interface1_n230, oc8051_memory_interface1_n229,
         oc8051_memory_interface1_n228, oc8051_memory_interface1_n227,
         oc8051_memory_interface1_n226, oc8051_memory_interface1_n225,
         oc8051_memory_interface1_n224, oc8051_memory_interface1_n223,
         oc8051_memory_interface1_n222, oc8051_memory_interface1_n221,
         oc8051_memory_interface1_n220, oc8051_memory_interface1_n219,
         oc8051_memory_interface1_n218, oc8051_memory_interface1_n217,
         oc8051_memory_interface1_n216, oc8051_memory_interface1_n215,
         oc8051_memory_interface1_n214, oc8051_memory_interface1_n213,
         oc8051_memory_interface1_n212, oc8051_memory_interface1_n211,
         oc8051_memory_interface1_n210, oc8051_memory_interface1_n209,
         oc8051_memory_interface1_n208, oc8051_memory_interface1_n207,
         oc8051_memory_interface1_n206, oc8051_memory_interface1_n205,
         oc8051_memory_interface1_n204, oc8051_memory_interface1_n203,
         oc8051_memory_interface1_n202, oc8051_memory_interface1_n201,
         oc8051_memory_interface1_n200, oc8051_memory_interface1_n199,
         oc8051_memory_interface1_n198, oc8051_memory_interface1_n197,
         oc8051_memory_interface1_n196, oc8051_memory_interface1_n195,
         oc8051_memory_interface1_n194, oc8051_memory_interface1_n193,
         oc8051_memory_interface1_n192, oc8051_memory_interface1_n191,
         oc8051_memory_interface1_n190, oc8051_memory_interface1_n189,
         oc8051_memory_interface1_n188, oc8051_memory_interface1_n187,
         oc8051_memory_interface1_n186, oc8051_memory_interface1_n185,
         oc8051_memory_interface1_n184, oc8051_memory_interface1_n183,
         oc8051_memory_interface1_n182, oc8051_memory_interface1_n181,
         oc8051_memory_interface1_n180, oc8051_memory_interface1_n179,
         oc8051_memory_interface1_n178, oc8051_memory_interface1_n177,
         oc8051_memory_interface1_n176, oc8051_memory_interface1_n175,
         oc8051_memory_interface1_n174, oc8051_memory_interface1_n173,
         oc8051_memory_interface1_n172, oc8051_memory_interface1_n171,
         oc8051_memory_interface1_n170, oc8051_memory_interface1_n169,
         oc8051_memory_interface1_n168, oc8051_memory_interface1_n167,
         oc8051_memory_interface1_n166, oc8051_memory_interface1_n165,
         oc8051_memory_interface1_n164, oc8051_memory_interface1_n163,
         oc8051_memory_interface1_n162, oc8051_memory_interface1_n161,
         oc8051_memory_interface1_n160, oc8051_memory_interface1_n159,
         oc8051_memory_interface1_n158, oc8051_memory_interface1_n157,
         oc8051_memory_interface1_n156, oc8051_memory_interface1_n155,
         oc8051_memory_interface1_n154, oc8051_memory_interface1_n153,
         oc8051_memory_interface1_n152, oc8051_memory_interface1_n151,
         oc8051_memory_interface1_n150, oc8051_memory_interface1_n149,
         oc8051_memory_interface1_n148, oc8051_memory_interface1_n147,
         oc8051_memory_interface1_n146, oc8051_memory_interface1_n145,
         oc8051_memory_interface1_n144, oc8051_memory_interface1_n143,
         oc8051_memory_interface1_n142, oc8051_memory_interface1_n141,
         oc8051_memory_interface1_n140, oc8051_memory_interface1_n139,
         oc8051_memory_interface1_n138, oc8051_memory_interface1_n137,
         oc8051_memory_interface1_n136, oc8051_memory_interface1_n135,
         oc8051_memory_interface1_n134, oc8051_memory_interface1_n133,
         oc8051_memory_interface1_n132, oc8051_memory_interface1_n131,
         oc8051_memory_interface1_n130, oc8051_memory_interface1_n129,
         oc8051_memory_interface1_n128, oc8051_memory_interface1_n127,
         oc8051_memory_interface1_n126, oc8051_memory_interface1_n125,
         oc8051_memory_interface1_n124, oc8051_memory_interface1_n123,
         oc8051_memory_interface1_n122, oc8051_memory_interface1_n121,
         oc8051_memory_interface1_n120, oc8051_memory_interface1_n119,
         oc8051_memory_interface1_n118, oc8051_memory_interface1_n117,
         oc8051_memory_interface1_n116, oc8051_memory_interface1_n115,
         oc8051_memory_interface1_n114, oc8051_memory_interface1_n113,
         oc8051_memory_interface1_n112, oc8051_memory_interface1_n111,
         oc8051_memory_interface1_n110, oc8051_memory_interface1_n109,
         oc8051_memory_interface1_n108, oc8051_memory_interface1_n107,
         oc8051_memory_interface1_n106, oc8051_memory_interface1_n105,
         oc8051_memory_interface1_n104, oc8051_memory_interface1_n103,
         oc8051_memory_interface1_n102, oc8051_memory_interface1_n101,
         oc8051_memory_interface1_n100, oc8051_memory_interface1_n99,
         oc8051_memory_interface1_n98, oc8051_memory_interface1_n97,
         oc8051_memory_interface1_n96, oc8051_memory_interface1_n95,
         oc8051_memory_interface1_n94, oc8051_memory_interface1_n93,
         oc8051_memory_interface1_n92, oc8051_memory_interface1_n91,
         oc8051_memory_interface1_n90, oc8051_memory_interface1_n89,
         oc8051_memory_interface1_n88, oc8051_memory_interface1_n87,
         oc8051_memory_interface1_n86, oc8051_memory_interface1_n85,
         oc8051_memory_interface1_n84, oc8051_memory_interface1_n83,
         oc8051_memory_interface1_n82, oc8051_memory_interface1_n81,
         oc8051_memory_interface1_n80, oc8051_memory_interface1_n79,
         oc8051_memory_interface1_n78, oc8051_memory_interface1_n77,
         oc8051_memory_interface1_n76, oc8051_memory_interface1_n75,
         oc8051_memory_interface1_n74, oc8051_memory_interface1_n73,
         oc8051_memory_interface1_n72, oc8051_memory_interface1_n71,
         oc8051_memory_interface1_n70, oc8051_memory_interface1_n69,
         oc8051_memory_interface1_n68, oc8051_memory_interface1_n67,
         oc8051_memory_interface1_n66, oc8051_memory_interface1_n65,
         oc8051_memory_interface1_n64, oc8051_memory_interface1_n63,
         oc8051_memory_interface1_n62, oc8051_memory_interface1_n61,
         oc8051_memory_interface1_n60, oc8051_memory_interface1_n59,
         oc8051_memory_interface1_n58, oc8051_memory_interface1_n57,
         oc8051_memory_interface1_n56, oc8051_memory_interface1_n55,
         oc8051_memory_interface1_n54, oc8051_memory_interface1_n53,
         oc8051_memory_interface1_n52, oc8051_memory_interface1_n51,
         oc8051_memory_interface1_n50, oc8051_memory_interface1_n49,
         oc8051_memory_interface1_n48, oc8051_memory_interface1_n47,
         oc8051_memory_interface1_n46, oc8051_memory_interface1_n45,
         oc8051_memory_interface1_n44, oc8051_memory_interface1_n43,
         oc8051_memory_interface1_n42, oc8051_memory_interface1_n41,
         oc8051_memory_interface1_n40, oc8051_memory_interface1_n39,
         oc8051_memory_interface1_n38, oc8051_memory_interface1_n37,
         oc8051_memory_interface1_n36, oc8051_memory_interface1_n35,
         oc8051_memory_interface1_n34, oc8051_memory_interface1_n33,
         oc8051_memory_interface1_n32, oc8051_memory_interface1_n31,
         oc8051_memory_interface1_n30, oc8051_memory_interface1_n29,
         oc8051_memory_interface1_n28, oc8051_memory_interface1_n27,
         oc8051_memory_interface1_n26, oc8051_memory_interface1_n25,
         oc8051_memory_interface1_n24, oc8051_memory_interface1_n23,
         oc8051_memory_interface1_n22, oc8051_memory_interface1_n21,
         oc8051_memory_interface1_n20, oc8051_memory_interface1_n19,
         oc8051_memory_interface1_n18, oc8051_memory_interface1_n17,
         oc8051_memory_interface1_n16, oc8051_memory_interface1_n15,
         oc8051_memory_interface1_n14, oc8051_memory_interface1_n13,
         oc8051_memory_interface1_n12, oc8051_memory_interface1_n11,
         oc8051_memory_interface1_n10, oc8051_memory_interface1_n9,
         oc8051_memory_interface1_n8, oc8051_memory_interface1_n7,
         oc8051_memory_interface1_n6, oc8051_memory_interface1_n5,
         oc8051_memory_interface1_n4, oc8051_memory_interface1_n3,
         oc8051_memory_interface1_n2, oc8051_memory_interface1_n1,
         oc8051_memory_interface1_n584, oc8051_memory_interface1_n583,
         oc8051_memory_interface1_n582, oc8051_memory_interface1_n581,
         oc8051_memory_interface1_n580, oc8051_memory_interface1_n579,
         oc8051_memory_interface1_n578, oc8051_memory_interface1_n577,
         oc8051_memory_interface1_n576, oc8051_memory_interface1_n575,
         oc8051_memory_interface1_n574, oc8051_memory_interface1_n573,
         oc8051_memory_interface1_n572, oc8051_memory_interface1_n571,
         oc8051_memory_interface1_n570, oc8051_memory_interface1_n569,
         oc8051_memory_interface1_n568, oc8051_memory_interface1_n567,
         oc8051_memory_interface1_n566, oc8051_memory_interface1_n565,
         oc8051_memory_interface1_n564, oc8051_memory_interface1_n563,
         oc8051_memory_interface1_n562, oc8051_memory_interface1_n561,
         oc8051_memory_interface1_n560, oc8051_memory_interface1_n559,
         oc8051_memory_interface1_n558, oc8051_memory_interface1_n557,
         oc8051_memory_interface1_n555, oc8051_memory_interface1_n553,
         oc8051_memory_interface1_n551, oc8051_memory_interface1_n549,
         oc8051_memory_interface1_n547, oc8051_memory_interface1_n545,
         oc8051_memory_interface1_n543, oc8051_memory_interface1_n541,
         oc8051_memory_interface1_n540, oc8051_memory_interface1_n539,
         oc8051_memory_interface1_n538, oc8051_memory_interface1_n537,
         oc8051_memory_interface1_n536, oc8051_memory_interface1_n535,
         oc8051_memory_interface1_n534, oc8051_memory_interface1_n533,
         oc8051_memory_interface1_n532, oc8051_memory_interface1_n531,
         oc8051_memory_interface1_n530, oc8051_memory_interface1_n529,
         oc8051_memory_interface1_n528, oc8051_memory_interface1_n527,
         oc8051_memory_interface1_n526, oc8051_memory_interface1_n525,
         oc8051_memory_interface1_n524, oc8051_memory_interface1_n523,
         oc8051_memory_interface1_n522, oc8051_memory_interface1_n521,
         oc8051_memory_interface1_n520, oc8051_memory_interface1_n519,
         oc8051_memory_interface1_n518, oc8051_memory_interface1_n517,
         oc8051_memory_interface1_n516, oc8051_memory_interface1_n515,
         oc8051_memory_interface1_n514, oc8051_memory_interface1_n513,
         oc8051_memory_interface1_n512, oc8051_memory_interface1_n511,
         oc8051_memory_interface1_n510, oc8051_memory_interface1_n509,
         oc8051_memory_interface1_n508, oc8051_memory_interface1_n507,
         oc8051_memory_interface1_n506, oc8051_memory_interface1_n505,
         oc8051_memory_interface1_n504, oc8051_memory_interface1_n503,
         oc8051_memory_interface1_n502, oc8051_memory_interface1_n501,
         oc8051_memory_interface1_n500, oc8051_memory_interface1_n499,
         oc8051_memory_interface1_n498, oc8051_memory_interface1_n497,
         oc8051_memory_interface1_n496, oc8051_memory_interface1_n495,
         oc8051_memory_interface1_n494, oc8051_memory_interface1_n493,
         oc8051_memory_interface1_n492, oc8051_memory_interface1_n491,
         oc8051_memory_interface1_n490, oc8051_memory_interface1_n489,
         oc8051_memory_interface1_n488, oc8051_memory_interface1_n487,
         oc8051_memory_interface1_n486, oc8051_memory_interface1_n485,
         oc8051_memory_interface1_n484, oc8051_memory_interface1_n483,
         oc8051_memory_interface1_n482, oc8051_memory_interface1_n481,
         oc8051_memory_interface1_n480, oc8051_memory_interface1_n479,
         oc8051_memory_interface1_n478, oc8051_memory_interface1_n477,
         oc8051_memory_interface1_n476, oc8051_memory_interface1_n475,
         oc8051_memory_interface1_n474, oc8051_memory_interface1_n473,
         oc8051_memory_interface1_n472, oc8051_memory_interface1_n471,
         oc8051_memory_interface1_n470, oc8051_memory_interface1_n469,
         oc8051_memory_interface1_n468, oc8051_memory_interface1_n467,
         oc8051_memory_interface1_n466, oc8051_memory_interface1_n465,
         oc8051_memory_interface1_n464, oc8051_memory_interface1_n463,
         oc8051_memory_interface1_n462, oc8051_memory_interface1_n461,
         oc8051_memory_interface1_n460, oc8051_memory_interface1_n459,
         oc8051_memory_interface1_n455, oc8051_memory_interface1_n454,
         oc8051_memory_interface1_n453, oc8051_memory_interface1_n452,
         oc8051_memory_interface1_n451, oc8051_memory_interface1_n450,
         oc8051_memory_interface1_n449, oc8051_memory_interface1_n448,
         oc8051_memory_interface1_n447, oc8051_memory_interface1_n446,
         oc8051_memory_interface1_n445, oc8051_memory_interface1_n444,
         oc8051_memory_interface1_n443, oc8051_memory_interface1_n442,
         oc8051_memory_interface1_n441, oc8051_memory_interface1_n440,
         oc8051_memory_interface1_n431, oc8051_memory_interface1_n430,
         oc8051_memory_interface1_n429, oc8051_memory_interface1_n428,
         oc8051_memory_interface1_n427, oc8051_memory_interface1_n426,
         oc8051_memory_interface1_n425, oc8051_memory_interface1_n424,
         oc8051_memory_interface1_n423, oc8051_memory_interface1_n422,
         oc8051_memory_interface1_n421, oc8051_memory_interface1_n420,
         oc8051_memory_interface1_n419, oc8051_memory_interface1_n418,
         oc8051_memory_interface1_n417, oc8051_memory_interface1_n416,
         oc8051_memory_interface1_n399, oc8051_memory_interface1_n398,
         oc8051_memory_interface1_n397, oc8051_memory_interface1_n396,
         oc8051_memory_interface1_n395, oc8051_memory_interface1_n394,
         oc8051_memory_interface1_n393, oc8051_memory_interface1_n392,
         oc8051_memory_interface1_n5530, oc8051_memory_interface1_pc_wr_r,
         oc8051_memory_interface1_pc_buf_0_,
         oc8051_memory_interface1_pc_buf_1_,
         oc8051_memory_interface1_pc_buf_2_,
         oc8051_memory_interface1_pc_buf_3_,
         oc8051_memory_interface1_pc_buf_4_,
         oc8051_memory_interface1_pc_buf_5_,
         oc8051_memory_interface1_pc_buf_6_,
         oc8051_memory_interface1_pc_buf_7_,
         oc8051_memory_interface1_pc_buf_8_,
         oc8051_memory_interface1_pc_buf_9_,
         oc8051_memory_interface1_pc_buf_10_,
         oc8051_memory_interface1_pc_buf_11_,
         oc8051_memory_interface1_pc_buf_12_,
         oc8051_memory_interface1_pc_buf_13_,
         oc8051_memory_interface1_pc_buf_14_,
         oc8051_memory_interface1_pc_buf_15_, oc8051_memory_interface1_n3720,
         oc8051_memory_interface1_int_ack_buff, oc8051_memory_interface1_n2000,
         oc8051_memory_interface1_int_vec_buff_0_,
         oc8051_memory_interface1_int_vec_buff_1_,
         oc8051_memory_interface1_int_vec_buff_2_,
         oc8051_memory_interface1_int_vec_buff_3_,
         oc8051_memory_interface1_int_vec_buff_4_,
         oc8051_memory_interface1_int_vec_buff_5_,
         oc8051_memory_interface1_int_vec_buff_6_,
         oc8051_memory_interface1_int_vec_buff_7_,
         oc8051_memory_interface1_int_ack_t,
         oc8051_memory_interface1_ddat_ir_0_,
         oc8051_memory_interface1_ddat_ir_1_,
         oc8051_memory_interface1_ddat_ir_2_,
         oc8051_memory_interface1_ddat_ir_3_,
         oc8051_memory_interface1_ddat_ir_4_,
         oc8051_memory_interface1_ddat_ir_5_,
         oc8051_memory_interface1_ddat_ir_6_,
         oc8051_memory_interface1_ddat_ir_7_, oc8051_memory_interface1_dack_ir,
         oc8051_memory_interface1_op1_0_, oc8051_memory_interface1_op1_1_,
         oc8051_memory_interface1_op1_2_, oc8051_memory_interface1_op1_3_,
         oc8051_memory_interface1_op1_4_, oc8051_memory_interface1_op1_5_,
         oc8051_memory_interface1_op1_6_, oc8051_memory_interface1_op1_7_,
         oc8051_memory_interface1_op_pos_0_,
         oc8051_memory_interface1_op_pos_1_,
         oc8051_memory_interface1_op_pos_2_, oc8051_memory_interface1_cdone,
         oc8051_memory_interface1_cdata_0_, oc8051_memory_interface1_cdata_1_,
         oc8051_memory_interface1_cdata_2_, oc8051_memory_interface1_cdata_3_,
         oc8051_memory_interface1_cdata_4_, oc8051_memory_interface1_cdata_5_,
         oc8051_memory_interface1_cdata_6_, oc8051_memory_interface1_cdata_7_,
         oc8051_memory_interface1_idat_cur_0_,
         oc8051_memory_interface1_idat_cur_1_,
         oc8051_memory_interface1_idat_cur_2_,
         oc8051_memory_interface1_idat_cur_3_,
         oc8051_memory_interface1_idat_cur_4_,
         oc8051_memory_interface1_idat_cur_5_,
         oc8051_memory_interface1_idat_cur_6_,
         oc8051_memory_interface1_idat_cur_7_,
         oc8051_memory_interface1_idat_cur_8_,
         oc8051_memory_interface1_idat_cur_9_,
         oc8051_memory_interface1_idat_cur_10_,
         oc8051_memory_interface1_idat_cur_11_,
         oc8051_memory_interface1_idat_cur_12_,
         oc8051_memory_interface1_idat_cur_13_,
         oc8051_memory_interface1_idat_cur_14_,
         oc8051_memory_interface1_idat_cur_15_,
         oc8051_memory_interface1_idat_cur_16_,
         oc8051_memory_interface1_idat_cur_17_,
         oc8051_memory_interface1_idat_cur_18_,
         oc8051_memory_interface1_idat_cur_19_,
         oc8051_memory_interface1_idat_cur_20_,
         oc8051_memory_interface1_idat_cur_21_,
         oc8051_memory_interface1_idat_cur_22_,
         oc8051_memory_interface1_idat_cur_23_,
         oc8051_memory_interface1_idat_cur_24_,
         oc8051_memory_interface1_idat_cur_25_,
         oc8051_memory_interface1_idat_cur_26_,
         oc8051_memory_interface1_idat_cur_27_,
         oc8051_memory_interface1_idat_cur_28_,
         oc8051_memory_interface1_idat_cur_29_,
         oc8051_memory_interface1_idat_cur_30_,
         oc8051_memory_interface1_idat_cur_31_,
         oc8051_memory_interface1_idat_old_0_,
         oc8051_memory_interface1_idat_old_1_,
         oc8051_memory_interface1_idat_old_2_,
         oc8051_memory_interface1_idat_old_3_,
         oc8051_memory_interface1_idat_old_4_,
         oc8051_memory_interface1_idat_old_5_,
         oc8051_memory_interface1_idat_old_6_,
         oc8051_memory_interface1_idat_old_7_,
         oc8051_memory_interface1_idat_old_8_,
         oc8051_memory_interface1_idat_old_9_,
         oc8051_memory_interface1_idat_old_10_,
         oc8051_memory_interface1_idat_old_11_,
         oc8051_memory_interface1_idat_old_12_,
         oc8051_memory_interface1_idat_old_13_,
         oc8051_memory_interface1_idat_old_14_,
         oc8051_memory_interface1_idat_old_15_,
         oc8051_memory_interface1_idat_old_16_,
         oc8051_memory_interface1_idat_old_17_,
         oc8051_memory_interface1_idat_old_18_,
         oc8051_memory_interface1_idat_old_19_,
         oc8051_memory_interface1_idat_old_20_,
         oc8051_memory_interface1_idat_old_21_,
         oc8051_memory_interface1_idat_old_22_,
         oc8051_memory_interface1_idat_old_23_,
         oc8051_memory_interface1_idat_old_24_,
         oc8051_memory_interface1_idat_old_25_,
         oc8051_memory_interface1_idat_old_26_,
         oc8051_memory_interface1_idat_old_27_,
         oc8051_memory_interface1_idat_old_28_,
         oc8051_memory_interface1_idat_old_29_,
         oc8051_memory_interface1_idat_old_30_,
         oc8051_memory_interface1_idat_old_31_, oc8051_memory_interface1_n1310,
         oc8051_memory_interface1_iadr_t_0_,
         oc8051_memory_interface1_iadr_t_1_,
         oc8051_memory_interface1_iadr_t_2_,
         oc8051_memory_interface1_iadr_t_3_,
         oc8051_memory_interface1_iadr_t_4_,
         oc8051_memory_interface1_iadr_t_5_,
         oc8051_memory_interface1_iadr_t_6_,
         oc8051_memory_interface1_iadr_t_7_,
         oc8051_memory_interface1_iadr_t_8_,
         oc8051_memory_interface1_iadr_t_9_,
         oc8051_memory_interface1_iadr_t_10_,
         oc8051_memory_interface1_iadr_t_11_,
         oc8051_memory_interface1_iadr_t_12_,
         oc8051_memory_interface1_iadr_t_13_,
         oc8051_memory_interface1_iadr_t_14_,
         oc8051_memory_interface1_iadr_t_15_, oc8051_memory_interface1_n830,
         oc8051_memory_interface1_rd_addr_r, oc8051_memory_interface1_istb_t,
         oc8051_memory_interface1_pc_wr_r2, oc8051_memory_interface1_imem_wait,
         oc8051_memory_interface1_dmem_wait, oc8051_memory_interface1_istb_o,
         oc8051_memory_interface1_rd_ind, oc8051_sfr1_n259, oc8051_sfr1_n258,
         oc8051_sfr1_n257, oc8051_sfr1_n256, oc8051_sfr1_n255,
         oc8051_sfr1_n254, oc8051_sfr1_n253, oc8051_sfr1_n252,
         oc8051_sfr1_n251, oc8051_sfr1_n250, oc8051_sfr1_n249,
         oc8051_sfr1_n248, oc8051_sfr1_n247, oc8051_sfr1_n246,
         oc8051_sfr1_n245, oc8051_sfr1_n236, oc8051_sfr1_n235,
         oc8051_sfr1_n234, oc8051_sfr1_n233, oc8051_sfr1_n232,
         oc8051_sfr1_n231, oc8051_sfr1_n230, oc8051_sfr1_n229,
         oc8051_sfr1_n228, oc8051_sfr1_n227, oc8051_sfr1_n226,
         oc8051_sfr1_n225, oc8051_sfr1_n224, oc8051_sfr1_n223,
         oc8051_sfr1_n222, oc8051_sfr1_n221, oc8051_sfr1_n220,
         oc8051_sfr1_n219, oc8051_sfr1_n218, oc8051_sfr1_n217,
         oc8051_sfr1_n216, oc8051_sfr1_n215, oc8051_sfr1_n214,
         oc8051_sfr1_n213, oc8051_sfr1_n212, oc8051_sfr1_n211,
         oc8051_sfr1_n210, oc8051_sfr1_n209, oc8051_sfr1_n208,
         oc8051_sfr1_n207, oc8051_sfr1_n206, oc8051_sfr1_n205,
         oc8051_sfr1_n204, oc8051_sfr1_n203, oc8051_sfr1_n202,
         oc8051_sfr1_n201, oc8051_sfr1_n200, oc8051_sfr1_n199,
         oc8051_sfr1_n198, oc8051_sfr1_n197, oc8051_sfr1_n196,
         oc8051_sfr1_n195, oc8051_sfr1_n194, oc8051_sfr1_n193,
         oc8051_sfr1_n192, oc8051_sfr1_n191, oc8051_sfr1_n190,
         oc8051_sfr1_n189, oc8051_sfr1_n188, oc8051_sfr1_n187,
         oc8051_sfr1_n186, oc8051_sfr1_n185, oc8051_sfr1_n184,
         oc8051_sfr1_n183, oc8051_sfr1_n182, oc8051_sfr1_n181,
         oc8051_sfr1_n180, oc8051_sfr1_n179, oc8051_sfr1_n178,
         oc8051_sfr1_n177, oc8051_sfr1_n176, oc8051_sfr1_n175,
         oc8051_sfr1_n174, oc8051_sfr1_n173, oc8051_sfr1_n172,
         oc8051_sfr1_n171, oc8051_sfr1_n170, oc8051_sfr1_n169,
         oc8051_sfr1_n168, oc8051_sfr1_n167, oc8051_sfr1_n166,
         oc8051_sfr1_n165, oc8051_sfr1_n164, oc8051_sfr1_n163,
         oc8051_sfr1_n162, oc8051_sfr1_n161, oc8051_sfr1_n160,
         oc8051_sfr1_n159, oc8051_sfr1_n158, oc8051_sfr1_n157,
         oc8051_sfr1_n156, oc8051_sfr1_n155, oc8051_sfr1_n154,
         oc8051_sfr1_n153, oc8051_sfr1_n152, oc8051_sfr1_n151,
         oc8051_sfr1_n150, oc8051_sfr1_n149, oc8051_sfr1_n148,
         oc8051_sfr1_n147, oc8051_sfr1_n146, oc8051_sfr1_n145,
         oc8051_sfr1_n144, oc8051_sfr1_n143, oc8051_sfr1_n142,
         oc8051_sfr1_n141, oc8051_sfr1_n140, oc8051_sfr1_n139,
         oc8051_sfr1_n138, oc8051_sfr1_n137, oc8051_sfr1_n136,
         oc8051_sfr1_n135, oc8051_sfr1_n134, oc8051_sfr1_n133,
         oc8051_sfr1_n132, oc8051_sfr1_n131, oc8051_sfr1_n130,
         oc8051_sfr1_n129, oc8051_sfr1_n128, oc8051_sfr1_n127,
         oc8051_sfr1_n126, oc8051_sfr1_n125, oc8051_sfr1_n124,
         oc8051_sfr1_n123, oc8051_sfr1_n122, oc8051_sfr1_n121,
         oc8051_sfr1_n120, oc8051_sfr1_n119, oc8051_sfr1_n118,
         oc8051_sfr1_n117, oc8051_sfr1_n116, oc8051_sfr1_n115,
         oc8051_sfr1_n114, oc8051_sfr1_n113, oc8051_sfr1_n112,
         oc8051_sfr1_n111, oc8051_sfr1_n110, oc8051_sfr1_n109,
         oc8051_sfr1_n108, oc8051_sfr1_n107, oc8051_sfr1_n106,
         oc8051_sfr1_n105, oc8051_sfr1_n104, oc8051_sfr1_n103,
         oc8051_sfr1_n102, oc8051_sfr1_n101, oc8051_sfr1_n100, oc8051_sfr1_n99,
         oc8051_sfr1_n98, oc8051_sfr1_n97, oc8051_sfr1_n96, oc8051_sfr1_n95,
         oc8051_sfr1_n94, oc8051_sfr1_n93, oc8051_sfr1_n92, oc8051_sfr1_n91,
         oc8051_sfr1_n90, oc8051_sfr1_n89, oc8051_sfr1_n88, oc8051_sfr1_n87,
         oc8051_sfr1_n86, oc8051_sfr1_n85, oc8051_sfr1_n84, oc8051_sfr1_n83,
         oc8051_sfr1_n82, oc8051_sfr1_n81, oc8051_sfr1_n80, oc8051_sfr1_n79,
         oc8051_sfr1_n78, oc8051_sfr1_n77, oc8051_sfr1_n76, oc8051_sfr1_n75,
         oc8051_sfr1_n74, oc8051_sfr1_n73, oc8051_sfr1_n72, oc8051_sfr1_n71,
         oc8051_sfr1_n70, oc8051_sfr1_n69, oc8051_sfr1_n68, oc8051_sfr1_n67,
         oc8051_sfr1_n66, oc8051_sfr1_n65, oc8051_sfr1_n64, oc8051_sfr1_n63,
         oc8051_sfr1_n62, oc8051_sfr1_n61, oc8051_sfr1_n60, oc8051_sfr1_n59,
         oc8051_sfr1_n58, oc8051_sfr1_n57, oc8051_sfr1_n56, oc8051_sfr1_n55,
         oc8051_sfr1_n54, oc8051_sfr1_n53, oc8051_sfr1_n52, oc8051_sfr1_n51,
         oc8051_sfr1_n50, oc8051_sfr1_n49, oc8051_sfr1_n48, oc8051_sfr1_n47,
         oc8051_sfr1_n46, oc8051_sfr1_n45, oc8051_sfr1_n44, oc8051_sfr1_n43,
         oc8051_sfr1_n42, oc8051_sfr1_n41, oc8051_sfr1_n40, oc8051_sfr1_n39,
         oc8051_sfr1_n38, oc8051_sfr1_n37, oc8051_sfr1_n36, oc8051_sfr1_n35,
         oc8051_sfr1_n34, oc8051_sfr1_n33, oc8051_sfr1_n32, oc8051_sfr1_n31,
         oc8051_sfr1_n30, oc8051_sfr1_n29, oc8051_sfr1_n28, oc8051_sfr1_n27,
         oc8051_sfr1_n26, oc8051_sfr1_n25, oc8051_sfr1_n24, oc8051_sfr1_n23,
         oc8051_sfr1_n22, oc8051_sfr1_n21, oc8051_sfr1_n20, oc8051_sfr1_n19,
         oc8051_sfr1_n18, oc8051_sfr1_n17, oc8051_sfr1_n16, oc8051_sfr1_n15,
         oc8051_sfr1_n14, oc8051_sfr1_n13, oc8051_sfr1_n12, oc8051_sfr1_n11,
         oc8051_sfr1_n10, oc8051_sfr1_n9, oc8051_sfr1_n8, oc8051_sfr1_n7,
         oc8051_sfr1_n6, oc8051_sfr1_n5, oc8051_sfr1_n4, oc8051_sfr1_n3,
         oc8051_sfr1_n2, oc8051_sfr1_int_src_2_, oc8051_sfr1_n244,
         oc8051_sfr1_n243, oc8051_sfr1_n242, oc8051_sfr1_n241,
         oc8051_sfr1_n240, oc8051_sfr1_n239, oc8051_sfr1_n238,
         oc8051_sfr1_n237, oc8051_sfr1_n1520, oc8051_sfr1_n1510,
         oc8051_sfr1_n1500, oc8051_sfr1_prescaler_0_, oc8051_sfr1_prescaler_1_,
         oc8051_sfr1_prescaler_2_, oc8051_sfr1_prescaler_3_, oc8051_sfr1_n1400,
         oc8051_sfr1_n1380, oc8051_sfr1_n1370, oc8051_sfr1_n1360,
         oc8051_sfr1_n1350, oc8051_sfr1_n1340, oc8051_sfr1_n1330,
         oc8051_sfr1_n1320, oc8051_sfr1_n1310, oc8051_sfr1_n1300,
         oc8051_sfr1_n1290, oc8051_sfr1_n1280, oc8051_sfr1_n1270,
         oc8051_sfr1_n1020, oc8051_sfr1_t2con_0_, oc8051_sfr1_t2con_1_,
         oc8051_sfr1_t2con_2_, oc8051_sfr1_t2con_3_, oc8051_sfr1_t2con_6_,
         oc8051_sfr1_t2con_7_, oc8051_sfr1_ip_0_, oc8051_sfr1_ip_1_,
         oc8051_sfr1_ip_2_, oc8051_sfr1_ip_3_, oc8051_sfr1_ip_4_,
         oc8051_sfr1_ip_5_, oc8051_sfr1_ip_6_, oc8051_sfr1_ip_7_,
         oc8051_sfr1_tcon_0_, oc8051_sfr1_tcon_1_, oc8051_sfr1_tcon_2_,
         oc8051_sfr1_tcon_3_, oc8051_sfr1_tcon_5_, oc8051_sfr1_tcon_7_,
         oc8051_sfr1_ie_0_, oc8051_sfr1_ie_1_, oc8051_sfr1_ie_2_,
         oc8051_sfr1_ie_3_, oc8051_sfr1_ie_4_, oc8051_sfr1_ie_5_,
         oc8051_sfr1_ie_6_, oc8051_sfr1_ie_7_, oc8051_sfr1_tr1,
         oc8051_sfr1_tr0, oc8051_sfr1_tc2_int, oc8051_sfr1_tf0,
         oc8051_sfr1_scon_0_, oc8051_sfr1_scon_1_, oc8051_sfr1_scon_2_,
         oc8051_sfr1_scon_3_, oc8051_sfr1_scon_4_, oc8051_sfr1_scon_5_,
         oc8051_sfr1_scon_6_, oc8051_sfr1_scon_7_, oc8051_sfr1_tclk,
         oc8051_sfr1_rclk, oc8051_sfr1_pres_ow, oc8051_sfr1_tf1,
         oc8051_sfr1_brate2, oc8051_sfr1_uart_int, oc8051_sfr1_p3_data_0_,
         oc8051_sfr1_p3_data_1_, oc8051_sfr1_p3_data_2_,
         oc8051_sfr1_p3_data_3_, oc8051_sfr1_p3_data_4_,
         oc8051_sfr1_p3_data_5_, oc8051_sfr1_p3_data_6_,
         oc8051_sfr1_p3_data_7_, oc8051_sfr1_p2_data_0_,
         oc8051_sfr1_p2_data_1_, oc8051_sfr1_p2_data_2_,
         oc8051_sfr1_p2_data_3_, oc8051_sfr1_p2_data_4_,
         oc8051_sfr1_p2_data_5_, oc8051_sfr1_p2_data_6_,
         oc8051_sfr1_p2_data_7_, oc8051_sfr1_p1_data_0_,
         oc8051_sfr1_p1_data_1_, oc8051_sfr1_p1_data_2_,
         oc8051_sfr1_p1_data_3_, oc8051_sfr1_p1_data_4_,
         oc8051_sfr1_p1_data_5_, oc8051_sfr1_p1_data_6_,
         oc8051_sfr1_p1_data_7_, oc8051_sfr1_p0_data_0_,
         oc8051_sfr1_p0_data_1_, oc8051_sfr1_p0_data_2_,
         oc8051_sfr1_p0_data_3_, oc8051_sfr1_p0_data_4_,
         oc8051_sfr1_p0_data_5_, oc8051_sfr1_p0_data_6_,
         oc8051_sfr1_p0_data_7_, oc8051_sfr1_b_reg_0_, oc8051_sfr1_b_reg_1_,
         oc8051_sfr1_b_reg_2_, oc8051_sfr1_b_reg_3_, oc8051_sfr1_b_reg_4_,
         oc8051_sfr1_b_reg_5_, oc8051_sfr1_b_reg_6_, oc8051_sfr1_b_reg_7_,
         oc8051_sfr1_wr_bit_r, oc8051_sfr1_psw_0_, oc8051_sfr1_psw_1_,
         oc8051_sfr1_psw_2_, oc8051_sfr1_psw_3_, oc8051_sfr1_psw_4_,
         oc8051_sfr1_psw_5_, oc8051_sfr1_oc8051_acc1_n66,
         oc8051_sfr1_oc8051_acc1_n65, oc8051_sfr1_oc8051_acc1_n64,
         oc8051_sfr1_oc8051_acc1_n63, oc8051_sfr1_oc8051_acc1_n62,
         oc8051_sfr1_oc8051_acc1_n61, oc8051_sfr1_oc8051_acc1_n60,
         oc8051_sfr1_oc8051_acc1_n59, oc8051_sfr1_oc8051_acc1_n58,
         oc8051_sfr1_oc8051_acc1_n57, oc8051_sfr1_oc8051_acc1_n56,
         oc8051_sfr1_oc8051_acc1_n55, oc8051_sfr1_oc8051_acc1_n54,
         oc8051_sfr1_oc8051_acc1_n53, oc8051_sfr1_oc8051_acc1_n52,
         oc8051_sfr1_oc8051_acc1_n51, oc8051_sfr1_oc8051_acc1_n50,
         oc8051_sfr1_oc8051_acc1_n49, oc8051_sfr1_oc8051_acc1_n48,
         oc8051_sfr1_oc8051_acc1_n47, oc8051_sfr1_oc8051_acc1_n46,
         oc8051_sfr1_oc8051_acc1_n45, oc8051_sfr1_oc8051_acc1_n44,
         oc8051_sfr1_oc8051_acc1_n43, oc8051_sfr1_oc8051_acc1_n42,
         oc8051_sfr1_oc8051_acc1_n41, oc8051_sfr1_oc8051_acc1_n40,
         oc8051_sfr1_oc8051_acc1_n39, oc8051_sfr1_oc8051_acc1_n38,
         oc8051_sfr1_oc8051_acc1_n37, oc8051_sfr1_oc8051_acc1_n36,
         oc8051_sfr1_oc8051_acc1_n35, oc8051_sfr1_oc8051_acc1_n34,
         oc8051_sfr1_oc8051_acc1_n33, oc8051_sfr1_oc8051_acc1_n32,
         oc8051_sfr1_oc8051_acc1_n31, oc8051_sfr1_oc8051_acc1_n30,
         oc8051_sfr1_oc8051_acc1_n29, oc8051_sfr1_oc8051_acc1_n28,
         oc8051_sfr1_oc8051_acc1_n27, oc8051_sfr1_oc8051_acc1_n26,
         oc8051_sfr1_oc8051_acc1_n25, oc8051_sfr1_oc8051_acc1_n24,
         oc8051_sfr1_oc8051_acc1_n23, oc8051_sfr1_oc8051_acc1_n22,
         oc8051_sfr1_oc8051_acc1_n21, oc8051_sfr1_oc8051_acc1_n20,
         oc8051_sfr1_oc8051_acc1_n19, oc8051_sfr1_oc8051_acc1_n18,
         oc8051_sfr1_oc8051_acc1_n17, oc8051_sfr1_oc8051_acc1_n16,
         oc8051_sfr1_oc8051_acc1_n15, oc8051_sfr1_oc8051_acc1_n14,
         oc8051_sfr1_oc8051_acc1_n13, oc8051_sfr1_oc8051_acc1_n12,
         oc8051_sfr1_oc8051_acc1_n11, oc8051_sfr1_oc8051_acc1_n10,
         oc8051_sfr1_oc8051_acc1_n9, oc8051_sfr1_oc8051_acc1_n8,
         oc8051_sfr1_oc8051_acc1_n7, oc8051_sfr1_oc8051_acc1_n6,
         oc8051_sfr1_oc8051_acc1_n5, oc8051_sfr1_oc8051_acc1_n4,
         oc8051_sfr1_oc8051_acc1_n3, oc8051_sfr1_oc8051_acc1_n2,
         oc8051_sfr1_oc8051_acc1_n1, oc8051_sfr1_oc8051_acc1_acc_0_,
         oc8051_sfr1_oc8051_acc1_acc_1_, oc8051_sfr1_oc8051_acc1_acc_2_,
         oc8051_sfr1_oc8051_acc1_acc_3_, oc8051_sfr1_oc8051_acc1_acc_4_,
         oc8051_sfr1_oc8051_acc1_acc_5_, oc8051_sfr1_oc8051_acc1_acc_6_,
         oc8051_sfr1_oc8051_acc1_acc_7_, oc8051_sfr1_oc8051_b_register_n28,
         oc8051_sfr1_oc8051_b_register_n27, oc8051_sfr1_oc8051_b_register_n26,
         oc8051_sfr1_oc8051_b_register_n25, oc8051_sfr1_oc8051_b_register_n24,
         oc8051_sfr1_oc8051_b_register_n23, oc8051_sfr1_oc8051_b_register_n22,
         oc8051_sfr1_oc8051_b_register_n21, oc8051_sfr1_oc8051_b_register_n20,
         oc8051_sfr1_oc8051_b_register_n19, oc8051_sfr1_oc8051_b_register_n18,
         oc8051_sfr1_oc8051_b_register_n17, oc8051_sfr1_oc8051_b_register_n16,
         oc8051_sfr1_oc8051_b_register_n15, oc8051_sfr1_oc8051_b_register_n14,
         oc8051_sfr1_oc8051_b_register_n13, oc8051_sfr1_oc8051_b_register_n12,
         oc8051_sfr1_oc8051_b_register_n11, oc8051_sfr1_oc8051_b_register_n10,
         oc8051_sfr1_oc8051_b_register_n9, oc8051_sfr1_oc8051_b_register_n8,
         oc8051_sfr1_oc8051_b_register_n7, oc8051_sfr1_oc8051_b_register_n6,
         oc8051_sfr1_oc8051_b_register_n5, oc8051_sfr1_oc8051_b_register_n4,
         oc8051_sfr1_oc8051_b_register_n3, oc8051_sfr1_oc8051_b_register_n2,
         oc8051_sfr1_oc8051_b_register_n1, oc8051_sfr1_oc8051_b_register_n39,
         oc8051_sfr1_oc8051_b_register_n38, oc8051_sfr1_oc8051_b_register_n37,
         oc8051_sfr1_oc8051_b_register_n36, oc8051_sfr1_oc8051_b_register_n35,
         oc8051_sfr1_oc8051_b_register_n34, oc8051_sfr1_oc8051_b_register_n33,
         oc8051_sfr1_oc8051_b_register_n32, oc8051_sfr1_oc8051_sp1_n37,
         oc8051_sfr1_oc8051_sp1_n36, oc8051_sfr1_oc8051_sp1_n35,
         oc8051_sfr1_oc8051_sp1_n34, oc8051_sfr1_oc8051_sp1_n33,
         oc8051_sfr1_oc8051_sp1_n32, oc8051_sfr1_oc8051_sp1_n31,
         oc8051_sfr1_oc8051_sp1_n30, oc8051_sfr1_oc8051_sp1_n29,
         oc8051_sfr1_oc8051_sp1_n28, oc8051_sfr1_oc8051_sp1_n27,
         oc8051_sfr1_oc8051_sp1_n26, oc8051_sfr1_oc8051_sp1_n25,
         oc8051_sfr1_oc8051_sp1_n24, oc8051_sfr1_oc8051_sp1_n23,
         oc8051_sfr1_oc8051_sp1_n21, oc8051_sfr1_oc8051_sp1_n20,
         oc8051_sfr1_oc8051_sp1_n19, oc8051_sfr1_oc8051_sp1_n18,
         oc8051_sfr1_oc8051_sp1_n17, oc8051_sfr1_oc8051_sp1_n16,
         oc8051_sfr1_oc8051_sp1_n15, oc8051_sfr1_oc8051_sp1_n14,
         oc8051_sfr1_oc8051_sp1_n13, oc8051_sfr1_oc8051_sp1_n12,
         oc8051_sfr1_oc8051_sp1_n11, oc8051_sfr1_oc8051_sp1_n10,
         oc8051_sfr1_oc8051_sp1_n9, oc8051_sfr1_oc8051_sp1_n8,
         oc8051_sfr1_oc8051_sp1_n7, oc8051_sfr1_oc8051_sp1_n6,
         oc8051_sfr1_oc8051_sp1_n5, oc8051_sfr1_oc8051_sp1_n4,
         oc8051_sfr1_oc8051_sp1_n3, oc8051_sfr1_oc8051_sp1_n2,
         oc8051_sfr1_oc8051_sp1_n1, oc8051_sfr1_oc8051_sp1_n22,
         oc8051_sfr1_oc8051_sp1_pop, oc8051_sfr1_oc8051_sp1_n200,
         oc8051_sfr1_oc8051_sp1_n190, oc8051_sfr1_oc8051_sp1_n180,
         oc8051_sfr1_oc8051_sp1_n170, oc8051_sfr1_oc8051_sp1_n160,
         oc8051_sfr1_oc8051_sp1_n150, oc8051_sfr1_oc8051_sp1_n140,
         oc8051_sfr1_oc8051_sp1_n130, oc8051_sfr1_oc8051_sp1_sp_0_,
         oc8051_sfr1_oc8051_sp1_sp_1_, oc8051_sfr1_oc8051_sp1_sp_2_,
         oc8051_sfr1_oc8051_sp1_sp_3_, oc8051_sfr1_oc8051_sp1_sp_4_,
         oc8051_sfr1_oc8051_sp1_sp_5_, oc8051_sfr1_oc8051_sp1_sp_6_,
         oc8051_sfr1_oc8051_sp1_sp_7_, oc8051_sfr1_oc8051_dptr1_n15,
         oc8051_sfr1_oc8051_dptr1_n14, oc8051_sfr1_oc8051_dptr1_n13,
         oc8051_sfr1_oc8051_dptr1_n12, oc8051_sfr1_oc8051_dptr1_n11,
         oc8051_sfr1_oc8051_dptr1_n10, oc8051_sfr1_oc8051_dptr1_n9,
         oc8051_sfr1_oc8051_dptr1_n8, oc8051_sfr1_oc8051_dptr1_n7,
         oc8051_sfr1_oc8051_dptr1_n6, oc8051_sfr1_oc8051_dptr1_n5,
         oc8051_sfr1_oc8051_dptr1_n4, oc8051_sfr1_oc8051_dptr1_n3,
         oc8051_sfr1_oc8051_dptr1_n2, oc8051_sfr1_oc8051_dptr1_n1,
         oc8051_sfr1_oc8051_dptr1_n33, oc8051_sfr1_oc8051_dptr1_n32,
         oc8051_sfr1_oc8051_dptr1_n31, oc8051_sfr1_oc8051_dptr1_n30,
         oc8051_sfr1_oc8051_dptr1_n29, oc8051_sfr1_oc8051_dptr1_n28,
         oc8051_sfr1_oc8051_dptr1_n27, oc8051_sfr1_oc8051_dptr1_n26,
         oc8051_sfr1_oc8051_dptr1_n25, oc8051_sfr1_oc8051_dptr1_n24,
         oc8051_sfr1_oc8051_dptr1_n23, oc8051_sfr1_oc8051_dptr1_n22,
         oc8051_sfr1_oc8051_dptr1_n21, oc8051_sfr1_oc8051_dptr1_n20,
         oc8051_sfr1_oc8051_dptr1_n19, oc8051_sfr1_oc8051_dptr1_n18,
         oc8051_sfr1_oc8051_psw1_n40, oc8051_sfr1_oc8051_psw1_n39,
         oc8051_sfr1_oc8051_psw1_n38, oc8051_sfr1_oc8051_psw1_n37,
         oc8051_sfr1_oc8051_psw1_n36, oc8051_sfr1_oc8051_psw1_n35,
         oc8051_sfr1_oc8051_psw1_n34, oc8051_sfr1_oc8051_psw1_n33,
         oc8051_sfr1_oc8051_psw1_n32, oc8051_sfr1_oc8051_psw1_n31,
         oc8051_sfr1_oc8051_psw1_n30, oc8051_sfr1_oc8051_psw1_n29,
         oc8051_sfr1_oc8051_psw1_n28, oc8051_sfr1_oc8051_psw1_n27,
         oc8051_sfr1_oc8051_psw1_n26, oc8051_sfr1_oc8051_psw1_n25,
         oc8051_sfr1_oc8051_psw1_n24, oc8051_sfr1_oc8051_psw1_n23,
         oc8051_sfr1_oc8051_psw1_n22, oc8051_sfr1_oc8051_psw1_n21,
         oc8051_sfr1_oc8051_psw1_n20, oc8051_sfr1_oc8051_psw1_n19,
         oc8051_sfr1_oc8051_psw1_n18, oc8051_sfr1_oc8051_psw1_n17,
         oc8051_sfr1_oc8051_psw1_n16, oc8051_sfr1_oc8051_psw1_n15,
         oc8051_sfr1_oc8051_psw1_n14, oc8051_sfr1_oc8051_psw1_n13,
         oc8051_sfr1_oc8051_psw1_n12, oc8051_sfr1_oc8051_psw1_n11,
         oc8051_sfr1_oc8051_psw1_n10, oc8051_sfr1_oc8051_psw1_n9,
         oc8051_sfr1_oc8051_psw1_n8, oc8051_sfr1_oc8051_psw1_n7,
         oc8051_sfr1_oc8051_psw1_n6, oc8051_sfr1_oc8051_psw1_n5,
         oc8051_sfr1_oc8051_psw1_n4, oc8051_sfr1_oc8051_psw1_n3,
         oc8051_sfr1_oc8051_psw1_n2, oc8051_sfr1_oc8051_psw1_n49,
         oc8051_sfr1_oc8051_psw1_n48, oc8051_sfr1_oc8051_psw1_n47,
         oc8051_sfr1_oc8051_psw1_n46, oc8051_sfr1_oc8051_psw1_n45,
         oc8051_sfr1_oc8051_psw1_n44, oc8051_sfr1_oc8051_psw1_n43,
         oc8051_sfr1_oc8051_psw1_n1, oc8051_sfr1_oc8051_ports1_n106,
         oc8051_sfr1_oc8051_ports1_n105, oc8051_sfr1_oc8051_ports1_n104,
         oc8051_sfr1_oc8051_ports1_n103, oc8051_sfr1_oc8051_ports1_n102,
         oc8051_sfr1_oc8051_ports1_n101, oc8051_sfr1_oc8051_ports1_n100,
         oc8051_sfr1_oc8051_ports1_n99, oc8051_sfr1_oc8051_ports1_n98,
         oc8051_sfr1_oc8051_ports1_n97, oc8051_sfr1_oc8051_ports1_n96,
         oc8051_sfr1_oc8051_ports1_n95, oc8051_sfr1_oc8051_ports1_n94,
         oc8051_sfr1_oc8051_ports1_n93, oc8051_sfr1_oc8051_ports1_n92,
         oc8051_sfr1_oc8051_ports1_n91, oc8051_sfr1_oc8051_ports1_n90,
         oc8051_sfr1_oc8051_ports1_n89, oc8051_sfr1_oc8051_ports1_n88,
         oc8051_sfr1_oc8051_ports1_n87, oc8051_sfr1_oc8051_ports1_n86,
         oc8051_sfr1_oc8051_ports1_n85, oc8051_sfr1_oc8051_ports1_n84,
         oc8051_sfr1_oc8051_ports1_n83, oc8051_sfr1_oc8051_ports1_n82,
         oc8051_sfr1_oc8051_ports1_n81, oc8051_sfr1_oc8051_ports1_n80,
         oc8051_sfr1_oc8051_ports1_n79, oc8051_sfr1_oc8051_ports1_n78,
         oc8051_sfr1_oc8051_ports1_n77, oc8051_sfr1_oc8051_ports1_n76,
         oc8051_sfr1_oc8051_ports1_n75, oc8051_sfr1_oc8051_ports1_n74,
         oc8051_sfr1_oc8051_ports1_n73, oc8051_sfr1_oc8051_ports1_n72,
         oc8051_sfr1_oc8051_ports1_n71, oc8051_sfr1_oc8051_ports1_n70,
         oc8051_sfr1_oc8051_ports1_n69, oc8051_sfr1_oc8051_ports1_n68,
         oc8051_sfr1_oc8051_ports1_n67, oc8051_sfr1_oc8051_ports1_n66,
         oc8051_sfr1_oc8051_ports1_n65, oc8051_sfr1_oc8051_ports1_n64,
         oc8051_sfr1_oc8051_ports1_n63, oc8051_sfr1_oc8051_ports1_n62,
         oc8051_sfr1_oc8051_ports1_n61, oc8051_sfr1_oc8051_ports1_n60,
         oc8051_sfr1_oc8051_ports1_n59, oc8051_sfr1_oc8051_ports1_n58,
         oc8051_sfr1_oc8051_ports1_n57, oc8051_sfr1_oc8051_ports1_n56,
         oc8051_sfr1_oc8051_ports1_n55, oc8051_sfr1_oc8051_ports1_n54,
         oc8051_sfr1_oc8051_ports1_n53, oc8051_sfr1_oc8051_ports1_n52,
         oc8051_sfr1_oc8051_ports1_n51, oc8051_sfr1_oc8051_ports1_n50,
         oc8051_sfr1_oc8051_ports1_n49, oc8051_sfr1_oc8051_ports1_n48,
         oc8051_sfr1_oc8051_ports1_n47, oc8051_sfr1_oc8051_ports1_n46,
         oc8051_sfr1_oc8051_ports1_n45, oc8051_sfr1_oc8051_ports1_n44,
         oc8051_sfr1_oc8051_ports1_n43, oc8051_sfr1_oc8051_ports1_n42,
         oc8051_sfr1_oc8051_ports1_n41, oc8051_sfr1_oc8051_ports1_n40,
         oc8051_sfr1_oc8051_ports1_n39, oc8051_sfr1_oc8051_ports1_n38,
         oc8051_sfr1_oc8051_ports1_n37, oc8051_sfr1_oc8051_ports1_n36,
         oc8051_sfr1_oc8051_ports1_n35, oc8051_sfr1_oc8051_ports1_n34,
         oc8051_sfr1_oc8051_ports1_n33, oc8051_sfr1_oc8051_ports1_n32,
         oc8051_sfr1_oc8051_ports1_n31, oc8051_sfr1_oc8051_ports1_n30,
         oc8051_sfr1_oc8051_ports1_n29, oc8051_sfr1_oc8051_ports1_n28,
         oc8051_sfr1_oc8051_ports1_n27, oc8051_sfr1_oc8051_ports1_n26,
         oc8051_sfr1_oc8051_ports1_n25, oc8051_sfr1_oc8051_ports1_n24,
         oc8051_sfr1_oc8051_ports1_n23, oc8051_sfr1_oc8051_ports1_n22,
         oc8051_sfr1_oc8051_ports1_n21, oc8051_sfr1_oc8051_ports1_n20,
         oc8051_sfr1_oc8051_ports1_n19, oc8051_sfr1_oc8051_ports1_n18,
         oc8051_sfr1_oc8051_ports1_n17, oc8051_sfr1_oc8051_ports1_n16,
         oc8051_sfr1_oc8051_ports1_n15, oc8051_sfr1_oc8051_ports1_n14,
         oc8051_sfr1_oc8051_ports1_n13, oc8051_sfr1_oc8051_ports1_n12,
         oc8051_sfr1_oc8051_ports1_n11, oc8051_sfr1_oc8051_ports1_n10,
         oc8051_sfr1_oc8051_ports1_n9, oc8051_sfr1_oc8051_ports1_n8,
         oc8051_sfr1_oc8051_ports1_n7, oc8051_sfr1_oc8051_ports1_n6,
         oc8051_sfr1_oc8051_ports1_n5, oc8051_sfr1_oc8051_ports1_n4,
         oc8051_sfr1_oc8051_ports1_n3, oc8051_sfr1_oc8051_ports1_n2,
         oc8051_sfr1_oc8051_ports1_n1, oc8051_sfr1_oc8051_ports1_n163,
         oc8051_sfr1_oc8051_ports1_n162, oc8051_sfr1_oc8051_ports1_n161,
         oc8051_sfr1_oc8051_ports1_n160, oc8051_sfr1_oc8051_ports1_n159,
         oc8051_sfr1_oc8051_ports1_n158, oc8051_sfr1_oc8051_ports1_n157,
         oc8051_sfr1_oc8051_ports1_n156, oc8051_sfr1_oc8051_ports1_n155,
         oc8051_sfr1_oc8051_ports1_n154, oc8051_sfr1_oc8051_ports1_n153,
         oc8051_sfr1_oc8051_ports1_n152, oc8051_sfr1_oc8051_ports1_n151,
         oc8051_sfr1_oc8051_ports1_n150, oc8051_sfr1_oc8051_ports1_n149,
         oc8051_sfr1_oc8051_ports1_n148, oc8051_sfr1_oc8051_ports1_n147,
         oc8051_sfr1_oc8051_ports1_n146, oc8051_sfr1_oc8051_ports1_n145,
         oc8051_sfr1_oc8051_ports1_n144, oc8051_sfr1_oc8051_ports1_n143,
         oc8051_sfr1_oc8051_ports1_n142, oc8051_sfr1_oc8051_ports1_n141,
         oc8051_sfr1_oc8051_ports1_n140, oc8051_sfr1_oc8051_ports1_n139,
         oc8051_sfr1_oc8051_ports1_n138, oc8051_sfr1_oc8051_ports1_n137,
         oc8051_sfr1_oc8051_ports1_n136, oc8051_sfr1_oc8051_ports1_n135,
         oc8051_sfr1_oc8051_ports1_n134, oc8051_sfr1_oc8051_ports1_n133,
         oc8051_sfr1_oc8051_ports1_n132, oc8051_sfr1_oc8051_uatr1_n172,
         oc8051_sfr1_oc8051_uatr1_n170, oc8051_sfr1_oc8051_uatr1_n169,
         oc8051_sfr1_oc8051_uatr1_n168, oc8051_sfr1_oc8051_uatr1_n167,
         oc8051_sfr1_oc8051_uatr1_n166, oc8051_sfr1_oc8051_uatr1_n165,
         oc8051_sfr1_oc8051_uatr1_n164, oc8051_sfr1_oc8051_uatr1_n163,
         oc8051_sfr1_oc8051_uatr1_n162, oc8051_sfr1_oc8051_uatr1_n161,
         oc8051_sfr1_oc8051_uatr1_n160, oc8051_sfr1_oc8051_uatr1_n159,
         oc8051_sfr1_oc8051_uatr1_n158, oc8051_sfr1_oc8051_uatr1_n157,
         oc8051_sfr1_oc8051_uatr1_n156, oc8051_sfr1_oc8051_uatr1_n155,
         oc8051_sfr1_oc8051_uatr1_n154, oc8051_sfr1_oc8051_uatr1_n153,
         oc8051_sfr1_oc8051_uatr1_n152, oc8051_sfr1_oc8051_uatr1_n151,
         oc8051_sfr1_oc8051_uatr1_n150, oc8051_sfr1_oc8051_uatr1_n149,
         oc8051_sfr1_oc8051_uatr1_n148, oc8051_sfr1_oc8051_uatr1_n147,
         oc8051_sfr1_oc8051_uatr1_n146, oc8051_sfr1_oc8051_uatr1_n145,
         oc8051_sfr1_oc8051_uatr1_n144, oc8051_sfr1_oc8051_uatr1_n143,
         oc8051_sfr1_oc8051_uatr1_n142, oc8051_sfr1_oc8051_uatr1_n141,
         oc8051_sfr1_oc8051_uatr1_n140, oc8051_sfr1_oc8051_uatr1_n139,
         oc8051_sfr1_oc8051_uatr1_n138, oc8051_sfr1_oc8051_uatr1_n137,
         oc8051_sfr1_oc8051_uatr1_n136, oc8051_sfr1_oc8051_uatr1_n135,
         oc8051_sfr1_oc8051_uatr1_n134, oc8051_sfr1_oc8051_uatr1_n133,
         oc8051_sfr1_oc8051_uatr1_n132, oc8051_sfr1_oc8051_uatr1_n131,
         oc8051_sfr1_oc8051_uatr1_n130, oc8051_sfr1_oc8051_uatr1_n129,
         oc8051_sfr1_oc8051_uatr1_n128, oc8051_sfr1_oc8051_uatr1_n127,
         oc8051_sfr1_oc8051_uatr1_n126, oc8051_sfr1_oc8051_uatr1_n125,
         oc8051_sfr1_oc8051_uatr1_n124, oc8051_sfr1_oc8051_uatr1_n123,
         oc8051_sfr1_oc8051_uatr1_n122, oc8051_sfr1_oc8051_uatr1_n121,
         oc8051_sfr1_oc8051_uatr1_n120, oc8051_sfr1_oc8051_uatr1_n119,
         oc8051_sfr1_oc8051_uatr1_n118, oc8051_sfr1_oc8051_uatr1_n117,
         oc8051_sfr1_oc8051_uatr1_n116, oc8051_sfr1_oc8051_uatr1_n115,
         oc8051_sfr1_oc8051_uatr1_n114, oc8051_sfr1_oc8051_uatr1_n113,
         oc8051_sfr1_oc8051_uatr1_n112, oc8051_sfr1_oc8051_uatr1_n111,
         oc8051_sfr1_oc8051_uatr1_n110, oc8051_sfr1_oc8051_uatr1_n109,
         oc8051_sfr1_oc8051_uatr1_n108, oc8051_sfr1_oc8051_uatr1_n107,
         oc8051_sfr1_oc8051_uatr1_n106, oc8051_sfr1_oc8051_uatr1_n105,
         oc8051_sfr1_oc8051_uatr1_n104, oc8051_sfr1_oc8051_uatr1_n103,
         oc8051_sfr1_oc8051_uatr1_n102, oc8051_sfr1_oc8051_uatr1_n101,
         oc8051_sfr1_oc8051_uatr1_n100, oc8051_sfr1_oc8051_uatr1_n99,
         oc8051_sfr1_oc8051_uatr1_n98, oc8051_sfr1_oc8051_uatr1_n97,
         oc8051_sfr1_oc8051_uatr1_n96, oc8051_sfr1_oc8051_uatr1_n95,
         oc8051_sfr1_oc8051_uatr1_n94, oc8051_sfr1_oc8051_uatr1_n93,
         oc8051_sfr1_oc8051_uatr1_n92, oc8051_sfr1_oc8051_uatr1_n91,
         oc8051_sfr1_oc8051_uatr1_n90, oc8051_sfr1_oc8051_uatr1_n89,
         oc8051_sfr1_oc8051_uatr1_n88, oc8051_sfr1_oc8051_uatr1_n87,
         oc8051_sfr1_oc8051_uatr1_n86, oc8051_sfr1_oc8051_uatr1_n85,
         oc8051_sfr1_oc8051_uatr1_n84, oc8051_sfr1_oc8051_uatr1_n83,
         oc8051_sfr1_oc8051_uatr1_n82, oc8051_sfr1_oc8051_uatr1_n81,
         oc8051_sfr1_oc8051_uatr1_n80, oc8051_sfr1_oc8051_uatr1_n79,
         oc8051_sfr1_oc8051_uatr1_n78, oc8051_sfr1_oc8051_uatr1_n77,
         oc8051_sfr1_oc8051_uatr1_n76, oc8051_sfr1_oc8051_uatr1_n75,
         oc8051_sfr1_oc8051_uatr1_n74, oc8051_sfr1_oc8051_uatr1_n73,
         oc8051_sfr1_oc8051_uatr1_n72, oc8051_sfr1_oc8051_uatr1_n71,
         oc8051_sfr1_oc8051_uatr1_n70, oc8051_sfr1_oc8051_uatr1_n69,
         oc8051_sfr1_oc8051_uatr1_n68, oc8051_sfr1_oc8051_uatr1_n67,
         oc8051_sfr1_oc8051_uatr1_n66, oc8051_sfr1_oc8051_uatr1_n65,
         oc8051_sfr1_oc8051_uatr1_n64, oc8051_sfr1_oc8051_uatr1_n63,
         oc8051_sfr1_oc8051_uatr1_n62, oc8051_sfr1_oc8051_uatr1_n61,
         oc8051_sfr1_oc8051_uatr1_n60, oc8051_sfr1_oc8051_uatr1_n59,
         oc8051_sfr1_oc8051_uatr1_n58, oc8051_sfr1_oc8051_uatr1_n57,
         oc8051_sfr1_oc8051_uatr1_n56, oc8051_sfr1_oc8051_uatr1_n55,
         oc8051_sfr1_oc8051_uatr1_n54, oc8051_sfr1_oc8051_uatr1_n53,
         oc8051_sfr1_oc8051_uatr1_n52, oc8051_sfr1_oc8051_uatr1_n51,
         oc8051_sfr1_oc8051_uatr1_n50, oc8051_sfr1_oc8051_uatr1_n49,
         oc8051_sfr1_oc8051_uatr1_n48, oc8051_sfr1_oc8051_uatr1_n47,
         oc8051_sfr1_oc8051_uatr1_n46, oc8051_sfr1_oc8051_uatr1_n45,
         oc8051_sfr1_oc8051_uatr1_n44, oc8051_sfr1_oc8051_uatr1_n43,
         oc8051_sfr1_oc8051_uatr1_n42, oc8051_sfr1_oc8051_uatr1_n41,
         oc8051_sfr1_oc8051_uatr1_n40, oc8051_sfr1_oc8051_uatr1_n39,
         oc8051_sfr1_oc8051_uatr1_n38, oc8051_sfr1_oc8051_uatr1_n37,
         oc8051_sfr1_oc8051_uatr1_n36, oc8051_sfr1_oc8051_uatr1_n35,
         oc8051_sfr1_oc8051_uatr1_n34, oc8051_sfr1_oc8051_uatr1_n33,
         oc8051_sfr1_oc8051_uatr1_n32, oc8051_sfr1_oc8051_uatr1_n31,
         oc8051_sfr1_oc8051_uatr1_n30, oc8051_sfr1_oc8051_uatr1_n29,
         oc8051_sfr1_oc8051_uatr1_n28, oc8051_sfr1_oc8051_uatr1_n27,
         oc8051_sfr1_oc8051_uatr1_n26, oc8051_sfr1_oc8051_uatr1_n25,
         oc8051_sfr1_oc8051_uatr1_n24, oc8051_sfr1_oc8051_uatr1_n23,
         oc8051_sfr1_oc8051_uatr1_n22, oc8051_sfr1_oc8051_uatr1_n21,
         oc8051_sfr1_oc8051_uatr1_n20, oc8051_sfr1_oc8051_uatr1_n19,
         oc8051_sfr1_oc8051_uatr1_n18, oc8051_sfr1_oc8051_uatr1_n17,
         oc8051_sfr1_oc8051_uatr1_n16, oc8051_sfr1_oc8051_uatr1_n15,
         oc8051_sfr1_oc8051_uatr1_n14, oc8051_sfr1_oc8051_uatr1_n13,
         oc8051_sfr1_oc8051_uatr1_n12, oc8051_sfr1_oc8051_uatr1_n11,
         oc8051_sfr1_oc8051_uatr1_n10, oc8051_sfr1_oc8051_uatr1_n9,
         oc8051_sfr1_oc8051_uatr1_n8, oc8051_sfr1_oc8051_uatr1_n7,
         oc8051_sfr1_oc8051_uatr1_n6, oc8051_sfr1_oc8051_uatr1_n5,
         oc8051_sfr1_oc8051_uatr1_n4, oc8051_sfr1_oc8051_uatr1_n3,
         oc8051_sfr1_oc8051_uatr1_n2, oc8051_sfr1_oc8051_uatr1_n1,
         oc8051_sfr1_oc8051_uatr1_n254, oc8051_sfr1_oc8051_uatr1_n253,
         oc8051_sfr1_oc8051_uatr1_n252, oc8051_sfr1_oc8051_uatr1_n251,
         oc8051_sfr1_oc8051_uatr1_n250, oc8051_sfr1_oc8051_uatr1_n249,
         oc8051_sfr1_oc8051_uatr1_n248, oc8051_sfr1_oc8051_uatr1_n247,
         oc8051_sfr1_oc8051_uatr1_n246, oc8051_sfr1_oc8051_uatr1_n245,
         oc8051_sfr1_oc8051_uatr1_n244, oc8051_sfr1_oc8051_uatr1_n243,
         oc8051_sfr1_oc8051_uatr1_n242, oc8051_sfr1_oc8051_uatr1_n240,
         oc8051_sfr1_oc8051_uatr1_n239, oc8051_sfr1_oc8051_uatr1_n238,
         oc8051_sfr1_oc8051_uatr1_n237, oc8051_sfr1_oc8051_uatr1_n236,
         oc8051_sfr1_oc8051_uatr1_n235, oc8051_sfr1_oc8051_uatr1_n234,
         oc8051_sfr1_oc8051_uatr1_n233, oc8051_sfr1_oc8051_uatr1_n232,
         oc8051_sfr1_oc8051_uatr1_n231, oc8051_sfr1_oc8051_uatr1_n230,
         oc8051_sfr1_oc8051_uatr1_n229, oc8051_sfr1_oc8051_uatr1_n228,
         oc8051_sfr1_oc8051_uatr1_n227, oc8051_sfr1_oc8051_uatr1_n226,
         oc8051_sfr1_oc8051_uatr1_n225, oc8051_sfr1_oc8051_uatr1_n224,
         oc8051_sfr1_oc8051_uatr1_n223, oc8051_sfr1_oc8051_uatr1_n222,
         oc8051_sfr1_oc8051_uatr1_n221, oc8051_sfr1_oc8051_uatr1_n220,
         oc8051_sfr1_oc8051_uatr1_n219, oc8051_sfr1_oc8051_uatr1_n218,
         oc8051_sfr1_oc8051_uatr1_n217, oc8051_sfr1_oc8051_uatr1_n216,
         oc8051_sfr1_oc8051_uatr1_n215, oc8051_sfr1_oc8051_uatr1_n214,
         oc8051_sfr1_oc8051_uatr1_n213, oc8051_sfr1_oc8051_uatr1_n212,
         oc8051_sfr1_oc8051_uatr1_n211, oc8051_sfr1_oc8051_uatr1_n210,
         oc8051_sfr1_oc8051_uatr1_n209, oc8051_sfr1_oc8051_uatr1_n208,
         oc8051_sfr1_oc8051_uatr1_n207, oc8051_sfr1_oc8051_uatr1_n206,
         oc8051_sfr1_oc8051_uatr1_n205, oc8051_sfr1_oc8051_uatr1_n204,
         oc8051_sfr1_oc8051_uatr1_n203, oc8051_sfr1_oc8051_uatr1_n202,
         oc8051_sfr1_oc8051_uatr1_n201, oc8051_sfr1_oc8051_uatr1_n200,
         oc8051_sfr1_oc8051_uatr1_n199, oc8051_sfr1_oc8051_uatr1_n198,
         oc8051_sfr1_oc8051_uatr1_n197, oc8051_sfr1_oc8051_uatr1_n196,
         oc8051_sfr1_oc8051_uatr1_n195, oc8051_sfr1_oc8051_uatr1_n194,
         oc8051_sfr1_oc8051_uatr1_n193, oc8051_sfr1_oc8051_uatr1_n192,
         oc8051_sfr1_oc8051_uatr1_n191, oc8051_sfr1_oc8051_uatr1_n190,
         oc8051_sfr1_oc8051_uatr1_n188, oc8051_sfr1_oc8051_uatr1_n187,
         oc8051_sfr1_oc8051_uatr1_n186, oc8051_sfr1_oc8051_uatr1_n185,
         oc8051_sfr1_oc8051_uatr1_n184, oc8051_sfr1_oc8051_uatr1_n183,
         oc8051_sfr1_oc8051_uatr1_n182, oc8051_sfr1_oc8051_uatr1_n181,
         oc8051_sfr1_oc8051_uatr1_n180, oc8051_sfr1_oc8051_uatr1_n269,
         oc8051_sfr1_oc8051_uatr1_smod_clk_re, oc8051_sfr1_oc8051_uatr1_rxd_r,
         oc8051_sfr1_oc8051_uatr1_shift_re, oc8051_sfr1_oc8051_uatr1_rx_sam_0_,
         oc8051_sfr1_oc8051_uatr1_rx_sam_1_,
         oc8051_sfr1_oc8051_uatr1_re_count_0_,
         oc8051_sfr1_oc8051_uatr1_re_count_1_,
         oc8051_sfr1_oc8051_uatr1_re_count_2_,
         oc8051_sfr1_oc8051_uatr1_re_count_3_,
         oc8051_sfr1_oc8051_uatr1_receive, oc8051_sfr1_oc8051_uatr1_n174,
         oc8051_sfr1_oc8051_uatr1_smod_clk_tr,
         oc8051_sfr1_oc8051_uatr1_shift_tr,
         oc8051_sfr1_oc8051_uatr1_tr_count_0_,
         oc8051_sfr1_oc8051_uatr1_tr_count_1_,
         oc8051_sfr1_oc8051_uatr1_tr_count_2_, oc8051_sfr1_oc8051_uatr1_trans,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_6_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_7_,
         oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_,
         oc8051_sfr1_oc8051_uatr1_rx_done,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_,
         oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_,
         oc8051_sfr1_oc8051_int1_n209, oc8051_sfr1_oc8051_int1_n208,
         oc8051_sfr1_oc8051_int1_n207, oc8051_sfr1_oc8051_int1_n206,
         oc8051_sfr1_oc8051_int1_n205, oc8051_sfr1_oc8051_int1_n204,
         oc8051_sfr1_oc8051_int1_n203, oc8051_sfr1_oc8051_int1_n202,
         oc8051_sfr1_oc8051_int1_n201, oc8051_sfr1_oc8051_int1_n200,
         oc8051_sfr1_oc8051_int1_n199, oc8051_sfr1_oc8051_int1_n198,
         oc8051_sfr1_oc8051_int1_n197, oc8051_sfr1_oc8051_int1_n196,
         oc8051_sfr1_oc8051_int1_n195, oc8051_sfr1_oc8051_int1_n194,
         oc8051_sfr1_oc8051_int1_n193, oc8051_sfr1_oc8051_int1_n192,
         oc8051_sfr1_oc8051_int1_n191, oc8051_sfr1_oc8051_int1_n190,
         oc8051_sfr1_oc8051_int1_n189, oc8051_sfr1_oc8051_int1_n188,
         oc8051_sfr1_oc8051_int1_n187, oc8051_sfr1_oc8051_int1_n186,
         oc8051_sfr1_oc8051_int1_n185, oc8051_sfr1_oc8051_int1_n184,
         oc8051_sfr1_oc8051_int1_n183, oc8051_sfr1_oc8051_int1_n182,
         oc8051_sfr1_oc8051_int1_n181, oc8051_sfr1_oc8051_int1_n180,
         oc8051_sfr1_oc8051_int1_n179, oc8051_sfr1_oc8051_int1_n178,
         oc8051_sfr1_oc8051_int1_n177, oc8051_sfr1_oc8051_int1_n176,
         oc8051_sfr1_oc8051_int1_n175, oc8051_sfr1_oc8051_int1_n174,
         oc8051_sfr1_oc8051_int1_n173, oc8051_sfr1_oc8051_int1_n172,
         oc8051_sfr1_oc8051_int1_n171, oc8051_sfr1_oc8051_int1_n170,
         oc8051_sfr1_oc8051_int1_n169, oc8051_sfr1_oc8051_int1_n168,
         oc8051_sfr1_oc8051_int1_n167, oc8051_sfr1_oc8051_int1_n166,
         oc8051_sfr1_oc8051_int1_n165, oc8051_sfr1_oc8051_int1_n164,
         oc8051_sfr1_oc8051_int1_n163, oc8051_sfr1_oc8051_int1_n162,
         oc8051_sfr1_oc8051_int1_n161, oc8051_sfr1_oc8051_int1_n160,
         oc8051_sfr1_oc8051_int1_n159, oc8051_sfr1_oc8051_int1_n158,
         oc8051_sfr1_oc8051_int1_n157, oc8051_sfr1_oc8051_int1_n156,
         oc8051_sfr1_oc8051_int1_n155, oc8051_sfr1_oc8051_int1_n154,
         oc8051_sfr1_oc8051_int1_n153, oc8051_sfr1_oc8051_int1_n152,
         oc8051_sfr1_oc8051_int1_n151, oc8051_sfr1_oc8051_int1_n150,
         oc8051_sfr1_oc8051_int1_n149, oc8051_sfr1_oc8051_int1_n148,
         oc8051_sfr1_oc8051_int1_n147, oc8051_sfr1_oc8051_int1_n146,
         oc8051_sfr1_oc8051_int1_n145, oc8051_sfr1_oc8051_int1_n144,
         oc8051_sfr1_oc8051_int1_n143, oc8051_sfr1_oc8051_int1_n142,
         oc8051_sfr1_oc8051_int1_n141, oc8051_sfr1_oc8051_int1_n140,
         oc8051_sfr1_oc8051_int1_n139, oc8051_sfr1_oc8051_int1_n138,
         oc8051_sfr1_oc8051_int1_n137, oc8051_sfr1_oc8051_int1_n136,
         oc8051_sfr1_oc8051_int1_n135, oc8051_sfr1_oc8051_int1_n134,
         oc8051_sfr1_oc8051_int1_n133, oc8051_sfr1_oc8051_int1_n132,
         oc8051_sfr1_oc8051_int1_n131, oc8051_sfr1_oc8051_int1_n130,
         oc8051_sfr1_oc8051_int1_n129, oc8051_sfr1_oc8051_int1_n128,
         oc8051_sfr1_oc8051_int1_n127, oc8051_sfr1_oc8051_int1_n126,
         oc8051_sfr1_oc8051_int1_n125, oc8051_sfr1_oc8051_int1_n124,
         oc8051_sfr1_oc8051_int1_n123, oc8051_sfr1_oc8051_int1_n122,
         oc8051_sfr1_oc8051_int1_n121, oc8051_sfr1_oc8051_int1_n120,
         oc8051_sfr1_oc8051_int1_n119, oc8051_sfr1_oc8051_int1_n118,
         oc8051_sfr1_oc8051_int1_n117, oc8051_sfr1_oc8051_int1_n116,
         oc8051_sfr1_oc8051_int1_n115, oc8051_sfr1_oc8051_int1_n114,
         oc8051_sfr1_oc8051_int1_n113, oc8051_sfr1_oc8051_int1_n112,
         oc8051_sfr1_oc8051_int1_n111, oc8051_sfr1_oc8051_int1_n110,
         oc8051_sfr1_oc8051_int1_n109, oc8051_sfr1_oc8051_int1_n108,
         oc8051_sfr1_oc8051_int1_n107, oc8051_sfr1_oc8051_int1_n106,
         oc8051_sfr1_oc8051_int1_n105, oc8051_sfr1_oc8051_int1_n104,
         oc8051_sfr1_oc8051_int1_n103, oc8051_sfr1_oc8051_int1_n102,
         oc8051_sfr1_oc8051_int1_n101, oc8051_sfr1_oc8051_int1_n100,
         oc8051_sfr1_oc8051_int1_n99, oc8051_sfr1_oc8051_int1_n98,
         oc8051_sfr1_oc8051_int1_n97, oc8051_sfr1_oc8051_int1_n96,
         oc8051_sfr1_oc8051_int1_n95, oc8051_sfr1_oc8051_int1_n94,
         oc8051_sfr1_oc8051_int1_n93, oc8051_sfr1_oc8051_int1_n92,
         oc8051_sfr1_oc8051_int1_n91, oc8051_sfr1_oc8051_int1_n90,
         oc8051_sfr1_oc8051_int1_n89, oc8051_sfr1_oc8051_int1_n88,
         oc8051_sfr1_oc8051_int1_n87, oc8051_sfr1_oc8051_int1_n86,
         oc8051_sfr1_oc8051_int1_n85, oc8051_sfr1_oc8051_int1_n84,
         oc8051_sfr1_oc8051_int1_n83, oc8051_sfr1_oc8051_int1_n82,
         oc8051_sfr1_oc8051_int1_n81, oc8051_sfr1_oc8051_int1_n80,
         oc8051_sfr1_oc8051_int1_n79, oc8051_sfr1_oc8051_int1_n78,
         oc8051_sfr1_oc8051_int1_n77, oc8051_sfr1_oc8051_int1_n76,
         oc8051_sfr1_oc8051_int1_n75, oc8051_sfr1_oc8051_int1_n74,
         oc8051_sfr1_oc8051_int1_n73, oc8051_sfr1_oc8051_int1_n72,
         oc8051_sfr1_oc8051_int1_n71, oc8051_sfr1_oc8051_int1_n70,
         oc8051_sfr1_oc8051_int1_n69, oc8051_sfr1_oc8051_int1_n68,
         oc8051_sfr1_oc8051_int1_n67, oc8051_sfr1_oc8051_int1_n66,
         oc8051_sfr1_oc8051_int1_n65, oc8051_sfr1_oc8051_int1_n64,
         oc8051_sfr1_oc8051_int1_n63, oc8051_sfr1_oc8051_int1_n62,
         oc8051_sfr1_oc8051_int1_n61, oc8051_sfr1_oc8051_int1_n60,
         oc8051_sfr1_oc8051_int1_n59, oc8051_sfr1_oc8051_int1_n58,
         oc8051_sfr1_oc8051_int1_n57, oc8051_sfr1_oc8051_int1_n56,
         oc8051_sfr1_oc8051_int1_n55, oc8051_sfr1_oc8051_int1_n54,
         oc8051_sfr1_oc8051_int1_n51, oc8051_sfr1_oc8051_int1_n50,
         oc8051_sfr1_oc8051_int1_n44, oc8051_sfr1_oc8051_int1_n42,
         oc8051_sfr1_oc8051_int1_n41, oc8051_sfr1_oc8051_int1_n40,
         oc8051_sfr1_oc8051_int1_n39, oc8051_sfr1_oc8051_int1_n38,
         oc8051_sfr1_oc8051_int1_n37, oc8051_sfr1_oc8051_int1_n36,
         oc8051_sfr1_oc8051_int1_n35, oc8051_sfr1_oc8051_int1_n34,
         oc8051_sfr1_oc8051_int1_n33, oc8051_sfr1_oc8051_int1_n32,
         oc8051_sfr1_oc8051_int1_n31, oc8051_sfr1_oc8051_int1_n30,
         oc8051_sfr1_oc8051_int1_n29, oc8051_sfr1_oc8051_int1_n28,
         oc8051_sfr1_oc8051_int1_n27, oc8051_sfr1_oc8051_int1_n26,
         oc8051_sfr1_oc8051_int1_n25, oc8051_sfr1_oc8051_int1_n24,
         oc8051_sfr1_oc8051_int1_n23, oc8051_sfr1_oc8051_int1_n22,
         oc8051_sfr1_oc8051_int1_n21, oc8051_sfr1_oc8051_int1_n20,
         oc8051_sfr1_oc8051_int1_n19, oc8051_sfr1_oc8051_int1_n18,
         oc8051_sfr1_oc8051_int1_n17, oc8051_sfr1_oc8051_int1_n16,
         oc8051_sfr1_oc8051_int1_n15, oc8051_sfr1_oc8051_int1_n14,
         oc8051_sfr1_oc8051_int1_n13, oc8051_sfr1_oc8051_int1_n12,
         oc8051_sfr1_oc8051_int1_n11, oc8051_sfr1_oc8051_int1_n10,
         oc8051_sfr1_oc8051_int1_n3, oc8051_sfr1_oc8051_int1_n2,
         oc8051_sfr1_oc8051_int1_int_vec_2_, oc8051_sfr1_oc8051_int1_n274,
         oc8051_sfr1_oc8051_int1_n273, oc8051_sfr1_oc8051_int1_n272,
         oc8051_sfr1_oc8051_int1_n271, oc8051_sfr1_oc8051_int1_n270,
         oc8051_sfr1_oc8051_int1_n269, oc8051_sfr1_oc8051_int1_n268,
         oc8051_sfr1_oc8051_int1_n267, oc8051_sfr1_oc8051_int1_n266,
         oc8051_sfr1_oc8051_int1_n265, oc8051_sfr1_oc8051_int1_n264,
         oc8051_sfr1_oc8051_int1_n263, oc8051_sfr1_oc8051_int1_n262,
         oc8051_sfr1_oc8051_int1_n261, oc8051_sfr1_oc8051_int1_n260,
         oc8051_sfr1_oc8051_int1_n259, oc8051_sfr1_oc8051_int1_n258,
         oc8051_sfr1_oc8051_int1_n257, oc8051_sfr1_oc8051_int1_n256,
         oc8051_sfr1_oc8051_int1_n255, oc8051_sfr1_oc8051_int1_n254,
         oc8051_sfr1_oc8051_int1_n253, oc8051_sfr1_oc8051_int1_n252,
         oc8051_sfr1_oc8051_int1_n251, oc8051_sfr1_oc8051_int1_n250,
         oc8051_sfr1_oc8051_int1_n249, oc8051_sfr1_oc8051_int1_n248,
         oc8051_sfr1_oc8051_int1_n247, oc8051_sfr1_oc8051_int1_n246,
         oc8051_sfr1_oc8051_int1_n245, oc8051_sfr1_oc8051_int1_n244,
         oc8051_sfr1_oc8051_int1_n243, oc8051_sfr1_oc8051_int1_n242,
         oc8051_sfr1_oc8051_int1_n241, oc8051_sfr1_oc8051_int1_n240,
         oc8051_sfr1_oc8051_int1_n239, oc8051_sfr1_oc8051_int1_n238,
         oc8051_sfr1_oc8051_int1_n237, oc8051_sfr1_oc8051_int1_n236,
         oc8051_sfr1_oc8051_int1_n235, oc8051_sfr1_oc8051_int1_n53,
         oc8051_sfr1_oc8051_int1_n52, oc8051_sfr1_oc8051_int1_n49,
         oc8051_sfr1_oc8051_int1_n48, oc8051_sfr1_oc8051_int1_n47,
         oc8051_sfr1_oc8051_int1_n46, oc8051_sfr1_oc8051_int1_n45,
         oc8051_sfr1_oc8051_int1_n43, oc8051_sfr1_oc8051_int1_n9,
         oc8051_sfr1_oc8051_int1_n8, oc8051_sfr1_oc8051_int1_n7,
         oc8051_sfr1_oc8051_int1_n6, oc8051_sfr1_oc8051_int1_n5,
         oc8051_sfr1_oc8051_int1_n4, oc8051_sfr1_oc8051_int1_ie1_buff,
         oc8051_sfr1_oc8051_int1_ie0_buff, oc8051_sfr1_oc8051_int1_tf0_buff,
         oc8051_sfr1_oc8051_int1_tf1_buff, oc8051_sfr1_oc8051_int1_int_dept_0_,
         oc8051_sfr1_oc8051_int1_int_dept_1_, oc8051_sfr1_oc8051_int1_int_proc,
         oc8051_sfr1_oc8051_tc1_n164, oc8051_sfr1_oc8051_tc1_n163,
         oc8051_sfr1_oc8051_tc1_n162, oc8051_sfr1_oc8051_tc1_n161,
         oc8051_sfr1_oc8051_tc1_n160, oc8051_sfr1_oc8051_tc1_n159,
         oc8051_sfr1_oc8051_tc1_n158, oc8051_sfr1_oc8051_tc1_n157,
         oc8051_sfr1_oc8051_tc1_n156, oc8051_sfr1_oc8051_tc1_n155,
         oc8051_sfr1_oc8051_tc1_n154, oc8051_sfr1_oc8051_tc1_n153,
         oc8051_sfr1_oc8051_tc1_n152, oc8051_sfr1_oc8051_tc1_n151,
         oc8051_sfr1_oc8051_tc1_n150, oc8051_sfr1_oc8051_tc1_n149,
         oc8051_sfr1_oc8051_tc1_n148, oc8051_sfr1_oc8051_tc1_n147,
         oc8051_sfr1_oc8051_tc1_n146, oc8051_sfr1_oc8051_tc1_n145,
         oc8051_sfr1_oc8051_tc1_n144, oc8051_sfr1_oc8051_tc1_n143,
         oc8051_sfr1_oc8051_tc1_n142, oc8051_sfr1_oc8051_tc1_n141,
         oc8051_sfr1_oc8051_tc1_n140, oc8051_sfr1_oc8051_tc1_n139,
         oc8051_sfr1_oc8051_tc1_n138, oc8051_sfr1_oc8051_tc1_n137,
         oc8051_sfr1_oc8051_tc1_n136, oc8051_sfr1_oc8051_tc1_n135,
         oc8051_sfr1_oc8051_tc1_n134, oc8051_sfr1_oc8051_tc1_n133,
         oc8051_sfr1_oc8051_tc1_n132, oc8051_sfr1_oc8051_tc1_n131,
         oc8051_sfr1_oc8051_tc1_n130, oc8051_sfr1_oc8051_tc1_n129,
         oc8051_sfr1_oc8051_tc1_n128, oc8051_sfr1_oc8051_tc1_n127,
         oc8051_sfr1_oc8051_tc1_n126, oc8051_sfr1_oc8051_tc1_n125,
         oc8051_sfr1_oc8051_tc1_n124, oc8051_sfr1_oc8051_tc1_n123,
         oc8051_sfr1_oc8051_tc1_n122, oc8051_sfr1_oc8051_tc1_n121,
         oc8051_sfr1_oc8051_tc1_n120, oc8051_sfr1_oc8051_tc1_n119,
         oc8051_sfr1_oc8051_tc1_n118, oc8051_sfr1_oc8051_tc1_n117,
         oc8051_sfr1_oc8051_tc1_n116, oc8051_sfr1_oc8051_tc1_n115,
         oc8051_sfr1_oc8051_tc1_n114, oc8051_sfr1_oc8051_tc1_n113,
         oc8051_sfr1_oc8051_tc1_n112, oc8051_sfr1_oc8051_tc1_n111,
         oc8051_sfr1_oc8051_tc1_n110, oc8051_sfr1_oc8051_tc1_n109,
         oc8051_sfr1_oc8051_tc1_n108, oc8051_sfr1_oc8051_tc1_n107,
         oc8051_sfr1_oc8051_tc1_n106, oc8051_sfr1_oc8051_tc1_n105,
         oc8051_sfr1_oc8051_tc1_n104, oc8051_sfr1_oc8051_tc1_n103,
         oc8051_sfr1_oc8051_tc1_n102, oc8051_sfr1_oc8051_tc1_n101,
         oc8051_sfr1_oc8051_tc1_n100, oc8051_sfr1_oc8051_tc1_n99,
         oc8051_sfr1_oc8051_tc1_n98, oc8051_sfr1_oc8051_tc1_n97,
         oc8051_sfr1_oc8051_tc1_n96, oc8051_sfr1_oc8051_tc1_n95,
         oc8051_sfr1_oc8051_tc1_n94, oc8051_sfr1_oc8051_tc1_n93,
         oc8051_sfr1_oc8051_tc1_n92, oc8051_sfr1_oc8051_tc1_n91,
         oc8051_sfr1_oc8051_tc1_n90, oc8051_sfr1_oc8051_tc1_n89,
         oc8051_sfr1_oc8051_tc1_n88, oc8051_sfr1_oc8051_tc1_n87,
         oc8051_sfr1_oc8051_tc1_n86, oc8051_sfr1_oc8051_tc1_n85,
         oc8051_sfr1_oc8051_tc1_n84, oc8051_sfr1_oc8051_tc1_n83,
         oc8051_sfr1_oc8051_tc1_n82, oc8051_sfr1_oc8051_tc1_n81,
         oc8051_sfr1_oc8051_tc1_n80, oc8051_sfr1_oc8051_tc1_n79,
         oc8051_sfr1_oc8051_tc1_n78, oc8051_sfr1_oc8051_tc1_n77,
         oc8051_sfr1_oc8051_tc1_n76, oc8051_sfr1_oc8051_tc1_n75,
         oc8051_sfr1_oc8051_tc1_n74, oc8051_sfr1_oc8051_tc1_n73,
         oc8051_sfr1_oc8051_tc1_n72, oc8051_sfr1_oc8051_tc1_n71,
         oc8051_sfr1_oc8051_tc1_n70, oc8051_sfr1_oc8051_tc1_n69,
         oc8051_sfr1_oc8051_tc1_n68, oc8051_sfr1_oc8051_tc1_n67,
         oc8051_sfr1_oc8051_tc1_n66, oc8051_sfr1_oc8051_tc1_n65,
         oc8051_sfr1_oc8051_tc1_n64, oc8051_sfr1_oc8051_tc1_n63,
         oc8051_sfr1_oc8051_tc1_n62, oc8051_sfr1_oc8051_tc1_n61,
         oc8051_sfr1_oc8051_tc1_n60, oc8051_sfr1_oc8051_tc1_n59,
         oc8051_sfr1_oc8051_tc1_n58, oc8051_sfr1_oc8051_tc1_n57,
         oc8051_sfr1_oc8051_tc1_n56, oc8051_sfr1_oc8051_tc1_n55,
         oc8051_sfr1_oc8051_tc1_n54, oc8051_sfr1_oc8051_tc1_n53,
         oc8051_sfr1_oc8051_tc1_n52, oc8051_sfr1_oc8051_tc1_n51,
         oc8051_sfr1_oc8051_tc1_n50, oc8051_sfr1_oc8051_tc1_n49,
         oc8051_sfr1_oc8051_tc1_n48, oc8051_sfr1_oc8051_tc1_n47,
         oc8051_sfr1_oc8051_tc1_n46, oc8051_sfr1_oc8051_tc1_n45,
         oc8051_sfr1_oc8051_tc1_n44, oc8051_sfr1_oc8051_tc1_n43,
         oc8051_sfr1_oc8051_tc1_n42, oc8051_sfr1_oc8051_tc1_n41,
         oc8051_sfr1_oc8051_tc1_n40, oc8051_sfr1_oc8051_tc1_n39,
         oc8051_sfr1_oc8051_tc1_n38, oc8051_sfr1_oc8051_tc1_n37,
         oc8051_sfr1_oc8051_tc1_n36, oc8051_sfr1_oc8051_tc1_n35,
         oc8051_sfr1_oc8051_tc1_n34, oc8051_sfr1_oc8051_tc1_n33,
         oc8051_sfr1_oc8051_tc1_n32, oc8051_sfr1_oc8051_tc1_n31,
         oc8051_sfr1_oc8051_tc1_n30, oc8051_sfr1_oc8051_tc1_n29,
         oc8051_sfr1_oc8051_tc1_n28, oc8051_sfr1_oc8051_tc1_n27,
         oc8051_sfr1_oc8051_tc1_n26, oc8051_sfr1_oc8051_tc1_n25,
         oc8051_sfr1_oc8051_tc1_n24, oc8051_sfr1_oc8051_tc1_n23,
         oc8051_sfr1_oc8051_tc1_n22, oc8051_sfr1_oc8051_tc1_n21,
         oc8051_sfr1_oc8051_tc1_n20, oc8051_sfr1_oc8051_tc1_n19,
         oc8051_sfr1_oc8051_tc1_n18, oc8051_sfr1_oc8051_tc1_n17,
         oc8051_sfr1_oc8051_tc1_n16, oc8051_sfr1_oc8051_tc1_n15,
         oc8051_sfr1_oc8051_tc1_n14, oc8051_sfr1_oc8051_tc1_n13,
         oc8051_sfr1_oc8051_tc1_n12, oc8051_sfr1_oc8051_tc1_n11,
         oc8051_sfr1_oc8051_tc1_n10, oc8051_sfr1_oc8051_tc1_n9,
         oc8051_sfr1_oc8051_tc1_n8, oc8051_sfr1_oc8051_tc1_n7,
         oc8051_sfr1_oc8051_tc1_n6, oc8051_sfr1_oc8051_tc1_n4,
         oc8051_sfr1_oc8051_tc1_n3, oc8051_sfr1_oc8051_tc1_n2,
         oc8051_sfr1_oc8051_tc1_n1, oc8051_sfr1_oc8051_tc1_n268,
         oc8051_sfr1_oc8051_tc1_n267, oc8051_sfr1_oc8051_tc1_n266,
         oc8051_sfr1_oc8051_tc1_n265, oc8051_sfr1_oc8051_tc1_n264,
         oc8051_sfr1_oc8051_tc1_n263, oc8051_sfr1_oc8051_tc1_n262,
         oc8051_sfr1_oc8051_tc1_n261, oc8051_sfr1_oc8051_tc1_n260,
         oc8051_sfr1_oc8051_tc1_n259, oc8051_sfr1_oc8051_tc1_n258,
         oc8051_sfr1_oc8051_tc1_n257, oc8051_sfr1_oc8051_tc1_n256,
         oc8051_sfr1_oc8051_tc1_n255, oc8051_sfr1_oc8051_tc1_n254,
         oc8051_sfr1_oc8051_tc1_n253, oc8051_sfr1_oc8051_tc1_n252,
         oc8051_sfr1_oc8051_tc1_n251, oc8051_sfr1_oc8051_tc1_n250,
         oc8051_sfr1_oc8051_tc1_n249, oc8051_sfr1_oc8051_tc1_n248,
         oc8051_sfr1_oc8051_tc1_n247, oc8051_sfr1_oc8051_tc1_n246,
         oc8051_sfr1_oc8051_tc1_n245, oc8051_sfr1_oc8051_tc1_n244,
         oc8051_sfr1_oc8051_tc1_n243, oc8051_sfr1_oc8051_tc1_n242,
         oc8051_sfr1_oc8051_tc1_n241, oc8051_sfr1_oc8051_tc1_n240,
         oc8051_sfr1_oc8051_tc1_n239, oc8051_sfr1_oc8051_tc1_n238,
         oc8051_sfr1_oc8051_tc1_n237, oc8051_sfr1_oc8051_tc1_n236,
         oc8051_sfr1_oc8051_tc1_n235, oc8051_sfr1_oc8051_tc1_n234,
         oc8051_sfr1_oc8051_tc1_n233, oc8051_sfr1_oc8051_tc1_n232,
         oc8051_sfr1_oc8051_tc1_n231, oc8051_sfr1_oc8051_tc1_n230,
         oc8051_sfr1_oc8051_tc1_n229, oc8051_sfr1_oc8051_tc1_n228,
         oc8051_sfr1_oc8051_tc1_n227, oc8051_sfr1_oc8051_tc1_n226,
         oc8051_sfr1_oc8051_tc1_n225, oc8051_sfr1_oc8051_tc1_n224,
         oc8051_sfr1_oc8051_tc1_n223, oc8051_sfr1_oc8051_tc1_n222,
         oc8051_sfr1_oc8051_tc1_n221, oc8051_sfr1_oc8051_tc1_n220,
         oc8051_sfr1_oc8051_tc1_n219, oc8051_sfr1_oc8051_tc1_n218,
         oc8051_sfr1_oc8051_tc1_n217, oc8051_sfr1_oc8051_tc1_n216,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_15, oc8051_sfr1_oc8051_tc1_u3_u8_z_14,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_13, oc8051_sfr1_oc8051_tc1_u3_u8_z_12,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_11, oc8051_sfr1_oc8051_tc1_u3_u8_z_10,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_9, oc8051_sfr1_oc8051_tc1_u3_u8_z_8,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_7, oc8051_sfr1_oc8051_tc1_u3_u8_z_6,
         oc8051_sfr1_oc8051_tc1_u3_u8_z_5, oc8051_sfr1_oc8051_tc1_u3_u1_z_15,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_14, oc8051_sfr1_oc8051_tc1_u3_u1_z_13,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_12, oc8051_sfr1_oc8051_tc1_u3_u1_z_11,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_10, oc8051_sfr1_oc8051_tc1_u3_u1_z_9,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_8, oc8051_sfr1_oc8051_tc1_u3_u1_z_7,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_6, oc8051_sfr1_oc8051_tc1_u3_u1_z_5,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_4, oc8051_sfr1_oc8051_tc1_u3_u1_z_3,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_2, oc8051_sfr1_oc8051_tc1_u3_u1_z_1,
         oc8051_sfr1_oc8051_tc1_u3_u1_z_0, oc8051_sfr1_oc8051_tc1_n5,
         oc8051_sfr1_oc8051_tc1_n203, oc8051_sfr1_oc8051_tc1_n202,
         oc8051_sfr1_oc8051_tc1_n201, oc8051_sfr1_oc8051_tc1_n200,
         oc8051_sfr1_oc8051_tc1_n199, oc8051_sfr1_oc8051_tc1_n198,
         oc8051_sfr1_oc8051_tc1_n197, oc8051_sfr1_oc8051_tc1_n196,
         oc8051_sfr1_oc8051_tc1_n192, oc8051_sfr1_oc8051_tc1_n191,
         oc8051_sfr1_oc8051_tc1_n190, oc8051_sfr1_oc8051_tc1_n174,
         oc8051_sfr1_oc8051_tc1_n173, oc8051_sfr1_oc8051_tc1_n172,
         oc8051_sfr1_oc8051_tc1_n171, oc8051_sfr1_oc8051_tc1_n170,
         oc8051_sfr1_oc8051_tc1_n169, oc8051_sfr1_oc8051_tc1_n168,
         oc8051_sfr1_oc8051_tc1_n167, oc8051_sfr1_oc8051_tc1_n166,
         oc8051_sfr1_oc8051_tc1_n165, oc8051_sfr1_oc8051_tc1_n1640,
         oc8051_sfr1_oc8051_tc1_n1630, oc8051_sfr1_oc8051_tc1_n1620,
         oc8051_sfr1_oc8051_tc1_n1610, oc8051_sfr1_oc8051_tc1_n920,
         oc8051_sfr1_oc8051_tc1_n910, oc8051_sfr1_oc8051_tc1_n900,
         oc8051_sfr1_oc8051_tc1_n890, oc8051_sfr1_oc8051_tc1_n880,
         oc8051_sfr1_oc8051_tc1_n870, oc8051_sfr1_oc8051_tc1_n860,
         oc8051_sfr1_oc8051_tc1_n850, oc8051_sfr1_oc8051_tc1_n840,
         oc8051_sfr1_oc8051_tc1_n630, oc8051_sfr1_oc8051_tc1_n620,
         oc8051_sfr1_oc8051_tc1_n610, oc8051_sfr1_oc8051_tc1_n600,
         oc8051_sfr1_oc8051_tc1_n590, oc8051_sfr1_oc8051_tc1_n580,
         oc8051_sfr1_oc8051_tc1_n570, oc8051_sfr1_oc8051_tc1_n560,
         oc8051_sfr1_oc8051_tc1_n550, oc8051_sfr1_oc8051_tc1_n540,
         oc8051_sfr1_oc8051_tc1_n530, oc8051_sfr1_oc8051_tc1_n520,
         oc8051_sfr1_oc8051_tc1_n510, oc8051_sfr1_oc8051_tc1_n500,
         oc8051_sfr1_oc8051_tc1_n490, oc8051_sfr1_oc8051_tc1_n480,
         oc8051_sfr1_oc8051_tc1_n470, oc8051_sfr1_oc8051_tc1_t1_buff,
         oc8051_sfr1_oc8051_tc1_t0_buff, oc8051_sfr1_oc8051_tc21_n139,
         oc8051_sfr1_oc8051_tc21_n138, oc8051_sfr1_oc8051_tc21_n137,
         oc8051_sfr1_oc8051_tc21_n136, oc8051_sfr1_oc8051_tc21_n135,
         oc8051_sfr1_oc8051_tc21_n134, oc8051_sfr1_oc8051_tc21_n133,
         oc8051_sfr1_oc8051_tc21_n132, oc8051_sfr1_oc8051_tc21_n131,
         oc8051_sfr1_oc8051_tc21_n130, oc8051_sfr1_oc8051_tc21_n129,
         oc8051_sfr1_oc8051_tc21_n128, oc8051_sfr1_oc8051_tc21_n127,
         oc8051_sfr1_oc8051_tc21_n126, oc8051_sfr1_oc8051_tc21_n125,
         oc8051_sfr1_oc8051_tc21_n124, oc8051_sfr1_oc8051_tc21_n123,
         oc8051_sfr1_oc8051_tc21_n122, oc8051_sfr1_oc8051_tc21_n121,
         oc8051_sfr1_oc8051_tc21_n120, oc8051_sfr1_oc8051_tc21_n119,
         oc8051_sfr1_oc8051_tc21_n118, oc8051_sfr1_oc8051_tc21_n117,
         oc8051_sfr1_oc8051_tc21_n116, oc8051_sfr1_oc8051_tc21_n115,
         oc8051_sfr1_oc8051_tc21_n114, oc8051_sfr1_oc8051_tc21_n113,
         oc8051_sfr1_oc8051_tc21_n112, oc8051_sfr1_oc8051_tc21_n111,
         oc8051_sfr1_oc8051_tc21_n110, oc8051_sfr1_oc8051_tc21_n109,
         oc8051_sfr1_oc8051_tc21_n108, oc8051_sfr1_oc8051_tc21_n107,
         oc8051_sfr1_oc8051_tc21_n106, oc8051_sfr1_oc8051_tc21_n105,
         oc8051_sfr1_oc8051_tc21_n104, oc8051_sfr1_oc8051_tc21_n103,
         oc8051_sfr1_oc8051_tc21_n102, oc8051_sfr1_oc8051_tc21_n101,
         oc8051_sfr1_oc8051_tc21_n100, oc8051_sfr1_oc8051_tc21_n99,
         oc8051_sfr1_oc8051_tc21_n98, oc8051_sfr1_oc8051_tc21_n97,
         oc8051_sfr1_oc8051_tc21_n96, oc8051_sfr1_oc8051_tc21_n95,
         oc8051_sfr1_oc8051_tc21_n94, oc8051_sfr1_oc8051_tc21_n93,
         oc8051_sfr1_oc8051_tc21_n92, oc8051_sfr1_oc8051_tc21_n91,
         oc8051_sfr1_oc8051_tc21_n90, oc8051_sfr1_oc8051_tc21_n89,
         oc8051_sfr1_oc8051_tc21_n88, oc8051_sfr1_oc8051_tc21_n87,
         oc8051_sfr1_oc8051_tc21_n86, oc8051_sfr1_oc8051_tc21_n85,
         oc8051_sfr1_oc8051_tc21_n84, oc8051_sfr1_oc8051_tc21_n83,
         oc8051_sfr1_oc8051_tc21_n82, oc8051_sfr1_oc8051_tc21_n81,
         oc8051_sfr1_oc8051_tc21_n80, oc8051_sfr1_oc8051_tc21_n79,
         oc8051_sfr1_oc8051_tc21_n78, oc8051_sfr1_oc8051_tc21_n77,
         oc8051_sfr1_oc8051_tc21_n76, oc8051_sfr1_oc8051_tc21_n75,
         oc8051_sfr1_oc8051_tc21_n74, oc8051_sfr1_oc8051_tc21_n73,
         oc8051_sfr1_oc8051_tc21_n72, oc8051_sfr1_oc8051_tc21_n71,
         oc8051_sfr1_oc8051_tc21_n70, oc8051_sfr1_oc8051_tc21_n69,
         oc8051_sfr1_oc8051_tc21_n68, oc8051_sfr1_oc8051_tc21_n67,
         oc8051_sfr1_oc8051_tc21_n66, oc8051_sfr1_oc8051_tc21_n65,
         oc8051_sfr1_oc8051_tc21_n64, oc8051_sfr1_oc8051_tc21_n63,
         oc8051_sfr1_oc8051_tc21_n62, oc8051_sfr1_oc8051_tc21_n61,
         oc8051_sfr1_oc8051_tc21_n60, oc8051_sfr1_oc8051_tc21_n59,
         oc8051_sfr1_oc8051_tc21_n58, oc8051_sfr1_oc8051_tc21_n57,
         oc8051_sfr1_oc8051_tc21_n56, oc8051_sfr1_oc8051_tc21_n55,
         oc8051_sfr1_oc8051_tc21_n54, oc8051_sfr1_oc8051_tc21_n53,
         oc8051_sfr1_oc8051_tc21_n52, oc8051_sfr1_oc8051_tc21_n51,
         oc8051_sfr1_oc8051_tc21_n50, oc8051_sfr1_oc8051_tc21_n49,
         oc8051_sfr1_oc8051_tc21_n48, oc8051_sfr1_oc8051_tc21_n47,
         oc8051_sfr1_oc8051_tc21_n46, oc8051_sfr1_oc8051_tc21_n45,
         oc8051_sfr1_oc8051_tc21_n44, oc8051_sfr1_oc8051_tc21_n43,
         oc8051_sfr1_oc8051_tc21_n42, oc8051_sfr1_oc8051_tc21_n41,
         oc8051_sfr1_oc8051_tc21_n40, oc8051_sfr1_oc8051_tc21_n39,
         oc8051_sfr1_oc8051_tc21_n38, oc8051_sfr1_oc8051_tc21_n37,
         oc8051_sfr1_oc8051_tc21_n36, oc8051_sfr1_oc8051_tc21_n35,
         oc8051_sfr1_oc8051_tc21_n34, oc8051_sfr1_oc8051_tc21_n33,
         oc8051_sfr1_oc8051_tc21_n32, oc8051_sfr1_oc8051_tc21_n31,
         oc8051_sfr1_oc8051_tc21_n30, oc8051_sfr1_oc8051_tc21_n29,
         oc8051_sfr1_oc8051_tc21_n28, oc8051_sfr1_oc8051_tc21_n27,
         oc8051_sfr1_oc8051_tc21_n26, oc8051_sfr1_oc8051_tc21_n25,
         oc8051_sfr1_oc8051_tc21_n24, oc8051_sfr1_oc8051_tc21_n23,
         oc8051_sfr1_oc8051_tc21_n22, oc8051_sfr1_oc8051_tc21_n21,
         oc8051_sfr1_oc8051_tc21_n20, oc8051_sfr1_oc8051_tc21_n19,
         oc8051_sfr1_oc8051_tc21_n18, oc8051_sfr1_oc8051_tc21_n17,
         oc8051_sfr1_oc8051_tc21_n16, oc8051_sfr1_oc8051_tc21_n15,
         oc8051_sfr1_oc8051_tc21_n14, oc8051_sfr1_oc8051_tc21_n13,
         oc8051_sfr1_oc8051_tc21_n12, oc8051_sfr1_oc8051_tc21_n11,
         oc8051_sfr1_oc8051_tc21_n10, oc8051_sfr1_oc8051_tc21_n9,
         oc8051_sfr1_oc8051_tc21_n4, oc8051_sfr1_oc8051_tc21_n3,
         oc8051_sfr1_oc8051_tc21_n2, oc8051_sfr1_oc8051_tc21_n191,
         oc8051_sfr1_oc8051_tc21_n190, oc8051_sfr1_oc8051_tc21_n189,
         oc8051_sfr1_oc8051_tc21_n188, oc8051_sfr1_oc8051_tc21_n187,
         oc8051_sfr1_oc8051_tc21_n186, oc8051_sfr1_oc8051_tc21_n185,
         oc8051_sfr1_oc8051_tc21_n184, oc8051_sfr1_oc8051_tc21_n183,
         oc8051_sfr1_oc8051_tc21_n182, oc8051_sfr1_oc8051_tc21_n181,
         oc8051_sfr1_oc8051_tc21_n180, oc8051_sfr1_oc8051_tc21_n179,
         oc8051_sfr1_oc8051_tc21_n178, oc8051_sfr1_oc8051_tc21_n177,
         oc8051_sfr1_oc8051_tc21_n176, oc8051_sfr1_oc8051_tc21_n175,
         oc8051_sfr1_oc8051_tc21_n174, oc8051_sfr1_oc8051_tc21_n173,
         oc8051_sfr1_oc8051_tc21_n172, oc8051_sfr1_oc8051_tc21_n171,
         oc8051_sfr1_oc8051_tc21_n170, oc8051_sfr1_oc8051_tc21_n169,
         oc8051_sfr1_oc8051_tc21_n168, oc8051_sfr1_oc8051_tc21_n167,
         oc8051_sfr1_oc8051_tc21_n166, oc8051_sfr1_oc8051_tc21_n165,
         oc8051_sfr1_oc8051_tc21_n164, oc8051_sfr1_oc8051_tc21_n163,
         oc8051_sfr1_oc8051_tc21_n162, oc8051_sfr1_oc8051_tc21_n161,
         oc8051_sfr1_oc8051_tc21_n160, oc8051_sfr1_oc8051_tc21_n159,
         oc8051_sfr1_oc8051_tc21_n158, oc8051_sfr1_oc8051_tc21_n157,
         oc8051_sfr1_oc8051_tc21_n156, oc8051_sfr1_oc8051_tc21_n155,
         oc8051_sfr1_oc8051_tc21_n154, oc8051_sfr1_oc8051_tc21_n153,
         oc8051_sfr1_oc8051_tc21_n152, oc8051_sfr1_oc8051_tc21_n151,
         oc8051_sfr1_oc8051_tc21_n150, oc8051_sfr1_oc8051_tc21_n8,
         oc8051_sfr1_oc8051_tc21_n7, oc8051_sfr1_oc8051_tc21_n6,
         oc8051_sfr1_oc8051_tc21_n5, oc8051_sfr1_oc8051_tc21_n1,
         oc8051_sfr1_oc8051_tc21_n220, oc8051_sfr1_oc8051_tc21_t2_r,
         oc8051_sfr1_oc8051_tc21_n217, oc8051_sfr1_oc8051_tc21_t2ex_r,
         oc8051_sfr1_oc8051_tc21_n850, oc8051_sfr1_oc8051_tc21_n840,
         oc8051_sfr1_oc8051_tc21_n830, oc8051_sfr1_oc8051_tc21_n820,
         oc8051_sfr1_oc8051_tc21_n810, oc8051_sfr1_oc8051_tc21_n800,
         oc8051_sfr1_oc8051_tc21_n790, oc8051_sfr1_oc8051_tc21_n780,
         oc8051_sfr1_oc8051_tc21_n770, oc8051_sfr1_oc8051_tc21_n760,
         oc8051_sfr1_oc8051_tc21_n750, oc8051_sfr1_oc8051_tc21_n740,
         oc8051_sfr1_oc8051_tc21_n730, oc8051_sfr1_oc8051_tc21_n720,
         oc8051_sfr1_oc8051_tc21_n710, oc8051_sfr1_oc8051_tc21_n700,
         oc8051_sfr1_oc8051_tc21_n690, oc8051_sfr1_oc8051_tc21_tc2_event,
         oc8051_sfr1_oc8051_tc21_neg_trans, oc8051_sfr1_oc8051_tc21_tf2_set;
  wire   [7:0] op1_n;
  wire   [2:0] op1_cur;
  wire   [2:0] ram_rd_sel;
  wire   [2:0] ram_wr_sel;
  wire   [2:0] src_sel1;
  wire   [1:0] src_sel2;
  wire   [3:0] alu_op;
  wire   [1:0] psw_set;
  wire   [1:0] cy_sel;
  wire   [2:0] pc_wr_sel;
  wire   [1:0] comp_sel;
  wire   [1:0] wr_sfr;
  wire   [2:0] mem_act;
  wire   [7:0] src1;
  wire   [7:0] src2;
  wire   [7:0] src3;
  wire   [7:0] des_acc;
  wire   [7:0] sub_result;
  wire   [7:0] des2;
  wire   [7:0] rd_addr;
  wire   [7:0] ram_data;
  wire   [7:0] wr_addr;
  wire   [7:0] wr_dat;
  wire   [7:0] acc;
  wire   [7:0] ram_out;
  wire   [15:0] pc;
  wire   [7:0] op2_n;
  wire   [7:0] op3_n;
  wire   [7:0] dptr_hi;
  wire   [7:0] dptr_lo;
  wire   [7:0] ri;
  wire   [1:0] bank_sel;
  wire   [7:0] sfr_out;
  wire   [5:0] int_src;
  wire   [7:0] sp_w;
  wire   [7:0] sp;
  wire   [2:0] oc8051_decoder1_ram_rd_sel_r;
  wire   [7:0] oc8051_decoder1_op;
  wire   [7:0] oc8051_alu1_des_acc_1;
  wire   [15:0] oc8051_alu1_dec;
  wire   [15:0] oc8051_alu1_inc;
  wire   [7:0] oc8051_alu1_divsrc2;
  wire   [7:0] oc8051_alu1_divsrc1;
  wire   [7:0] oc8051_alu1_mulsrc2;
  wire   [7:0] oc8051_alu1_mulsrc1;
  wire   [8:0] oc8051_alu1_oc8051_div1_sub0;
  wire   [8:0] oc8051_alu1_oc8051_div1_sub1;
  wire   [7:0] oc8051_alu1_oc8051_div1_tmp_rem;
  wire   [8:2] oc8051_alu1_oc8051_div1_sub_98_carry;
  wire   [8:3] oc8051_alu1_oc8051_div1_sub_94_carry;
  wire   [15:2] oc8051_alu1_add_204_carry;
  wire   [7:0] oc8051_ram_top1_wr_data_m;
  wire   [7:0] oc8051_ram_top1_rd_data_m;
  wire   [7:0] oc8051_ram_top1_wr_data_r;
  wire   [7:0] oc8051_alu_src_sel1_op3_r;
  wire   [7:0] oc8051_alu_src_sel1_op1_r;
  wire   [7:0] oc8051_memory_interface1_op2_buff;
  wire   [7:0] oc8051_memory_interface1_op3_buff;
  wire   [7:0] oc8051_memory_interface1_op3;
  wire   [7:0] oc8051_memory_interface1_op2;
  wire   [7:0] oc8051_memory_interface1_imm2_r;
  wire   [7:0] oc8051_memory_interface1_imm_r;
  wire   [7:0] oc8051_memory_interface1_ri_r;
  wire   [4:0] oc8051_memory_interface1_rn_r;
  wire   [7:0] oc8051_sfr1_rcap2h;
  wire   [7:0] oc8051_sfr1_rcap2l;
  wire   [7:0] oc8051_sfr1_th2;
  wire   [7:0] oc8051_sfr1_tl2;
  wire   [7:0] oc8051_sfr1_th1;
  wire   [7:0] oc8051_sfr1_tl1;
  wire   [7:0] oc8051_sfr1_th0;
  wire   [7:0] oc8051_sfr1_tl0;
  wire   [7:0] oc8051_sfr1_tmod;
  wire   [7:0] oc8051_sfr1_sbuf;
  wire   [7:0] oc8051_sfr1_pcon;
  wire   [7:2] oc8051_sfr1_oc8051_sp1_add_102_s2_carry;
  wire   [15:2] oc8051_sfr1_oc8051_tc1_r372_carry;
  wire   [7:2] oc8051_sfr1_oc8051_tc1_add_220_carry;
  wire   [7:2] oc8051_sfr1_oc8051_tc1_r364_carry;
  wire   [15:2] oc8051_sfr1_oc8051_tc1_r360_carry;
  wire   [15:2] oc8051_sfr1_oc8051_tc21_r320_carry;
  assign wbd_stb_o = wbd_cyc_o;
  assign wbi_stb_o = wbi_cyc_o;

  TIELO_X1M_A12TS u6 ( .Y(n2) );
  TIEHI_X1M_A12TS u7 ( .Y(wbi_cyc_o) );
  NOR2_X0P5A_A12TS u8 ( .A(wr_ind), .B(n3), .Y(n_5_net_) );
  AND2_X0P5M_A12TS u9 ( .A(pc_wr), .B(comp_wait), .Y(n_3_net_) );
  AOI2XB1_X0P5M_A12TS u10 ( .A1N(wr_ind), .A0(wr_addr[7]), .B0(n3), .Y(
        n_0_net_) );
  INV_X0P5B_A12TS u11 ( .A(wr_o), .Y(n3) );
  INV_X0P5B_A12TS oc8051_decoder1_u472 ( .A(oc8051_decoder1_state_1_), .Y(
        oc8051_decoder1_n317) );
  INV_X0P5B_A12TS oc8051_decoder1_u471 ( .A(oc8051_decoder1_state_0_), .Y(
        oc8051_decoder1_n316) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u470 ( .A(oc8051_decoder1_n317), .B(
        oc8051_decoder1_n316), .Y(oc8051_decoder1_n303) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u469 ( .A(oc8051_decoder1_n303), .B(
        wait_data), .Y(rd) );
  INV_X0P5B_A12TS oc8051_decoder1_u468 ( .A(mem_wait), .Y(oc8051_decoder1_n435) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u467 ( .A(rd), .B(oc8051_decoder1_n435), 
        .Y(oc8051_decoder1_n318) );
  INV_X0P5B_A12TS oc8051_decoder1_u466 ( .A(op1_n[0]), .Y(oc8051_decoder1_n301) );
  OR2_X0P5M_A12TS oc8051_decoder1_u465 ( .A(rd), .B(mem_wait), .Y(
        oc8051_decoder1_n439) );
  INV_X0P5B_A12TS oc8051_decoder1_u464 ( .A(oc8051_decoder1_op[0]), .Y(
        oc8051_decoder1_n302) );
  INV_X0P5B_A12TS oc8051_decoder1_u463 ( .A(op1_n[1]), .Y(oc8051_decoder1_n304) );
  INV_X0P5B_A12TS oc8051_decoder1_u462 ( .A(oc8051_decoder1_op[1]), .Y(
        oc8051_decoder1_n305) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u461 ( .A0(oc8051_decoder1_n318), .A1(
        oc8051_decoder1_n304), .B0(oc8051_decoder1_n439), .B1(
        oc8051_decoder1_n305), .Y(op1_cur[1]) );
  INV_X0P5B_A12TS oc8051_decoder1_u460 ( .A(op1_cur[1]), .Y(
        oc8051_decoder1_n22) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u459 ( .A(op1_cur[0]), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n25) );
  INV_X0P5B_A12TS oc8051_decoder1_u458 ( .A(oc8051_decoder1_op[3]), .Y(
        oc8051_decoder1_n309) );
  INV_X0P5B_A12TS oc8051_decoder1_u457 ( .A(op1_n[3]), .Y(oc8051_decoder1_n308) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u456 ( .A(oc8051_decoder1_n309), .B(
        oc8051_decoder1_n308), .S0(rd), .Y(oc8051_decoder1_n440) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u455 ( .A(oc8051_decoder1_n440), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n69) );
  INV_X0P5B_A12TS oc8051_decoder1_u454 ( .A(op1_n[2]), .Y(oc8051_decoder1_n306) );
  INV_X0P5B_A12TS oc8051_decoder1_u453 ( .A(oc8051_decoder1_op[2]), .Y(
        oc8051_decoder1_n307) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u452 ( .A0(oc8051_decoder1_n318), .A1(
        oc8051_decoder1_n306), .B0(oc8051_decoder1_n439), .B1(
        oc8051_decoder1_n307), .Y(op1_cur[2]) );
  INV_X0P5B_A12TS oc8051_decoder1_u451 ( .A(op1_cur[2]), .Y(
        oc8051_decoder1_n131) );
  INV_X0P5B_A12TS oc8051_decoder1_u450 ( .A(oc8051_decoder1_op[7]), .Y(
        oc8051_decoder1_n315) );
  INV_X0P5B_A12TS oc8051_decoder1_u449 ( .A(op1_n[7]), .Y(oc8051_decoder1_n314) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u448 ( .A(oc8051_decoder1_n315), .B(
        oc8051_decoder1_n314), .S0(rd), .Y(oc8051_decoder1_n438) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u447 ( .A(oc8051_decoder1_n438), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n185) );
  INV_X0P5B_A12TS oc8051_decoder1_u446 ( .A(oc8051_decoder1_n185), .Y(
        oc8051_decoder1_n54) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u445 ( .A(oc8051_decoder1_n69), .B(
        oc8051_decoder1_n131), .C(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n334) );
  INV_X0P5B_A12TS oc8051_decoder1_u444 ( .A(oc8051_decoder1_n334), .Y(
        oc8051_decoder1_n224) );
  AND3_X0P5M_A12TS oc8051_decoder1_u443 ( .A(rd), .B(oc8051_decoder1_n25), .C(
        oc8051_decoder1_n224), .Y(oc8051_decoder1_n432) );
  INV_X0P5B_A12TS oc8051_decoder1_u442 ( .A(oc8051_decoder1_op[4]), .Y(
        oc8051_decoder1_n310) );
  INV_X0P5B_A12TS oc8051_decoder1_u441 ( .A(op1_n[4]), .Y(oc8051_decoder1_n300) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u440 ( .A(oc8051_decoder1_n310), .B(
        oc8051_decoder1_n300), .S0(rd), .Y(oc8051_decoder1_n437) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u439 ( .A(oc8051_decoder1_n437), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n82) );
  INV_X0P5B_A12TS oc8051_decoder1_u438 ( .A(oc8051_decoder1_n82), .Y(
        oc8051_decoder1_n165) );
  INV_X0P5B_A12TS oc8051_decoder1_u437 ( .A(oc8051_decoder1_op[5]), .Y(
        oc8051_decoder1_n312) );
  INV_X0P5B_A12TS oc8051_decoder1_u436 ( .A(op1_n[5]), .Y(oc8051_decoder1_n311) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u435 ( .A(oc8051_decoder1_n312), .B(
        oc8051_decoder1_n311), .S0(rd), .Y(oc8051_decoder1_n436) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u434 ( .A(oc8051_decoder1_n436), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n71) );
  INV_X0P5B_A12TS oc8051_decoder1_u433 ( .A(oc8051_decoder1_n71), .Y(
        oc8051_decoder1_n161) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u432 ( .A(oc8051_decoder1_n165), .B(
        oc8051_decoder1_n161), .Y(oc8051_decoder1_n59) );
  INV_X0P5B_A12TS oc8051_decoder1_u431 ( .A(op1_cur[0]), .Y(
        oc8051_decoder1_n137) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u430 ( .A(oc8051_decoder1_n71), .B(
        oc8051_decoder1_n137), .Y(oc8051_decoder1_n55) );
  INV_X0P5B_A12TS oc8051_decoder1_u429 ( .A(oc8051_decoder1_op[6]), .Y(
        oc8051_decoder1_n313) );
  INV_X0P5B_A12TS oc8051_decoder1_u428 ( .A(op1_n[6]), .Y(oc8051_decoder1_n299) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u427 ( .A(oc8051_decoder1_n313), .B(
        oc8051_decoder1_n299), .S0(rd), .Y(oc8051_decoder1_n434) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u426 ( .A(oc8051_decoder1_n434), .B(
        oc8051_decoder1_n435), .Y(oc8051_decoder1_n21) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u425 ( .A(oc8051_decoder1_n21), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n431) );
  INV_X0P5B_A12TS oc8051_decoder1_u424 ( .A(oc8051_decoder1_n21), .Y(
        oc8051_decoder1_n14) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u423 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n275) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u422 ( .A(oc8051_decoder1_n431), .B(
        oc8051_decoder1_n275), .Y(oc8051_decoder1_n141) );
  INV_X0P5B_A12TS oc8051_decoder1_u421 ( .A(oc8051_decoder1_n141), .Y(
        oc8051_decoder1_n118) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u420 ( .A(oc8051_decoder1_n432), .B(
        oc8051_decoder1_n59), .C(oc8051_decoder1_n55), .D(oc8051_decoder1_n118), .Y(oc8051_decoder1_n1804) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u419 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n225) );
  INV_X0P5B_A12TS oc8051_decoder1_u418 ( .A(oc8051_decoder1_n225), .Y(
        oc8051_decoder1_n139) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u417 ( .A0(oc8051_decoder1_n21), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n139), .Y(
        oc8051_decoder1_n433) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u416 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n432), .C0(
        oc8051_decoder1_n433), .Y(oc8051_decoder1_n1805) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u415 ( .A(oc8051_decoder1_n431), .B(
        oc8051_decoder1_n432), .Y(oc8051_decoder1_n1806) );
  INV_X0P5B_A12TS oc8051_decoder1_u414 ( .A(oc8051_decoder1_alu_op_0_), .Y(
        oc8051_decoder1_n124) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u413 ( .A(wait_data), .B(
        oc8051_decoder1_n124), .Y(alu_op[0]) );
  INV_X0P5B_A12TS oc8051_decoder1_u412 ( .A(oc8051_decoder1_alu_op_1_), .Y(
        oc8051_decoder1_n145) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u411 ( .A(wait_data), .B(
        oc8051_decoder1_n145), .Y(alu_op[1]) );
  NOR2B_X0P5M_A12TS oc8051_decoder1_u410 ( .AN(oc8051_decoder1_alu_op_2_), .B(
        wait_data), .Y(alu_op[2]) );
  INV_X0P5B_A12TS oc8051_decoder1_u409 ( .A(oc8051_decoder1_alu_op_3_), .Y(
        oc8051_decoder1_n379) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u408 ( .A(wait_data), .B(
        oc8051_decoder1_n379), .Y(alu_op[3]) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u407 ( .A(op1_cur[1]), .B(
        oc8051_decoder1_n137), .Y(oc8051_decoder1_n193) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u406 ( .A(oc8051_decoder1_n71), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n375) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u405 ( .A(oc8051_decoder1_n375), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n52) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u404 ( .A0(oc8051_decoder1_n161), .A1(
        oc8051_decoder1_n193), .B0(oc8051_decoder1_n52), .Y(
        oc8051_decoder1_n430) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u403 ( .A(op1_cur[1]), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n66) );
  INV_X0P5B_A12TS oc8051_decoder1_u402 ( .A(oc8051_decoder1_n66), .Y(
        oc8051_decoder1_n425) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u401 ( .A(oc8051_decoder1_n69), .B(
        oc8051_decoder1_n131), .Y(oc8051_decoder1_n36) );
  INV_X0P5B_A12TS oc8051_decoder1_u400 ( .A(oc8051_decoder1_n36), .Y(
        oc8051_decoder1_n90) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u399 ( .A(oc8051_decoder1_n425), .B(
        oc8051_decoder1_n90), .Y(oc8051_decoder1_n257) );
  INV_X0P5B_A12TS oc8051_decoder1_u398 ( .A(oc8051_decoder1_n257), .Y(
        oc8051_decoder1_n75) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u397 ( .A(oc8051_decoder1_n75), .B(
        oc8051_decoder1_n137), .Y(oc8051_decoder1_n270) );
  INV_X0P5B_A12TS oc8051_decoder1_u396 ( .A(oc8051_decoder1_n270), .Y(
        oc8051_decoder1_n109) );
  INV_X0P5B_A12TS oc8051_decoder1_u395 ( .A(oc8051_decoder1_n59), .Y(
        oc8051_decoder1_n53) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u394 ( .A(oc8051_decoder1_n53), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n283) );
  INV_X0P5B_A12TS oc8051_decoder1_u393 ( .A(oc8051_decoder1_n283), .Y(
        oc8051_decoder1_n221) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u392 ( .A0(oc8051_decoder1_n224), .A1(
        oc8051_decoder1_n430), .B0(oc8051_decoder1_n109), .B1(
        oc8051_decoder1_n221), .Y(oc8051_decoder1_n428) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u391 ( .A(oc8051_decoder1_n53), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n115) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u390 ( .A(oc8051_decoder1_n137), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n50) );
  INV_X0P5B_A12TS oc8051_decoder1_u389 ( .A(oc8051_decoder1_n50), .Y(
        oc8051_decoder1_n178) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u388 ( .A(oc8051_decoder1_n90), .B(
        oc8051_decoder1_n185), .C(oc8051_decoder1_n178), .Y(
        oc8051_decoder1_n322) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u387 ( .A(oc8051_decoder1_n115), .B(
        oc8051_decoder1_n322), .Y(oc8051_decoder1_n85) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u386 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n58) );
  INV_X0P5B_A12TS oc8051_decoder1_u385 ( .A(oc8051_decoder1_n58), .Y(
        oc8051_decoder1_n42) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u384 ( .A(oc8051_decoder1_n42), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n236) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u383 ( .A(oc8051_decoder1_n236), .B(
        oc8051_decoder1_n322), .Y(oc8051_decoder1_n84) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u382 ( .A(oc8051_decoder1_n85), .B(
        oc8051_decoder1_n84), .Y(oc8051_decoder1_n92) );
  INV_X0P5B_A12TS oc8051_decoder1_u381 ( .A(oc8051_decoder1_n92), .Y(
        oc8051_decoder1_n117) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u380 ( .A(oc8051_decoder1_n165), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n265) );
  INV_X0P5B_A12TS oc8051_decoder1_u379 ( .A(oc8051_decoder1_n265), .Y(
        oc8051_decoder1_n156) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u378 ( .A(oc8051_decoder1_n156), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n226) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u377 ( .A(oc8051_decoder1_n226), .B(
        oc8051_decoder1_n322), .Y(oc8051_decoder1_n83) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u376 ( .A(oc8051_decoder1_n117), .B(
        oc8051_decoder1_n83), .Y(oc8051_decoder1_n112) );
  INV_X0P5B_A12TS oc8051_decoder1_u375 ( .A(wait_data), .Y(
        oc8051_decoder1_n125) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u374 ( .A(oc8051_decoder1_n125), .B(
        oc8051_decoder1_n303), .Y(oc8051_decoder1_n33) );
  INV_X0P5B_A12TS oc8051_decoder1_u373 ( .A(oc8051_decoder1_n33), .Y(
        oc8051_decoder1_n5) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u372 ( .A(oc8051_decoder1_n316), .B(
        oc8051_decoder1_n125), .C(oc8051_decoder1_state_1_), .Y(
        oc8051_decoder1_n30) );
  INV_X0P5B_A12TS oc8051_decoder1_u371 ( .A(oc8051_decoder1_n30), .Y(
        oc8051_decoder1_n111) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u370 ( .A0(oc8051_decoder1_n85), .A1(
        oc8051_decoder1_n83), .B0(oc8051_decoder1_n111), .Y(
        oc8051_decoder1_n429) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u369 ( .A0(oc8051_decoder1_n428), .A1(
        oc8051_decoder1_n112), .B0(oc8051_decoder1_n5), .C0(
        oc8051_decoder1_n429), .Y(bit_addr_o) );
  INV_X0P5B_A12TS oc8051_decoder1_u368 ( .A(oc8051_decoder1_n322), .Y(
        oc8051_decoder1_n427) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u367 ( .A(oc8051_decoder1_n427), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n29) );
  INV_X0P5B_A12TS oc8051_decoder1_u366 ( .A(oc8051_decoder1_n29), .Y(
        oc8051_decoder1_n81) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u365 ( .A(oc8051_decoder1_n111), .B(
        oc8051_decoder1_n81), .Y(comp_sel[0]) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u364 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n156), .Y(oc8051_decoder1_n11) );
  INV_X0P5B_A12TS oc8051_decoder1_u363 ( .A(oc8051_decoder1_n11), .Y(
        oc8051_decoder1_n61) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u362 ( .A(oc8051_decoder1_n427), .B(
        oc8051_decoder1_n61), .Y(oc8051_decoder1_n99) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u361 ( .A(oc8051_decoder1_n111), .B(
        oc8051_decoder1_n33), .Y(oc8051_decoder1_n426) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u360 ( .A(oc8051_decoder1_n71), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n105) );
  OAI222_X0P5M_A12TS oc8051_decoder1_u359 ( .A0(oc8051_decoder1_n30), .A1(
        oc8051_decoder1_n99), .B0(oc8051_decoder1_n112), .B1(
        oc8051_decoder1_n426), .C0(comp_sel[0]), .C1(oc8051_decoder1_n105), 
        .Y(comp_sel[1]) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u358 ( .A(oc8051_decoder1_n317), .B(
        oc8051_decoder1_n125), .C(oc8051_decoder1_state_0_), .Y(
        oc8051_decoder1_n277) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u357 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n132) );
  INV_X0P5B_A12TS oc8051_decoder1_u356 ( .A(oc8051_decoder1_n132), .Y(
        oc8051_decoder1_n281) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u355 ( .A(op1_cur[0]), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n23) );
  INV_X0P5B_A12TS oc8051_decoder1_u354 ( .A(oc8051_decoder1_n23), .Y(
        oc8051_decoder1_n244) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u353 ( .A(oc8051_decoder1_n54), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n155) );
  INV_X0P5B_A12TS oc8051_decoder1_u352 ( .A(oc8051_decoder1_n155), .Y(
        oc8051_decoder1_n40) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u351 ( .A(oc8051_decoder1_n21), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n48) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u350 ( .A(oc8051_decoder1_n132), .B(
        oc8051_decoder1_n48), .Y(oc8051_decoder1_n164) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u349 ( .A0(oc8051_decoder1_n105), .A1(
        oc8051_decoder1_n22), .A2(oc8051_decoder1_n164), .B0(
        oc8051_decoder1_n425), .B1(oc8051_decoder1_n137), .Y(
        oc8051_decoder1_n411) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u348 ( .A(oc8051_decoder1_n221), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n104) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u347 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n411), .B0(oc8051_decoder1_n25), .C0(
        oc8051_decoder1_n104), .Y(oc8051_decoder1_n410) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u346 ( .A0(oc8051_decoder1_n281), .A1(
        oc8051_decoder1_n161), .B0(oc8051_decoder1_n244), .B1(
        oc8051_decoder1_n40), .C0(oc8051_decoder1_n410), .Y(
        oc8051_decoder1_n386) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u345 ( .A0(oc8051_decoder1_n156), .A1(
        oc8051_decoder1_n50), .B0(oc8051_decoder1_n59), .Y(oc8051_decoder1_n24) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u344 ( .A(op1_cur[2]), .B(
        oc8051_decoder1_n69), .Y(oc8051_decoder1_n26) );
  INV_X0P5B_A12TS oc8051_decoder1_u343 ( .A(oc8051_decoder1_n26), .Y(
        oc8051_decoder1_n67) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u342 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n24), .A2(oc8051_decoder1_n67), .B0(
        oc8051_decoder1_state_1_), .Y(oc8051_decoder1_n387) );
  INV_X0P5B_A12TS oc8051_decoder1_u341 ( .A(oc8051_decoder1_n69), .Y(
        oc8051_decoder1_n9) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u340 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n265), .Y(oc8051_decoder1_n186) );
  INV_X0P5B_A12TS oc8051_decoder1_u339 ( .A(oc8051_decoder1_n186), .Y(
        oc8051_decoder1_n373) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u338 ( .A0(oc8051_decoder1_n59), .A1(
        oc8051_decoder1_n21), .B0(oc8051_decoder1_n373), .Y(
        oc8051_decoder1_n409) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u337 ( .A(oc8051_decoder1_n61), .B(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n98) );
  INV_X0P5B_A12TS oc8051_decoder1_u336 ( .A(oc8051_decoder1_n98), .Y(
        oc8051_decoder1_n353) );
  INV_X0P5B_A12TS oc8051_decoder1_u335 ( .A(oc8051_decoder1_n25), .Y(
        oc8051_decoder1_n44) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u334 ( .A0(oc8051_decoder1_n9), .A1(
        oc8051_decoder1_n54), .A2(oc8051_decoder1_n409), .B0(
        oc8051_decoder1_n353), .B1(oc8051_decoder1_n44), .Y(
        oc8051_decoder1_n404) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u333 ( .A0(oc8051_decoder1_n386), .A1(
        oc8051_decoder1_n36), .B0(oc8051_decoder1_n387), .C0(
        oc8051_decoder1_n404), .Y(oc8051_decoder1_n385) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u332 ( .A(oc8051_decoder1_n277), .B(
        oc8051_decoder1_n385), .Y(istb) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u331 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n18) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u330 ( .A0(oc8051_decoder1_n82), .A1(
        oc8051_decoder1_n21), .B0(oc8051_decoder1_n18), .Y(
        oc8051_decoder1_n251) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u329 ( .A(oc8051_decoder1_n251), .B(
        oc8051_decoder1_n161), .S0(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n380) );
  INV_X0P5B_A12TS oc8051_decoder1_u328 ( .A(oc8051_decoder1_n105), .Y(
        oc8051_decoder1_n47) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u327 ( .A(oc8051_decoder1_n185), .B(
        oc8051_decoder1_n47), .Y(oc8051_decoder1_n138) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u326 ( .A0(oc8051_decoder1_n138), .A1(
        oc8051_decoder1_n178), .B0(oc8051_decoder1_n40), .Y(
        oc8051_decoder1_n381) );
  INV_X0P5B_A12TS oc8051_decoder1_u325 ( .A(oc8051_decoder1_n193), .Y(
        oc8051_decoder1_n8) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u324 ( .A(oc8051_decoder1_n165), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n136) );
  INV_X0P5B_A12TS oc8051_decoder1_u323 ( .A(oc8051_decoder1_n136), .Y(
        oc8051_decoder1_n154) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u322 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n375), .B0(op1_cur[1]), .Y(oc8051_decoder1_n384) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u321 ( .A0(oc8051_decoder1_n8), .A1(
        oc8051_decoder1_n186), .B0(oc8051_decoder1_n154), .B1(
        oc8051_decoder1_n14), .C0(oc8051_decoder1_n384), .Y(
        oc8051_decoder1_n382) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u320 ( .A(oc8051_decoder1_n54), .B(
        op1_cur[1]), .Y(oc8051_decoder1_n245) );
  INV_X0P5B_A12TS oc8051_decoder1_u319 ( .A(oc8051_decoder1_n245), .Y(
        oc8051_decoder1_n142) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u318 ( .A(oc8051_decoder1_n9), .B(
        op1_cur[2]), .C(oc8051_decoder1_n142), .Y(oc8051_decoder1_n383) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u317 ( .A0(oc8051_decoder1_n380), .A1(
        oc8051_decoder1_n67), .A2(oc8051_decoder1_n381), .B0(
        oc8051_decoder1_n382), .B1(oc8051_decoder1_n383), .Y(
        oc8051_decoder1_n377) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u316 ( .A(oc8051_decoder1_n125), .B(
        oc8051_decoder1_n33), .Y(oc8051_decoder1_n144) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u315 ( .A(oc8051_decoder1_n139), .B(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n49) );
  INV_X0P5B_A12TS oc8051_decoder1_u314 ( .A(oc8051_decoder1_n49), .Y(
        oc8051_decoder1_n176) );
  INV_X0P5B_A12TS oc8051_decoder1_u313 ( .A(oc8051_decoder1_n144), .Y(
        oc8051_decoder1_n126) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u312 ( .A(oc8051_decoder1_n126), .B(
        oc8051_decoder1_n9), .Y(oc8051_decoder1_n166) );
  INV_X0P5B_A12TS oc8051_decoder1_u311 ( .A(oc8051_decoder1_n166), .Y(
        oc8051_decoder1_n330) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u310 ( .A(oc8051_decoder1_n176), .B(
        oc8051_decoder1_n330), .Y(oc8051_decoder1_n182) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u309 ( .A(oc8051_decoder1_n330), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n119) );
  OA22_X0P5M_A12TS oc8051_decoder1_u308 ( .A0(oc8051_decoder1_n251), .A1(
        oc8051_decoder1_n119), .B0(oc8051_decoder1_n379), .B1(
        oc8051_decoder1_n125), .Y(oc8051_decoder1_n378) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u307 ( .A0(oc8051_decoder1_n377), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n182), .C0(
        oc8051_decoder1_n378), .Y(oc8051_decoder1_n388) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u306 ( .A(oc8051_decoder1_n90), .B(
        op1_cur[1]), .Y(oc8051_decoder1_n355) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u305 ( .A(oc8051_decoder1_n244), .B(
        oc8051_decoder1_n281), .Y(oc8051_decoder1_n150) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u304 ( .A(oc8051_decoder1_n21), .B(
        oc8051_decoder1_n53), .Y(oc8051_decoder1_n217) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u303 ( .A(oc8051_decoder1_n257), .B(
        oc8051_decoder1_n136), .Y(oc8051_decoder1_n376) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u302 ( .A(oc8051_decoder1_n109), .B(
        oc8051_decoder1_n376), .S0(oc8051_decoder1_n21), .Y(
        oc8051_decoder1_n374) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u301 ( .A(oc8051_decoder1_n375), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n326) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u300 ( .A(oc8051_decoder1_n90), .B(
        oc8051_decoder1_n40), .Y(oc8051_decoder1_n157) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u299 ( .A(oc8051_decoder1_n326), .B(
        oc8051_decoder1_n157), .Y(oc8051_decoder1_n20) );
  AOI2XB1_X0P5M_A12TS oc8051_decoder1_u298 ( .A1N(oc8051_decoder1_n217), .A0(
        oc8051_decoder1_n374), .B0(oc8051_decoder1_n20), .Y(
        oc8051_decoder1_n351) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u297 ( .A0(oc8051_decoder1_n155), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n71), .B1(
        oc8051_decoder1_n48), .Y(oc8051_decoder1_n367) );
  INV_X0P5B_A12TS oc8051_decoder1_u296 ( .A(oc8051_decoder1_n367), .Y(
        oc8051_decoder1_n201) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u295 ( .A(oc8051_decoder1_n67), .B(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n37) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u294 ( .A0(oc8051_decoder1_n201), .A1(
        oc8051_decoder1_n131), .B0(oc8051_decoder1_n37), .C0(
        oc8051_decoder1_n373), .Y(oc8051_decoder1_n369) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u293 ( .A(oc8051_decoder1_n40), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n370) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u292 ( .A0(oc8051_decoder1_n185), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n14), .B1(op1_cur[0]), .Y(
        oc8051_decoder1_n371) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u291 ( .A(oc8051_decoder1_n59), .B(
        oc8051_decoder1_n165), .S0(oc8051_decoder1_n137), .Y(
        oc8051_decoder1_n372) );
  INV_X0P5B_A12TS oc8051_decoder1_u290 ( .A(oc8051_decoder1_n157), .Y(
        oc8051_decoder1_n6) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u289 ( .A(oc8051_decoder1_n6), .B(
        op1_cur[1]), .Y(oc8051_decoder1_n350) );
  INV_X0P5B_A12TS oc8051_decoder1_u288 ( .A(oc8051_decoder1_n350), .Y(
        oc8051_decoder1_n146) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u287 ( .A0(oc8051_decoder1_n369), .A1(
        oc8051_decoder1_n370), .A2(oc8051_decoder1_n371), .B0(
        oc8051_decoder1_n372), .B1(oc8051_decoder1_n146), .Y(
        oc8051_decoder1_n368) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u286 ( .A0(oc8051_decoder1_n355), .A1(
        oc8051_decoder1_n150), .B0(oc8051_decoder1_n351), .C0(
        oc8051_decoder1_n368), .Y(oc8051_decoder1_n366) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u285 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n366), .B0(oc8051_decoder1_n330), .B1(
        oc8051_decoder1_n367), .Y(oc8051_decoder1_n365) );
  AO1B2_X0P5M_A12TS oc8051_decoder1_u284 ( .B0(psw_set[0]), .B1(wait_data), 
        .A0N(oc8051_decoder1_n365), .Y(oc8051_decoder1_n389) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u283 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n82), .Y(oc8051_decoder1_n356) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u282 ( .A(oc8051_decoder1_n281), .B(
        oc8051_decoder1_n47), .Y(oc8051_decoder1_n292) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u281 ( .A(oc8051_decoder1_n292), .B(
        oc8051_decoder1_n166), .Y(oc8051_decoder1_n128) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u280 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n40), .A2(oc8051_decoder1_n330), .B0(
        oc8051_decoder1_n128), .Y(oc8051_decoder1_n357) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u279 ( .A(oc8051_decoder1_n281), .B(
        oc8051_decoder1_n42), .Y(oc8051_decoder1_n202) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u278 ( .A(oc8051_decoder1_n217), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n13) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u277 ( .A0(oc8051_decoder1_n155), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n202), .C0(
        oc8051_decoder1_n13), .Y(oc8051_decoder1_n362) );
  INV_X0P5B_A12TS oc8051_decoder1_u276 ( .A(oc8051_decoder1_n356), .Y(
        oc8051_decoder1_n70) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u275 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n40), .B0(oc8051_decoder1_n176), .C0(op1_cur[1]), .Y(
        oc8051_decoder1_n364) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u274 ( .A0(oc8051_decoder1_n25), .A1(
        oc8051_decoder1_n292), .B0(oc8051_decoder1_n326), .B1(
        oc8051_decoder1_n48), .C0(oc8051_decoder1_n364), .Y(
        oc8051_decoder1_n363) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u273 ( .A0(oc8051_decoder1_n178), .A1(
        oc8051_decoder1_n362), .B0(oc8051_decoder1_n70), .B1(
        oc8051_decoder1_n185), .C0(oc8051_decoder1_n363), .Y(
        oc8051_decoder1_n360) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u272 ( .A(oc8051_decoder1_n50), .B(
        oc8051_decoder1_n157), .C(oc8051_decoder1_n265), .Y(
        oc8051_decoder1_n279) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u271 ( .A0(oc8051_decoder1_n47), .A1(
        op1_cur[0]), .A2(oc8051_decoder1_n146), .B0(oc8051_decoder1_n279), .Y(
        oc8051_decoder1_n361) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u270 ( .A0(oc8051_decoder1_n360), .A1(
        oc8051_decoder1_n26), .B0(oc8051_decoder1_n270), .B1(
        oc8051_decoder1_n356), .C0(oc8051_decoder1_n361), .Y(
        oc8051_decoder1_n359) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u269 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n359), .B0(src_sel2[0]), .B1(wait_data), .Y(
        oc8051_decoder1_n358) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u268 ( .A0(oc8051_decoder1_n119), .A1(
        oc8051_decoder1_n356), .B0(oc8051_decoder1_n357), .C0(
        oc8051_decoder1_n358), .Y(oc8051_decoder1_n390) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u267 ( .A(op1_cur[2]), .B(
        oc8051_decoder1_n69), .C(oc8051_decoder1_n54), .Y(oc8051_decoder1_n116) );
  INV_X0P5B_A12TS oc8051_decoder1_u266 ( .A(oc8051_decoder1_n116), .Y(
        oc8051_decoder1_n293) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u265 ( .A(oc8051_decoder1_n126), .B(
        oc8051_decoder1_n293), .Y(oc8051_decoder1_n212) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u264 ( .A0(oc8051_decoder1_n155), .A1(
        oc8051_decoder1_n166), .B0(oc8051_decoder1_n50), .B1(
        oc8051_decoder1_n212), .Y(oc8051_decoder1_n347) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u263 ( .A0(oc8051_decoder1_n137), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n55), .Y(
        oc8051_decoder1_n262) );
  INV_X0P5B_A12TS oc8051_decoder1_u262 ( .A(oc8051_decoder1_n262), .Y(
        oc8051_decoder1_n349) );
  INV_X0P5B_A12TS oc8051_decoder1_u261 ( .A(oc8051_decoder1_n355), .Y(
        oc8051_decoder1_n16) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u260 ( .A(oc8051_decoder1_n265), .B(
        oc8051_decoder1_n155), .C(oc8051_decoder1_n26), .Y(
        oc8051_decoder1_n287) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u259 ( .A(oc8051_decoder1_n67), .B(
        oc8051_decoder1_n185), .Y(oc8051_decoder1_n27) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u258 ( .A(oc8051_decoder1_n27), .B(
        oc8051_decoder1_n14), .C(oc8051_decoder1_n82), .Y(oc8051_decoder1_n354) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u257 ( .A0(oc8051_decoder1_n353), .A1(
        oc8051_decoder1_n16), .B0(oc8051_decoder1_n287), .C0(
        oc8051_decoder1_n354), .Y(oc8051_decoder1_n352) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u256 ( .A0(oc8051_decoder1_n349), .A1(
        oc8051_decoder1_n350), .B0(oc8051_decoder1_n351), .C0(
        oc8051_decoder1_n352), .Y(oc8051_decoder1_n348) );
  AOI222_X0P5M_A12TS oc8051_decoder1_u255 ( .A0(cy_sel[0]), .A1(wait_data), 
        .B0(oc8051_decoder1_n156), .B1(oc8051_decoder1_n347), .C0(
        oc8051_decoder1_n126), .C1(oc8051_decoder1_n348), .Y(
        oc8051_decoder1_n342) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u254 ( .A(oc8051_decoder1_n47), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n211) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u253 ( .A0(op1_cur[1]), .A1(
        oc8051_decoder1_n225), .B0(oc8051_decoder1_n211), .C0(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n344) );
  INV_X0P5B_A12TS oc8051_decoder1_u252 ( .A(oc8051_decoder1_n212), .Y(
        oc8051_decoder1_n273) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u251 ( .A(oc8051_decoder1_n166), .B(
        oc8051_decoder1_n82), .C(oc8051_decoder1_n48), .Y(oc8051_decoder1_n345) );
  INV_X0P5B_A12TS oc8051_decoder1_u250 ( .A(oc8051_decoder1_n182), .Y(
        oc8051_decoder1_n346) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u249 ( .A0(oc8051_decoder1_n344), .A1(
        oc8051_decoder1_n273), .B0(oc8051_decoder1_n345), .C0(
        oc8051_decoder1_n346), .Y(oc8051_decoder1_n343) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u248 ( .A(oc8051_decoder1_n342), .B(
        oc8051_decoder1_n343), .Y(oc8051_decoder1_n391) );
  INV_X0P5B_A12TS oc8051_decoder1_u247 ( .A(oc8051_decoder1_n27), .Y(
        oc8051_decoder1_n189) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u246 ( .A(oc8051_decoder1_n44), .B(
        oc8051_decoder1_n61), .C(oc8051_decoder1_n293), .Y(
        oc8051_decoder1_n114) );
  INV_X0P5B_A12TS oc8051_decoder1_u245 ( .A(oc8051_decoder1_n115), .Y(
        oc8051_decoder1_n341) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u244 ( .A(oc8051_decoder1_n9), .B(
        oc8051_decoder1_n54), .C(oc8051_decoder1_n341), .Y(
        oc8051_decoder1_n113) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u243 ( .A(oc8051_decoder1_n341), .B(
        oc8051_decoder1_n54), .C(oc8051_decoder1_n25), .D(op1_cur[2]), .Y(
        oc8051_decoder1_n340) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u242 ( .A(oc8051_decoder1_n114), .B(
        oc8051_decoder1_n113), .C(oc8051_decoder1_n340), .Y(
        oc8051_decoder1_n339) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u241 ( .A(oc8051_decoder1_n224), .B(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n325) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u240 ( .A(op1_cur[0]), .B(op1_cur[1]), .C(
        oc8051_decoder1_n224), .Y(oc8051_decoder1_n102) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u239 ( .A0(oc8051_decoder1_n325), .A1(
        oc8051_decoder1_n226), .B0(oc8051_decoder1_n102), .B1(
        oc8051_decoder1_n236), .Y(oc8051_decoder1_n291) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u238 ( .A0(oc8051_decoder1_n275), .A1(
        oc8051_decoder1_n189), .B0(oc8051_decoder1_n339), .C0(
        oc8051_decoder1_n291), .Y(oc8051_decoder1_n335) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u237 ( .A(src_sel2[1]), .B(wait_data), .Y(
        oc8051_decoder1_n336) );
  INV_X0P5B_A12TS oc8051_decoder1_u236 ( .A(oc8051_decoder1_n226), .Y(
        oc8051_decoder1_n207) );
  INV_X0P5B_A12TS oc8051_decoder1_u235 ( .A(oc8051_decoder1_n48), .Y(
        oc8051_decoder1_n135) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u234 ( .A(oc8051_decoder1_n135), .B(
        oc8051_decoder1_n71), .Y(oc8051_decoder1_n12) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u233 ( .A0(oc8051_decoder1_n98), .A1(
        oc8051_decoder1_n12), .B0(oc8051_decoder1_n166), .Y(
        oc8051_decoder1_n338) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u232 ( .A0(oc8051_decoder1_n207), .A1(
        oc8051_decoder1_n178), .A2(oc8051_decoder1_n273), .B0(
        oc8051_decoder1_n338), .Y(oc8051_decoder1_n337) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u231 ( .A0(oc8051_decoder1_n335), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n336), .C0(
        oc8051_decoder1_n337), .Y(oc8051_decoder1_n392) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u230 ( .A0(oc8051_decoder1_n115), .A1(
        oc8051_decoder1_n193), .A2(oc8051_decoder1_n334), .B0(
        oc8051_decoder1_n114), .Y(oc8051_decoder1_n332) );
  INV_X0P5B_A12TS oc8051_decoder1_u229 ( .A(oc8051_decoder1_n102), .Y(
        oc8051_decoder1_n269) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u228 ( .A0(oc8051_decoder1_n8), .A1(
        oc8051_decoder1_n224), .B0(oc8051_decoder1_n269), .Y(
        oc8051_decoder1_n324) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u227 ( .A0(oc8051_decoder1_n82), .A1(
        oc8051_decoder1_n225), .B0(oc8051_decoder1_n236), .C0(
        oc8051_decoder1_n324), .Y(oc8051_decoder1_n333) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u226 ( .A0(oc8051_decoder1_n189), .A1(
        oc8051_decoder1_n207), .B0(oc8051_decoder1_n332), .C0(
        oc8051_decoder1_n333), .Y(oc8051_decoder1_n327) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u225 ( .A(oc8051_decoder1_n225), .B(
        oc8051_decoder1_n212), .Y(oc8051_decoder1_n331) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u224 ( .A0(op1_cur[1]), .A1(
        oc8051_decoder1_n44), .B0(oc8051_decoder1_n82), .C0(
        oc8051_decoder1_n331), .Y(oc8051_decoder1_n328) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u223 ( .A0(oc8051_decoder1_n54), .A1(
        oc8051_decoder1_n226), .B0(oc8051_decoder1_n49), .Y(
        oc8051_decoder1_n197) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u222 ( .A0(oc8051_decoder1_n330), .A1(
        oc8051_decoder1_n197), .B0(cy_sel[1]), .B1(wait_data), .Y(
        oc8051_decoder1_n329) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u221 ( .A0(oc8051_decoder1_n327), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n328), .C0(
        oc8051_decoder1_n329), .Y(oc8051_decoder1_n393) );
  INV_X0P5B_A12TS oc8051_decoder1_u220 ( .A(oc8051_decoder1_n326), .Y(
        oc8051_decoder1_n320) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u219 ( .A(oc8051_decoder1_n47), .B(
        oc8051_decoder1_n21), .Y(oc8051_decoder1_n181) );
  INV_X0P5B_A12TS oc8051_decoder1_u218 ( .A(oc8051_decoder1_n181), .Y(
        oc8051_decoder1_n219) );
  INV_X0P5B_A12TS oc8051_decoder1_u217 ( .A(oc8051_decoder1_n325), .Y(
        oc8051_decoder1_n60) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u216 ( .A(oc8051_decoder1_n219), .B(
        oc8051_decoder1_n60), .Y(oc8051_decoder1_n78) );
  OA22_X0P5M_A12TS oc8051_decoder1_u215 ( .A0(oc8051_decoder1_n225), .A1(
        oc8051_decoder1_n324), .B0(oc8051_decoder1_n105), .B1(
        oc8051_decoder1_n102), .Y(oc8051_decoder1_n323) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u214 ( .A0(oc8051_decoder1_n219), .A1(
        oc8051_decoder1_n322), .B0(oc8051_decoder1_n78), .C0(
        oc8051_decoder1_n323), .Y(oc8051_decoder1_n321) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u213 ( .A0(oc8051_decoder1_n273), .A1(
        oc8051_decoder1_n320), .A2(oc8051_decoder1_n70), .B0(
        oc8051_decoder1_n126), .B1(oc8051_decoder1_n321), .Y(
        oc8051_decoder1_n319) );
  AO1B2_X0P5M_A12TS oc8051_decoder1_u212 ( .B0(src_sel3), .B1(wait_data), 
        .A0N(oc8051_decoder1_n319), .Y(oc8051_decoder1_n394) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u211 ( .A(wait_data), .B(mem_wait), .Y(
        oc8051_decoder1_n296) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u210 ( .A0(oc8051_decoder1_n296), .A1(
        oc8051_decoder1_n316), .B0(oc8051_decoder1_n317), .C0(
        oc8051_decoder1_n318), .Y(oc8051_decoder1_n395) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u209 ( .A(oc8051_decoder1_n314), .B(
        oc8051_decoder1_n315), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n396) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u208 ( .A(oc8051_decoder1_n299), .B(
        oc8051_decoder1_n313), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n397) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u207 ( .A(oc8051_decoder1_n311), .B(
        oc8051_decoder1_n312), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n398) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u206 ( .A(oc8051_decoder1_n300), .B(
        oc8051_decoder1_n310), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n399) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u205 ( .A(oc8051_decoder1_n308), .B(
        oc8051_decoder1_n309), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n400) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u204 ( .A(oc8051_decoder1_n306), .B(
        oc8051_decoder1_n307), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n401) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u203 ( .A(oc8051_decoder1_n304), .B(
        oc8051_decoder1_n305), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n402) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u202 ( .A(oc8051_decoder1_n301), .B(
        oc8051_decoder1_n302), .S0(oc8051_decoder1_n303), .Y(
        oc8051_decoder1_n403) );
  XOR2_X0P5M_A12TS oc8051_decoder1_u201 ( .A(op1_n[7]), .B(op1_n[5]), .Y(
        oc8051_decoder1_n298) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u200 ( .A0(oc8051_decoder1_n298), .A1(
        oc8051_decoder1_n299), .A2(op1_n[1]), .B0(op1_n[2]), .B1(
        oc8051_decoder1_n300), .Y(oc8051_decoder1_n297) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u199 ( .A(oc8051_decoder1_state_0_), .B(
        oc8051_decoder1_n297), .Y(oc8051_decoder1_n295) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u198 ( .A(oc8051_decoder1_state_0_), .B(
        oc8051_decoder1_n295), .S0(oc8051_decoder1_n296), .Y(
        oc8051_decoder1_n294) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u197 ( .A0(mem_wait), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n294), .Y(
        oc8051_decoder1_n405) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u196 ( .A(oc8051_decoder1_n293), .B(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n180) );
  INV_X0P5B_A12TS oc8051_decoder1_u195 ( .A(oc8051_decoder1_n52), .Y(
        oc8051_decoder1_n68) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u194 ( .A(oc8051_decoder1_n68), .B(
        oc8051_decoder1_n293), .C(oc8051_decoder1_n82), .D(oc8051_decoder1_n22), .Y(oc8051_decoder1_n122) );
  OA21_X0P5M_A12TS oc8051_decoder1_u193 ( .A0(oc8051_decoder1_n180), .A1(
        oc8051_decoder1_n181), .B0(oc8051_decoder1_n122), .Y(
        oc8051_decoder1_n255) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u192 ( .A(oc8051_decoder1_n277), .B(
        oc8051_decoder1_n255), .Y(oc8051_decoder1_n228) );
  INV_X0P5B_A12TS oc8051_decoder1_u191 ( .A(oc8051_decoder1_n228), .Y(
        oc8051_decoder1_n229) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u190 ( .A(oc8051_decoder1_n219), .B(
        oc8051_decoder1_n44), .C(oc8051_decoder1_n273), .Y(
        oc8051_decoder1_n213) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u189 ( .A0(oc8051_decoder1_n408), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n229), .C0(
        oc8051_decoder1_n213), .Y(oc8051_decoder1_n412) );
  INV_X0P5B_A12TS oc8051_decoder1_u188 ( .A(oc8051_decoder1_n292), .Y(
        oc8051_decoder1_n290) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u187 ( .A0(oc8051_decoder1_n290), .A1(
        oc8051_decoder1_n36), .B0(oc8051_decoder1_n291), .C0(
        oc8051_decoder1_n126), .Y(oc8051_decoder1_n288) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u186 ( .A0(oc8051_decoder1_n61), .A1(
        op1_cur[1]), .A2(oc8051_decoder1_n273), .B0(oc8051_decoder1_n228), .Y(
        oc8051_decoder1_n289) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u185 ( .A0(oc8051_decoder1_n406), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n288), .C0(
        oc8051_decoder1_n289), .Y(oc8051_decoder1_n413) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u184 ( .A0(oc8051_decoder1_n42), .A1(
        oc8051_decoder1_n16), .B0(oc8051_decoder1_n75), .Y(
        oc8051_decoder1_n284) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u183 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n23), .B0(oc8051_decoder1_n104), .Y(
        oc8051_decoder1_n190) );
  INV_X0P5B_A12TS oc8051_decoder1_u182 ( .A(oc8051_decoder1_n190), .Y(
        oc8051_decoder1_n286) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u181 ( .A0(oc8051_decoder1_n286), .A1(
        oc8051_decoder1_n189), .B0(oc8051_decoder1_n287), .C0(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n285) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u180 ( .A0(oc8051_decoder1_n284), .A1(
        oc8051_decoder1_n14), .A2(oc8051_decoder1_n137), .B0(
        oc8051_decoder1_n285), .Y(oc8051_decoder1_n278) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u179 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n131), .B0(oc8051_decoder1_n69), .Y(
        oc8051_decoder1_n41) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u178 ( .A(oc8051_decoder1_n283), .B(
        oc8051_decoder1_n12), .C(oc8051_decoder1_n41), .Y(oc8051_decoder1_n282) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u177 ( .A0(oc8051_decoder1_n281), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n40), .B1(
        oc8051_decoder1_n265), .C0(oc8051_decoder1_n282), .Y(
        oc8051_decoder1_n280) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u176 ( .A0(oc8051_decoder1_n278), .A1(
        oc8051_decoder1_n279), .A2(oc8051_decoder1_n280), .B0(
        oc8051_decoder1_n126), .Y(oc8051_decoder1_n271) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u175 ( .A0(oc8051_decoder1_n50), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n47), .Y(
        oc8051_decoder1_n274) );
  AND4_X0P5M_A12TS oc8051_decoder1_u174 ( .A(oc8051_decoder1_n42), .B(
        oc8051_decoder1_n224), .C(oc8051_decoder1_n14), .D(oc8051_decoder1_n25), .Y(oc8051_decoder1_n276) );
  INV_X0P5B_A12TS oc8051_decoder1_u173 ( .A(oc8051_decoder1_n277), .Y(
        oc8051_decoder1_n183) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u172 ( .A0(oc8051_decoder1_n275), .A1(
        oc8051_decoder1_n269), .B0(oc8051_decoder1_n276), .C0(
        oc8051_decoder1_n183), .Y(oc8051_decoder1_n267) );
  INV_X0P5B_A12TS oc8051_decoder1_u171 ( .A(oc8051_decoder1_n267), .Y(
        oc8051_decoder1_n241) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u170 ( .A0(oc8051_decoder1_n273), .A1(
        oc8051_decoder1_n14), .A2(oc8051_decoder1_n274), .B0(
        oc8051_decoder1_n241), .Y(oc8051_decoder1_n272) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u169 ( .A0(oc8051_decoder1_n407), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n271), .C0(
        oc8051_decoder1_n272), .Y(oc8051_decoder1_n414) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u168 ( .A(oc8051_decoder1_n165), .B(
        oc8051_decoder1_n90), .C(oc8051_decoder1_n44), .Y(oc8051_decoder1_n200) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u167 ( .A0(oc8051_decoder1_n270), .A1(
        oc8051_decoder1_n226), .B0(oc8051_decoder1_n200), .Y(
        oc8051_decoder1_n218) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u166 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n111), .B0(oc8051_decoder1_n218), .Y(
        oc8051_decoder1_n230) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u165 ( .A0(oc8051_decoder1_n219), .A1(
        oc8051_decoder1_n269), .A2(oc8051_decoder1_n126), .B0(src_sel1[2]), 
        .B1(wait_data), .Y(oc8051_decoder1_n268) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u164 ( .A(oc8051_decoder1_n267), .B(
        oc8051_decoder1_n230), .C(oc8051_decoder1_n268), .Y(
        oc8051_decoder1_n415) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u163 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n185), .B0(oc8051_decoder1_n161), .Y(
        oc8051_decoder1_n266) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u162 ( .A(oc8051_decoder1_n265), .B(
        oc8051_decoder1_n266), .S0(oc8051_decoder1_n164), .Y(
        oc8051_decoder1_n252) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u161 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n185), .B1(
        oc8051_decoder1_n50), .Y(oc8051_decoder1_n259) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u160 ( .A(oc8051_decoder1_n154), .B(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n264) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u159 ( .A(oc8051_decoder1_n217), .B(
        op1_cur[0]), .Y(oc8051_decoder1_n38) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u158 ( .A0(oc8051_decoder1_n137), .A1(
        oc8051_decoder1_n165), .B0(oc8051_decoder1_n38), .Y(
        oc8051_decoder1_n250) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u157 ( .A(oc8051_decoder1_n264), .B(
        oc8051_decoder1_n250), .S0(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n263) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u156 ( .A0(oc8051_decoder1_n135), .A1(
        oc8051_decoder1_n262), .B0(oc8051_decoder1_n263), .Y(
        oc8051_decoder1_n261) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u155 ( .A(oc8051_decoder1_n252), .B(
        oc8051_decoder1_n261), .S0(oc8051_decoder1_n22), .Y(
        oc8051_decoder1_n260) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u154 ( .A0(oc8051_decoder1_n90), .A1(
        oc8051_decoder1_n259), .A2(oc8051_decoder1_n207), .B0(
        oc8051_decoder1_n260), .B1(oc8051_decoder1_n67), .Y(
        oc8051_decoder1_n258) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u153 ( .A0(oc8051_decoder1_n11), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n257), .C0(
        oc8051_decoder1_n258), .Y(oc8051_decoder1_n256) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u152 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n256), .B0(oc8051_decoder1_n241), .Y(
        oc8051_decoder1_n253) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u151 ( .A(oc8051_decoder1_state_1_), .B(
        oc8051_decoder1_n125), .C(oc8051_decoder1_state_0_), .Y(
        oc8051_decoder1_n184) );
  NAND3B_X0P5M_A12TS oc8051_decoder1_u150 ( .AN(oc8051_decoder1_n180), .B(
        oc8051_decoder1_n82), .C(oc8051_decoder1_n21), .Y(oc8051_decoder1_n101) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u149 ( .A0(oc8051_decoder1_n184), .A1(
        oc8051_decoder1_n101), .B0(oc8051_decoder1_n255), .B1(
        oc8051_decoder1_n30), .C0(oc8051_decoder1_n229), .Y(
        oc8051_decoder1_n203) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u148 ( .A0(src_sel1[1]), .A1(wait_data), 
        .B0(oc8051_decoder1_n203), .Y(oc8051_decoder1_n254) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u147 ( .A0(oc8051_decoder1_n166), .A1(
        oc8051_decoder1_n252), .B0(oc8051_decoder1_n253), .C0(
        oc8051_decoder1_n254), .Y(oc8051_decoder1_n416) );
  OAI222_X0P5M_A12TS oc8051_decoder1_u146 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n132), .B0(oc8051_decoder1_n54), .B1(
        oc8051_decoder1_n251), .C0(oc8051_decoder1_n156), .C1(
        oc8051_decoder1_n155), .Y(oc8051_decoder1_n237) );
  INV_X0P5B_A12TS oc8051_decoder1_u145 ( .A(oc8051_decoder1_n237), .Y(
        oc8051_decoder1_n247) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u144 ( .A(oc8051_decoder1_n25), .B(
        oc8051_decoder1_n186), .Y(oc8051_decoder1_n249) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u143 ( .A(oc8051_decoder1_n249), .B(
        oc8051_decoder1_n250), .S0(oc8051_decoder1_n54), .Y(
        oc8051_decoder1_n248) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u142 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n247), .B0(oc8051_decoder1_n48), .B1(
        oc8051_decoder1_n23), .C0(oc8051_decoder1_n248), .Y(
        oc8051_decoder1_n242) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u141 ( .A(oc8051_decoder1_n154), .B(
        oc8051_decoder1_n38), .S0(op1_cur[1]), .Y(oc8051_decoder1_n246) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u140 ( .A0(op1_cur[0]), .A1(
        oc8051_decoder1_n156), .B0(oc8051_decoder1_n244), .B1(
        oc8051_decoder1_n245), .C0(oc8051_decoder1_n246), .Y(
        oc8051_decoder1_n243) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u139 ( .A(oc8051_decoder1_n242), .B(
        oc8051_decoder1_n243), .S0(oc8051_decoder1_n131), .Y(
        oc8051_decoder1_n240) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u138 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n69), .A2(oc8051_decoder1_n240), .B0(
        oc8051_decoder1_n241), .Y(oc8051_decoder1_n238) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u137 ( .A0(src_sel1[0]), .A1(wait_data), 
        .B0(oc8051_decoder1_n203), .Y(oc8051_decoder1_n239) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u136 ( .A0(oc8051_decoder1_n166), .A1(
        oc8051_decoder1_n237), .B0(oc8051_decoder1_n238), .C0(
        oc8051_decoder1_n239), .Y(oc8051_decoder1_n417) );
  INV_X0P5B_A12TS oc8051_decoder1_u135 ( .A(oc8051_decoder1_n211), .Y(
        oc8051_decoder1_n222) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u134 ( .A(oc8051_decoder1_n126), .B(
        oc8051_decoder1_n60), .C(oc8051_decoder1_n222), .Y(
        oc8051_decoder1_n231) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u133 ( .A(oc8051_decoder1_n226), .B(
        oc8051_decoder1_n181), .Y(oc8051_decoder1_n108) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u132 ( .A0(oc8051_decoder1_n189), .A1(
        oc8051_decoder1_n108), .B0(oc8051_decoder1_n221), .B1(
        oc8051_decoder1_n67), .Y(oc8051_decoder1_n234) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u131 ( .A0(oc8051_decoder1_n11), .A1(
        oc8051_decoder1_n211), .A2(oc8051_decoder1_n236), .B0(
        oc8051_decoder1_n212), .Y(oc8051_decoder1_n235) );
  OAI21B_X0P5M_A12TS oc8051_decoder1_u130 ( .A0(oc8051_decoder1_n234), .A1(
        oc8051_decoder1_n144), .B0N(oc8051_decoder1_n235), .Y(
        oc8051_decoder1_n233) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u129 ( .A0(oc8051_decoder1_n233), .A1(
        op1_cur[1]), .B0(wait_data), .B1(oc8051_decoder1_ram_wr_sel_1_), .Y(
        oc8051_decoder1_n232) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u128 ( .A(oc8051_decoder1_n229), .B(
        oc8051_decoder1_n230), .C(oc8051_decoder1_n231), .D(
        oc8051_decoder1_n232), .Y(oc8051_decoder1_n418) );
  INV_X0P5B_A12TS oc8051_decoder1_u127 ( .A(oc8051_decoder1_ram_wr_sel_0_), 
        .Y(oc8051_decoder1_n28) );
  AND4_X0P5M_A12TS oc8051_decoder1_u126 ( .A(oc8051_decoder1_n207), .B(
        oc8051_decoder1_n90), .C(oc8051_decoder1_n185), .D(oc8051_decoder1_n22), .Y(oc8051_decoder1_n227) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u125 ( .A0(oc8051_decoder1_n218), .A1(
        oc8051_decoder1_n227), .B0(oc8051_decoder1_n111), .C0(
        oc8051_decoder1_n228), .Y(oc8051_decoder1_n188) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u124 ( .A0(oc8051_decoder1_n115), .A1(
        oc8051_decoder1_n225), .A2(oc8051_decoder1_n226), .B0(
        oc8051_decoder1_n22), .Y(oc8051_decoder1_n223) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u123 ( .A0(oc8051_decoder1_n222), .A1(
        oc8051_decoder1_n223), .B0(oc8051_decoder1_n137), .C0(
        oc8051_decoder1_n224), .Y(oc8051_decoder1_n214) );
  AO22_X0P5M_A12TS oc8051_decoder1_u122 ( .A0(oc8051_decoder1_n69), .A1(
        oc8051_decoder1_n221), .B0(oc8051_decoder1_n108), .B1(
        oc8051_decoder1_n189), .Y(oc8051_decoder1_n220) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u121 ( .A0(oc8051_decoder1_n54), .A1(
        oc8051_decoder1_n41), .A2(oc8051_decoder1_n219), .B0(
        oc8051_decoder1_n44), .B1(oc8051_decoder1_n220), .Y(
        oc8051_decoder1_n215) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u120 ( .A0(oc8051_decoder1_n60), .A1(
        oc8051_decoder1_n61), .B0(oc8051_decoder1_n75), .B1(
        oc8051_decoder1_n217), .C0(oc8051_decoder1_n218), .Y(
        oc8051_decoder1_n216) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u119 ( .A(oc8051_decoder1_n214), .B(
        oc8051_decoder1_n114), .C(oc8051_decoder1_n215), .D(
        oc8051_decoder1_n216), .Y(oc8051_decoder1_n209) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u118 ( .A0(oc8051_decoder1_n211), .A1(
        oc8051_decoder1_n25), .A2(oc8051_decoder1_n212), .B0(
        oc8051_decoder1_n213), .Y(oc8051_decoder1_n210) );
  AOI21_X0P5M_A12TS oc8051_decoder1_u117 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n209), .B0(oc8051_decoder1_n210), .Y(
        oc8051_decoder1_n208) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u116 ( .A0(oc8051_decoder1_n28), .A1(
        oc8051_decoder1_n125), .B0(oc8051_decoder1_n188), .C0(
        oc8051_decoder1_n208), .Y(oc8051_decoder1_n419) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u115 ( .A0(oc8051_decoder1_n135), .A1(
        oc8051_decoder1_n161), .B0(oc8051_decoder1_n207), .B1(
        oc8051_decoder1_n54), .Y(oc8051_decoder1_n206) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u114 ( .A0(oc8051_decoder1_n90), .A1(
        oc8051_decoder1_n206), .B0(oc8051_decoder1_n101), .Y(
        oc8051_decoder1_n205) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u113 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n205), .B0(psw_set[1]), .B1(wait_data), .Y(
        oc8051_decoder1_n204) );
  NAND2B_X0P5M_A12TS oc8051_decoder1_u112 ( .AN(oc8051_decoder1_n203), .B(
        oc8051_decoder1_n204), .Y(oc8051_decoder1_n420) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u111 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n47), .C0(
        oc8051_decoder1_n44), .Y(oc8051_decoder1_n198) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u110 ( .A(oc8051_decoder1_n201), .B(
        oc8051_decoder1_n202), .C(oc8051_decoder1_n41), .D(oc8051_decoder1_n13), .Y(oc8051_decoder1_n199) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u109 ( .A0(oc8051_decoder1_n116), .A1(
        oc8051_decoder1_n198), .B0(oc8051_decoder1_n199), .C0(
        oc8051_decoder1_n200), .Y(oc8051_decoder1_n191) );
  INV_X0P5B_A12TS oc8051_decoder1_u108 ( .A(oc8051_decoder1_n197), .Y(
        oc8051_decoder1_n196) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u107 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n13), .B0(oc8051_decoder1_n196), .B1(
        oc8051_decoder1_n193), .Y(oc8051_decoder1_n195) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u106 ( .A0(oc8051_decoder1_n176), .A1(
        oc8051_decoder1_n178), .B0(oc8051_decoder1_n195), .C0(
        oc8051_decoder1_n90), .Y(oc8051_decoder1_n194) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u105 ( .A0(oc8051_decoder1_n193), .A1(
        oc8051_decoder1_n157), .A2(oc8051_decoder1_n82), .B0(
        oc8051_decoder1_n194), .Y(oc8051_decoder1_n192) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u104 ( .A0(oc8051_decoder1_n189), .A1(
        oc8051_decoder1_n190), .B0(oc8051_decoder1_n191), .C0(
        oc8051_decoder1_n192), .Y(oc8051_decoder1_n187) );
  INV_X0P5B_A12TS oc8051_decoder1_u103 ( .A(oc8051_decoder1_wr), .Y(
        oc8051_decoder1_n1) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u102 ( .A0(oc8051_decoder1_n187), .A1(
        oc8051_decoder1_n144), .B0(oc8051_decoder1_n1), .B1(
        oc8051_decoder1_n125), .C0(oc8051_decoder1_n188), .Y(
        oc8051_decoder1_n421) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u101 ( .A(oc8051_decoder1_n185), .B(
        oc8051_decoder1_n18), .C(oc8051_decoder1_n186), .Y(
        oc8051_decoder1_n151) );
  INV_X0P5B_A12TS oc8051_decoder1_u100 ( .A(oc8051_decoder1_n184), .Y(
        oc8051_decoder1_n110) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u99 ( .A(oc8051_decoder1_n110), .B(
        oc8051_decoder1_n183), .C(oc8051_decoder1_n111), .Y(
        oc8051_decoder1_n123) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u98 ( .A0(oc8051_decoder1_n180), .A1(
        oc8051_decoder1_n123), .A2(oc8051_decoder1_n181), .B0(
        oc8051_decoder1_n182), .Y(oc8051_decoder1_n179) );
  INV_X0P5B_A12TS oc8051_decoder1_u97 ( .A(oc8051_decoder1_n179), .Y(
        oc8051_decoder1_n167) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u96 ( .A0(op1_cur[0]), .A1(
        oc8051_decoder1_n105), .B0(oc8051_decoder1_n59), .Y(
        oc8051_decoder1_n147) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u95 ( .A0(oc8051_decoder1_n132), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n105), .B1(
        oc8051_decoder1_n155), .Y(oc8051_decoder1_n177) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u94 ( .A0(op1_cur[1]), .A1(
        oc8051_decoder1_n176), .B0(oc8051_decoder1_n177), .B1(
        oc8051_decoder1_n178), .Y(oc8051_decoder1_n175) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u93 ( .A0(oc8051_decoder1_n175), .A1(
        oc8051_decoder1_n151), .A2(oc8051_decoder1_n150), .B0(
        oc8051_decoder1_n26), .Y(oc8051_decoder1_n171) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u92 ( .A0(oc8051_decoder1_n14), .A1(
        oc8051_decoder1_n23), .B0(oc8051_decoder1_n11), .Y(
        oc8051_decoder1_n174) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u91 ( .A0(oc8051_decoder1_n6), .A1(
        oc8051_decoder1_n137), .A2(oc8051_decoder1_n53), .B0(
        oc8051_decoder1_n75), .B1(oc8051_decoder1_n174), .Y(
        oc8051_decoder1_n173) );
  INV_X0P5B_A12TS oc8051_decoder1_u90 ( .A(oc8051_decoder1_n173), .Y(
        oc8051_decoder1_n172) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u89 ( .A0(oc8051_decoder1_n147), .A1(
        oc8051_decoder1_n146), .B0(oc8051_decoder1_n171), .C0(
        oc8051_decoder1_n172), .Y(oc8051_decoder1_n170) );
  INV_X0P5B_A12TS oc8051_decoder1_u88 ( .A(oc8051_decoder1_n170), .Y(
        oc8051_decoder1_n169) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u87 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n169), .B0(oc8051_decoder1_alu_op_2_), .B1(wait_data), 
        .Y(oc8051_decoder1_n168) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u86 ( .A0(oc8051_decoder1_n166), .A1(
        oc8051_decoder1_n151), .B0(oc8051_decoder1_n167), .C0(
        oc8051_decoder1_n168), .Y(oc8051_decoder1_n422) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u85 ( .A(oc8051_decoder1_n137), .B(
        oc8051_decoder1_n82), .S0(oc8051_decoder1_n14), .Y(
        oc8051_decoder1_n159) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u84 ( .A0(oc8051_decoder1_n156), .A1(
        oc8051_decoder1_n54), .B0(oc8051_decoder1_n165), .Y(
        oc8051_decoder1_n162) );
  INV_X0P5B_A12TS oc8051_decoder1_u83 ( .A(oc8051_decoder1_n164), .Y(
        oc8051_decoder1_n163) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u82 ( .A(oc8051_decoder1_n161), .B(
        oc8051_decoder1_n162), .S0(oc8051_decoder1_n163), .Y(
        oc8051_decoder1_n160) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u81 ( .A0(oc8051_decoder1_n141), .A1(
        oc8051_decoder1_n75), .A2(oc8051_decoder1_n159), .B0(
        oc8051_decoder1_n160), .B1(oc8051_decoder1_n41), .Y(
        oc8051_decoder1_n158) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u80 ( .A0(oc8051_decoder1_n58), .A1(
        oc8051_decoder1_n157), .A2(oc8051_decoder1_n50), .B0(
        oc8051_decoder1_n158), .Y(oc8051_decoder1_n148) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u79 ( .A0(oc8051_decoder1_n47), .A1(
        oc8051_decoder1_n155), .B0(oc8051_decoder1_n156), .B1(
        oc8051_decoder1_n132), .Y(oc8051_decoder1_n153) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u78 ( .A0(oc8051_decoder1_n153), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n154), .B1(
        oc8051_decoder1_n40), .Y(oc8051_decoder1_n152) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u77 ( .A0(oc8051_decoder1_n150), .A1(
        oc8051_decoder1_n151), .A2(oc8051_decoder1_n152), .B0(
        oc8051_decoder1_n37), .Y(oc8051_decoder1_n149) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u76 ( .A0(oc8051_decoder1_n146), .A1(
        oc8051_decoder1_n147), .B0(oc8051_decoder1_n148), .C0(
        oc8051_decoder1_n149), .Y(oc8051_decoder1_n143) );
  OAI222_X0P5M_A12TS oc8051_decoder1_u75 ( .A0(oc8051_decoder1_n123), .A1(
        oc8051_decoder1_n122), .B0(oc8051_decoder1_n143), .B1(
        oc8051_decoder1_n144), .C0(oc8051_decoder1_n125), .C1(
        oc8051_decoder1_n145), .Y(oc8051_decoder1_n423) );
  AOI221_X0P5M_A12TS oc8051_decoder1_u74 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n58), .B0(oc8051_decoder1_n138), .B1(op1_cur[0]), .C0(
        oc8051_decoder1_n142), .Y(oc8051_decoder1_n140) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u73 ( .A0(oc8051_decoder1_n139), .A1(
        op1_cur[1]), .B0(oc8051_decoder1_n140), .C0(oc8051_decoder1_n141), .Y(
        oc8051_decoder1_n129) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u72 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n137), .B0(oc8051_decoder1_n138), .Y(
        oc8051_decoder1_n133) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u71 ( .A0(oc8051_decoder1_n135), .A1(
        oc8051_decoder1_n136), .B0(oc8051_decoder1_n42), .B1(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n134) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u70 ( .A(oc8051_decoder1_n132), .B(
        op1_cur[1]), .C(oc8051_decoder1_n133), .D(oc8051_decoder1_n134), .Y(
        oc8051_decoder1_n130) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u69 ( .A(oc8051_decoder1_n129), .B(
        oc8051_decoder1_n130), .S0(oc8051_decoder1_n131), .Y(
        oc8051_decoder1_n127) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u68 ( .A0(oc8051_decoder1_n126), .A1(
        oc8051_decoder1_n69), .A2(oc8051_decoder1_n127), .B0(
        oc8051_decoder1_n128), .Y(oc8051_decoder1_n120) );
  OA22_X0P5M_A12TS oc8051_decoder1_u67 ( .A0(oc8051_decoder1_n122), .A1(
        oc8051_decoder1_n123), .B0(oc8051_decoder1_n124), .B1(
        oc8051_decoder1_n125), .Y(oc8051_decoder1_n121) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u66 ( .A0(oc8051_decoder1_n118), .A1(
        oc8051_decoder1_n119), .B0(oc8051_decoder1_n120), .C0(
        oc8051_decoder1_n121), .Y(oc8051_decoder1_n424) );
  INV_X0P5B_A12TS oc8051_decoder1_u65 ( .A(wb_rst_i), .Y(oc8051_decoder1_n444)
         );
  NAND2_X0P5A_A12TS oc8051_decoder1_u64 ( .A(oc8051_decoder1_n117), .B(
        oc8051_decoder1_n33), .Y(oc8051_decoder1_n106) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u63 ( .A(oc8051_decoder1_n115), .B(
        oc8051_decoder1_n116), .Y(oc8051_decoder1_n72) );
  NAND3B_X0P5M_A12TS oc8051_decoder1_u62 ( .AN(oc8051_decoder1_n72), .B(
        oc8051_decoder1_n113), .C(oc8051_decoder1_n114), .Y(
        oc8051_decoder1_n96) );
  INV_X0P5B_A12TS oc8051_decoder1_u61 ( .A(oc8051_decoder1_n112), .Y(
        oc8051_decoder1_n94) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u60 ( .A0(oc8051_decoder1_n96), .A1(
        oc8051_decoder1_n94), .B0(oc8051_decoder1_n111), .Y(
        oc8051_decoder1_n107) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u59 ( .A(oc8051_decoder1_n68), .B(
        oc8051_decoder1_n75), .C(oc8051_decoder1_n110), .Y(oc8051_decoder1_n34) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u58 ( .A(oc8051_decoder1_n108), .B(
        oc8051_decoder1_n33), .C(oc8051_decoder1_n109), .Y(oc8051_decoder1_n89) );
  NAND4_X0P5A_A12TS oc8051_decoder1_u57 ( .A(oc8051_decoder1_n106), .B(
        oc8051_decoder1_n107), .C(oc8051_decoder1_n34), .D(oc8051_decoder1_n89), .Y(pc_wr_sel[0]) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u56 ( .A(oc8051_decoder1_n59), .B(
        oc8051_decoder1_n105), .Y(oc8051_decoder1_n7) );
  INV_X0P5B_A12TS oc8051_decoder1_u55 ( .A(oc8051_decoder1_n104), .Y(
        oc8051_decoder1_n103) );
  NAND2_X0P5A_A12TS oc8051_decoder1_u54 ( .A(oc8051_decoder1_n103), .B(
        oc8051_decoder1_n75), .Y(oc8051_decoder1_n87) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u53 ( .A0(oc8051_decoder1_n7), .A1(
        oc8051_decoder1_n14), .A2(oc8051_decoder1_n102), .B0(
        oc8051_decoder1_n87), .Y(oc8051_decoder1_n63) );
  INV_X0P5B_A12TS oc8051_decoder1_u52 ( .A(oc8051_decoder1_n63), .Y(
        oc8051_decoder1_n100) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u51 ( .A0(oc8051_decoder1_n5), .A1(
        oc8051_decoder1_n100), .B0(oc8051_decoder1_n29), .B1(
        oc8051_decoder1_n30), .C0(oc8051_decoder1_n101), .Y(
        oc8051_decoder1_n441) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u50 ( .A(oc8051_decoder1_n78), .B(
        oc8051_decoder1_n87), .C(oc8051_decoder1_n29), .Y(oc8051_decoder1_n93)
         );
  OAI21_X0P5M_A12TS oc8051_decoder1_u49 ( .A0(oc8051_decoder1_n98), .A1(
        oc8051_decoder1_n69), .B0(oc8051_decoder1_n99), .Y(oc8051_decoder1_n97) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u48 ( .A0(oc8051_decoder1_n53), .A1(
        oc8051_decoder1_n81), .B0(oc8051_decoder1_n96), .C0(
        oc8051_decoder1_n97), .Y(oc8051_decoder1_n95) );
  INV_X0P5B_A12TS oc8051_decoder1_u47 ( .A(oc8051_decoder1_n95), .Y(
        oc8051_decoder1_n86) );
  NOR3_X0P5A_A12TS oc8051_decoder1_u46 ( .A(oc8051_decoder1_n93), .B(
        oc8051_decoder1_n86), .C(oc8051_decoder1_n94), .Y(oc8051_decoder1_n91)
         );
  OAI22_X0P5M_A12TS oc8051_decoder1_u45 ( .A0(oc8051_decoder1_n91), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n5), .B1(oc8051_decoder1_n92), .Y(pc_wr_sel[1]) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u44 ( .A(oc8051_decoder1_n90), .B(
        oc8051_decoder1_n33), .C(oc8051_decoder1_n44), .Y(oc8051_decoder1_n88)
         );
  OAI211_X0P5M_A12TS oc8051_decoder1_u43 ( .A0(oc8051_decoder1_n30), .A1(
        oc8051_decoder1_n87), .B0(oc8051_decoder1_n88), .C0(
        oc8051_decoder1_n89), .Y(pc_wr_sel[2]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u42 ( .A(oc8051_decoder1_n85), .B(
        oc8051_decoder1_n86), .Y(oc8051_decoder1_n79) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u41 ( .A0(oc8051_decoder1_n81), .A1(
        oc8051_decoder1_n82), .B0(oc8051_decoder1_n83), .C0(
        oc8051_decoder1_n84), .Y(oc8051_decoder1_n80) );
  MXIT2_X0P5M_A12TS oc8051_decoder1_u40 ( .A(oc8051_decoder1_n79), .B(
        oc8051_decoder1_n80), .S0(eq), .Y(oc8051_decoder1_n76) );
  INV_X0P5B_A12TS oc8051_decoder1_u39 ( .A(oc8051_decoder1_n78), .Y(
        oc8051_decoder1_n77) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u38 ( .A0(oc8051_decoder1_n68), .A1(
        oc8051_decoder1_n75), .B0(oc8051_decoder1_n76), .C0(
        oc8051_decoder1_n77), .Y(oc8051_decoder1_n73) );
  INV_X0P5B_A12TS oc8051_decoder1_u37 ( .A(pc_wr_sel[2]), .Y(
        oc8051_decoder1_n74) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u36 ( .A0(oc8051_decoder1_n73), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n34), .C0(
        oc8051_decoder1_n74), .Y(pc_wr) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u35 ( .A0(oc8051_decoder1_n70), .A1(
        oc8051_decoder1_n71), .B0(oc8051_decoder1_n67), .C0(
        oc8051_decoder1_n72), .Y(oc8051_decoder1_n64) );
  AOI22_X0P5M_A12TS oc8051_decoder1_u34 ( .A0(oc8051_decoder1_n67), .A1(
        oc8051_decoder1_n21), .B0(oc8051_decoder1_n68), .B1(
        oc8051_decoder1_n69), .Y(oc8051_decoder1_n65) );
  OAI22_X0P5M_A12TS oc8051_decoder1_u33 ( .A0(oc8051_decoder1_n22), .A1(
        oc8051_decoder1_n64), .B0(oc8051_decoder1_n65), .B1(
        oc8051_decoder1_n66), .Y(oc8051_decoder1_n62) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u32 ( .A0(oc8051_decoder1_n60), .A1(
        oc8051_decoder1_n61), .B0(oc8051_decoder1_n62), .C0(
        oc8051_decoder1_n63), .Y(oc8051_decoder1_n56) );
  AO21_X0P5M_A12TS oc8051_decoder1_u31 ( .A0(oc8051_decoder1_n58), .A1(
        oc8051_decoder1_n59), .B0(comp_sel[0]), .Y(oc8051_decoder1_n57) );
  OAI211_X0P5M_A12TS oc8051_decoder1_u30 ( .A0(oc8051_decoder1_n5), .A1(
        oc8051_decoder1_n56), .B0(oc8051_decoder1_n57), .C0(
        oc8051_decoder1_n34), .Y(oc8051_decoder1_ram_rd_sel_0_) );
  AO21A1AI2_X0P5M_A12TS oc8051_decoder1_u29 ( .A0(oc8051_decoder1_n53), .A1(
        op1_cur[0]), .B0(oc8051_decoder1_n54), .C0(oc8051_decoder1_n55), .Y(
        oc8051_decoder1_n15) );
  INV_X0P5B_A12TS oc8051_decoder1_u28 ( .A(oc8051_decoder1_n15), .Y(
        oc8051_decoder1_n51) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u27 ( .A0(oc8051_decoder1_n21), .A1(
        oc8051_decoder1_n22), .A2(oc8051_decoder1_n51), .B0(
        oc8051_decoder1_n52), .Y(oc8051_decoder1_n45) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u26 ( .A0(oc8051_decoder1_n47), .A1(
        oc8051_decoder1_n48), .B0(oc8051_decoder1_n49), .C0(
        oc8051_decoder1_n50), .Y(oc8051_decoder1_n46) );
  AOI211_X0P5M_A12TS oc8051_decoder1_u25 ( .A0(oc8051_decoder1_n8), .A1(
        oc8051_decoder1_n40), .B0(oc8051_decoder1_n45), .C0(
        oc8051_decoder1_n46), .Y(oc8051_decoder1_n35) );
  OA21A1OI2_X0P5M_A12TS oc8051_decoder1_u24 ( .A0(oc8051_decoder1_n42), .A1(
        oc8051_decoder1_n26), .B0(oc8051_decoder1_n27), .C0(
        oc8051_decoder1_n14), .Y(oc8051_decoder1_n43) );
  AOI32_X0P5M_A12TS oc8051_decoder1_u23 ( .A0(oc8051_decoder1_n40), .A1(
        oc8051_decoder1_n41), .A2(oc8051_decoder1_n42), .B0(
        oc8051_decoder1_n43), .B1(oc8051_decoder1_n44), .Y(oc8051_decoder1_n39) );
  OAI221_X0P5M_A12TS oc8051_decoder1_u22 ( .A0(oc8051_decoder1_n35), .A1(
        oc8051_decoder1_n36), .B0(oc8051_decoder1_n37), .B1(
        oc8051_decoder1_n38), .C0(oc8051_decoder1_n39), .Y(oc8051_decoder1_n32) );
  AOI21B_X0P5M_A12TS oc8051_decoder1_u21 ( .A0(oc8051_decoder1_n32), .A1(
        oc8051_decoder1_n33), .B0N(oc8051_decoder1_n34), .Y(
        oc8051_decoder1_n31) );
  OAI21_X0P5M_A12TS oc8051_decoder1_u20 ( .A0(oc8051_decoder1_n29), .A1(
        oc8051_decoder1_n30), .B0(oc8051_decoder1_n31), .Y(
        oc8051_decoder1_ram_rd_sel_1_) );
  MXT2_X0P5M_A12TS oc8051_decoder1_u19 ( .A(oc8051_decoder1_ram_rd_sel_0_), 
        .B(oc8051_decoder1_ram_rd_sel_r[0]), .S0(wait_data), .Y(ram_rd_sel[0])
         );
  MXT2_X0P5M_A12TS oc8051_decoder1_u18 ( .A(oc8051_decoder1_ram_rd_sel_1_), 
        .B(oc8051_decoder1_ram_rd_sel_r[1]), .S0(wait_data), .Y(ram_rd_sel[1])
         );
  MXT2_X0P5M_A12TS oc8051_decoder1_u17 ( .A(oc8051_decoder1_n441), .B(
        oc8051_decoder1_ram_rd_sel_r[2]), .S0(wait_data), .Y(ram_rd_sel[2]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u16 ( .A(wait_data), .B(oc8051_decoder1_n28), .Y(ram_wr_sel[0]) );
  NOR2B_X0P5M_A12TS oc8051_decoder1_u15 ( .AN(oc8051_decoder1_ram_wr_sel_1_), 
        .B(wait_data), .Y(ram_wr_sel[1]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u14 ( .A(wait_data), .B(
        oc8051_decoder1_n408), .Y(ram_wr_sel[2]) );
  OAI31_X0P5M_A12TS oc8051_decoder1_u13 ( .A0(oc8051_decoder1_n25), .A1(
        oc8051_decoder1_n26), .A2(oc8051_decoder1_n11), .B0(
        oc8051_decoder1_n27), .Y(oc8051_decoder1_n17) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u12 ( .A0(oc8051_decoder1_n21), .A1(
        oc8051_decoder1_n22), .A2(oc8051_decoder1_n23), .B0(
        oc8051_decoder1_n24), .Y(oc8051_decoder1_n19) );
  AOI31_X0P5M_A12TS oc8051_decoder1_u11 ( .A0(oc8051_decoder1_n17), .A1(
        oc8051_decoder1_n18), .A2(oc8051_decoder1_n19), .B0(
        oc8051_decoder1_n20), .Y(oc8051_decoder1_n2) );
  NAND3_X0P5A_A12TS oc8051_decoder1_u10 ( .A(oc8051_decoder1_n14), .B(
        oc8051_decoder1_n15), .C(oc8051_decoder1_n16), .Y(oc8051_decoder1_n3)
         );
  NAND3_X0P5A_A12TS oc8051_decoder1_u9 ( .A(oc8051_decoder1_n11), .B(
        oc8051_decoder1_n12), .C(oc8051_decoder1_n13), .Y(oc8051_decoder1_n10)
         );
  AOI32_X0P5M_A12TS oc8051_decoder1_u8 ( .A0(oc8051_decoder1_n6), .A1(
        oc8051_decoder1_n7), .A2(oc8051_decoder1_n8), .B0(oc8051_decoder1_n9), 
        .B1(oc8051_decoder1_n10), .Y(oc8051_decoder1_n4) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u7 ( .A(wait_data), .B(oc8051_decoder1_n1), 
        .Y(wr_o) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u6 ( .A(wait_data), .B(oc8051_decoder1_n407), .Y(wr_sfr[0]) );
  NOR2_X0P5A_A12TS oc8051_decoder1_u5 ( .A(wait_data), .B(oc8051_decoder1_n406), .Y(wr_sfr[1]) );
  OAI22_X1M_A12TS oc8051_decoder1_u4 ( .A0(oc8051_decoder1_n318), .A1(
        oc8051_decoder1_n301), .B0(oc8051_decoder1_n439), .B1(
        oc8051_decoder1_n302), .Y(op1_cur[0]) );
  AOI31_X2M_A12TS oc8051_decoder1_u3 ( .A0(oc8051_decoder1_n2), .A1(
        oc8051_decoder1_n3), .A2(oc8051_decoder1_n4), .B0(oc8051_decoder1_n5), 
        .Y(rmw) );
  DFFRPQN_X1M_A12TS oc8051_decoder1_ram_wr_sel_reg_2_ ( .D(
        oc8051_decoder1_n412), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_decoder1_n408) );
  DFFRPQN_X1M_A12TS oc8051_decoder1_wr_sfr_reg_0_ ( .D(oc8051_decoder1_n414), 
        .CK(wb_clk_i), .R(wb_rst_i), .QN(oc8051_decoder1_n407) );
  DFFRPQN_X1M_A12TS oc8051_decoder1_wr_sfr_reg_1_ ( .D(oc8051_decoder1_n413), 
        .CK(wb_clk_i), .R(wb_rst_i), .QN(oc8051_decoder1_n406) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel3_reg ( .D(oc8051_decoder1_n394), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel3) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel1_reg_0_ ( .D(oc8051_decoder1_n417), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel1[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel1_reg_1_ ( .D(oc8051_decoder1_n416), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel1[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel1_reg_2_ ( .D(oc8051_decoder1_n415), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel1[2]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_psw_set_reg_1_ ( .D(oc8051_decoder1_n420), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(psw_set[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel2_reg_0_ ( .D(oc8051_decoder1_n390), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel2[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_src_sel2_reg_1_ ( .D(oc8051_decoder1_n392), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(src_sel2[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_psw_set_reg_0_ ( .D(oc8051_decoder1_n389), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(psw_set[0]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_state_reg_0_ ( .D(oc8051_decoder1_n405), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(oc8051_decoder1_state_0_)
         );
  DFFRPQ_X1M_A12TS oc8051_decoder1_cy_sel_reg_0_ ( .D(oc8051_decoder1_n391), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(cy_sel[0]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_state_reg_1_ ( .D(oc8051_decoder1_n395), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(oc8051_decoder1_state_1_)
         );
  DFFRPQ_X1M_A12TS oc8051_decoder1_cy_sel_reg_1_ ( .D(oc8051_decoder1_n393), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(cy_sel[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_wr_sel_reg_1_ ( .D(oc8051_decoder1_n418), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_ram_wr_sel_1_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_2_ ( .D(oc8051_decoder1_n422), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_2_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_3_ ( .D(oc8051_decoder1_n388), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_3_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_0_ ( .D(oc8051_decoder1_n424), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_0_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_alu_op_reg_1_ ( .D(oc8051_decoder1_n423), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_alu_op_1_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_wr_reg ( .D(oc8051_decoder1_n421), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_wr) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_wr_sel_reg_0_ ( .D(oc8051_decoder1_n419), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_ram_wr_sel_0_) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_7_ ( .D(oc8051_decoder1_n396), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[7]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_6_ ( .D(oc8051_decoder1_n397), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[6]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_5_ ( .D(oc8051_decoder1_n398), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[5]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_4_ ( .D(oc8051_decoder1_n399), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[4]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_3_ ( .D(oc8051_decoder1_n400), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[3]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_2_ ( .D(oc8051_decoder1_n401), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[2]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_1_ ( .D(oc8051_decoder1_n402), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_op_reg_0_ ( .D(oc8051_decoder1_n403), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_decoder1_op[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_rd_sel_r_reg_0_ ( .D(
        oc8051_decoder1_ram_rd_sel_0_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_decoder1_ram_rd_sel_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_rd_sel_r_reg_1_ ( .D(
        oc8051_decoder1_ram_rd_sel_1_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_decoder1_ram_rd_sel_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_decoder1_ram_rd_sel_r_reg_2_ ( .D(
        oc8051_decoder1_n441), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_decoder1_ram_rd_sel_r[2]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_mem_act_reg_1_ ( .D(oc8051_decoder1_n1805), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(mem_act[1]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_mem_act_reg_0_ ( .D(oc8051_decoder1_n1804), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(mem_act[0]) );
  DFFSQ_X1M_A12TS oc8051_decoder1_mem_act_reg_2_ ( .D(oc8051_decoder1_n1806), 
        .CK(wb_clk_i), .SN(oc8051_decoder1_n444), .Q(mem_act[2]) );
  INV_X0P5B_A12TS oc8051_alu1_u332 ( .A(alu_op[2]), .Y(oc8051_alu1_n281) );
  NOR2_X0P5A_A12TS oc8051_alu1_u331 ( .A(oc8051_alu1_n281), .B(alu_op[3]), .Y(
        oc8051_alu1_n277) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u330 ( .AN(alu_op[0]), .B(alu_op[1]), .Y(
        oc8051_alu1_n269) );
  NAND2_X0P5A_A12TS oc8051_alu1_u329 ( .A(oc8051_alu1_n277), .B(
        oc8051_alu1_n269), .Y(oc8051_alu1_n47) );
  INV_X0P5B_A12TS oc8051_alu1_u328 ( .A(oc8051_alu1_n47), .Y(oc8051_alu1_n41)
         );
  INV_X0P5B_A12TS oc8051_alu1_u327 ( .A(src1[3]), .Y(oc8051_alu1_n4) );
  NOR2_X0P5A_A12TS oc8051_alu1_u326 ( .A(src1[2]), .B(src1[1]), .Y(
        oc8051_alu1_n227) );
  NOR2_X0P5A_A12TS oc8051_alu1_u325 ( .A(oc8051_alu1_n4), .B(oc8051_alu1_n227), 
        .Y(oc8051_alu1_n180) );
  INV_X0P5B_A12TS oc8051_alu1_u324 ( .A(oc8051_alu1_n180), .Y(oc8051_alu1_n29)
         );
  NAND2B_X0P5M_A12TS oc8051_alu1_u323 ( .AN(srcac), .B(oc8051_alu1_n29), .Y(
        oc8051_alu1_n283) );
  NAND2_X0P5A_A12TS oc8051_alu1_u322 ( .A(oc8051_alu1_n41), .B(
        oc8051_alu1_n283), .Y(oc8051_alu1_n30) );
  NOR2_X0P5A_A12TS oc8051_alu1_u321 ( .A(alu_op[1]), .B(alu_op[0]), .Y(
        oc8051_alu1_n270) );
  NOR2_X0P5A_A12TS oc8051_alu1_u320 ( .A(alu_op[3]), .B(alu_op[2]), .Y(
        oc8051_alu1_n272) );
  NAND2_X0P5A_A12TS oc8051_alu1_u319 ( .A(oc8051_alu1_n270), .B(
        oc8051_alu1_n272), .Y(oc8051_alu1_n35) );
  OAI21_X0P5M_A12TS oc8051_alu1_u318 ( .A0(oc8051_alu1_n47), .A1(
        oc8051_alu1_n283), .B0(oc8051_alu1_n35), .Y(oc8051_alu1_n261) );
  INV_X0P5B_A12TS oc8051_alu1_u317 ( .A(oc8051_alu1_n261), .Y(oc8051_alu1_n225) );
  INV_X0P5B_A12TS oc8051_alu1_u316 ( .A(src1[0]), .Y(oc8051_alu1_n27) );
  NAND2_X0P5A_A12TS oc8051_alu1_u315 ( .A(oc8051_alu1_n269), .B(
        oc8051_alu1_n272), .Y(oc8051_alu1_n111) );
  INV_X0P5B_A12TS oc8051_alu1_u314 ( .A(oc8051_alu1_n111), .Y(oc8051_alu1_n289) );
  INV_X0P5B_A12TS oc8051_alu1_u313 ( .A(alu_op[1]), .Y(oc8051_alu1_n278) );
  NOR2_X0P5A_A12TS oc8051_alu1_u312 ( .A(oc8051_alu1_n278), .B(alu_op[0]), .Y(
        oc8051_alu1_n267) );
  NAND2_X0P5A_A12TS oc8051_alu1_u311 ( .A(oc8051_alu1_n267), .B(
        oc8051_alu1_n272), .Y(oc8051_alu1_n11) );
  INV_X0P5B_A12TS oc8051_alu1_u310 ( .A(oc8051_alu1_n11), .Y(oc8051_alu1_n24)
         );
  INV_X0P5B_A12TS oc8051_alu1_u309 ( .A(alu_cy), .Y(oc8051_alu1_n133) );
  XOR2_X0P5M_A12TS oc8051_alu1_u308 ( .A(src2[0]), .B(src1[0]), .Y(
        oc8051_alu1_n275) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u307 ( .A(oc8051_alu1_n133), .B(
        oc8051_alu1_n275), .Y(sub_result[0]) );
  OAI21_X0P5M_A12TS oc8051_alu1_u306 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n24), .B0(sub_result[0]), .Y(oc8051_alu1_n282) );
  AO21A1AI2_X0P5M_A12TS oc8051_alu1_u305 ( .A0(oc8051_alu1_n30), .A1(
        oc8051_alu1_n225), .B0(oc8051_alu1_n27), .C0(oc8051_alu1_n282), .Y(
        oc8051_alu1_n262) );
  NAND2_X0P5A_A12TS oc8051_alu1_u304 ( .A(oc8051_alu1_n270), .B(
        oc8051_alu1_n277), .Y(oc8051_alu1_n128) );
  INV_X0P5B_A12TS oc8051_alu1_u303 ( .A(oc8051_alu1_n128), .Y(oc8051_alu1_n288) );
  INV_X0P5B_A12TS oc8051_alu1_u302 ( .A(alu_op[3]), .Y(oc8051_alu1_n280) );
  NOR2_X0P5A_A12TS oc8051_alu1_u301 ( .A(oc8051_alu1_n280), .B(
        oc8051_alu1_n281), .Y(oc8051_alu1_n268) );
  AND3_X0P5M_A12TS oc8051_alu1_u300 ( .A(oc8051_alu1_n268), .B(alu_cy), .C(
        oc8051_alu1_n267), .Y(oc8051_alu1_n67) );
  NAND2_X0P5A_A12TS oc8051_alu1_u299 ( .A(oc8051_alu1_n267), .B(
        oc8051_alu1_n277), .Y(oc8051_alu1_n50) );
  NOR2_X0P5A_A12TS oc8051_alu1_u298 ( .A(oc8051_alu1_n280), .B(alu_op[2]), .Y(
        oc8051_alu1_n266) );
  NAND2_X0P5A_A12TS oc8051_alu1_u297 ( .A(oc8051_alu1_n266), .B(
        oc8051_alu1_n269), .Y(oc8051_alu1_n36) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u296 ( .A(oc8051_alu1_n50), .B(oc8051_alu1_n36), .S0(src1[0]), .Y(oc8051_alu1_n279) );
  AOI21_X0P5M_A12TS oc8051_alu1_u295 ( .A0(oc8051_alu1_dec[0]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_n279), .Y(oc8051_alu1_n273) );
  AND3_X0P5M_A12TS oc8051_alu1_u294 ( .A(oc8051_alu1_n268), .B(
        oc8051_alu1_n133), .C(oc8051_alu1_n267), .Y(oc8051_alu1_n66) );
  NAND2_X0P5A_A12TS oc8051_alu1_u293 ( .A(oc8051_alu1_n266), .B(
        oc8051_alu1_n270), .Y(oc8051_alu1_n48) );
  INV_X0P5B_A12TS oc8051_alu1_u292 ( .A(oc8051_alu1_n48), .Y(oc8051_alu1_n46)
         );
  NOR2B_X0P5M_A12TS oc8051_alu1_u291 ( .AN(alu_op[0]), .B(oc8051_alu1_n278), 
        .Y(oc8051_alu1_n271) );
  NAND2_X0P5A_A12TS oc8051_alu1_u290 ( .A(oc8051_alu1_n271), .B(
        oc8051_alu1_n277), .Y(oc8051_alu1_n44) );
  NAND2_X0P5A_A12TS oc8051_alu1_u289 ( .A(oc8051_alu1_n268), .B(
        oc8051_alu1_n271), .Y(oc8051_alu1_n204) );
  INV_X0P5B_A12TS oc8051_alu1_u288 ( .A(oc8051_alu1_n204), .Y(oc8051_alu1_n92)
         );
  NOR2B_X0P5M_A12TS oc8051_alu1_u287 ( .AN(oc8051_alu1_n36), .B(
        oc8051_alu1_n92), .Y(oc8051_alu1_n221) );
  INV_X0P5B_A12TS oc8051_alu1_u286 ( .A(src2[0]), .Y(oc8051_alu1_n256) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u285 ( .A0(oc8051_alu1_n27), .A1(
        oc8051_alu1_n44), .B0(oc8051_alu1_n221), .C0(oc8051_alu1_n256), .Y(
        oc8051_alu1_n276) );
  AOI221_X0P5M_A12TS oc8051_alu1_u284 ( .A0(oc8051_alu1_inc[0]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_n46), .B1(oc8051_alu1_n275), .C0(
        oc8051_alu1_n276), .Y(oc8051_alu1_n274) );
  NAND2_X0P5A_A12TS oc8051_alu1_u283 ( .A(oc8051_alu1_n273), .B(
        oc8051_alu1_n274), .Y(oc8051_alu1_n9) );
  AOI21_X0P5M_A12TS oc8051_alu1_u282 ( .A0(oc8051_alu1_divsrc1[0]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n9), .Y(oc8051_alu1_n263) );
  AND2_X0P5M_A12TS oc8051_alu1_u281 ( .A(oc8051_alu1_n266), .B(
        oc8051_alu1_n271), .Y(oc8051_alu1_n51) );
  NAND2_X0P5A_A12TS oc8051_alu1_u280 ( .A(oc8051_alu1_n271), .B(
        oc8051_alu1_n272), .Y(oc8051_alu1_n127) );
  INV_X0P5B_A12TS oc8051_alu1_u279 ( .A(oc8051_alu1_n127), .Y(oc8051_alu1_n290) );
  AOI22_X0P5M_A12TS oc8051_alu1_u278 ( .A0(oc8051_alu1_n51), .A1(alu_cy), .B0(
        oc8051_alu1_mulsrc1[0]), .B1(oc8051_alu1_n290), .Y(oc8051_alu1_n264)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_u277 ( .A(oc8051_alu1_n268), .B(
        oc8051_alu1_n270), .Y(oc8051_alu1_n134) );
  NAND2_X0P5A_A12TS oc8051_alu1_u276 ( .A(oc8051_alu1_n268), .B(
        oc8051_alu1_n269), .Y(oc8051_alu1_n28) );
  NAND2_X0P5A_A12TS oc8051_alu1_u275 ( .A(oc8051_alu1_n134), .B(
        oc8051_alu1_n28), .Y(oc8051_alu1_n124) );
  NAND2_X0P5A_A12TS oc8051_alu1_u274 ( .A(oc8051_alu1_n266), .B(
        oc8051_alu1_n267), .Y(oc8051_alu1_n37) );
  INV_X0P5B_A12TS oc8051_alu1_u273 ( .A(oc8051_alu1_n37), .Y(oc8051_alu1_n254)
         );
  AOI22_X0P5M_A12TS oc8051_alu1_u272 ( .A0(src1[1]), .A1(oc8051_alu1_n124), 
        .B0(oc8051_alu1_n254), .B1(src1[7]), .Y(oc8051_alu1_n265) );
  NAND4B_X0P5M_A12TS oc8051_alu1_u271 ( .AN(oc8051_alu1_n262), .B(
        oc8051_alu1_n263), .C(oc8051_alu1_n264), .D(oc8051_alu1_n265), .Y(
        oc8051_alu1_n2130) );
  INV_X0P5B_A12TS oc8051_alu1_u270 ( .A(oc8051_alu1_n30), .Y(oc8051_alu1_n235)
         );
  MXIT2_X0P5M_A12TS oc8051_alu1_u269 ( .A(oc8051_alu1_n235), .B(
        oc8051_alu1_n261), .S0(src1[1]), .Y(oc8051_alu1_n248) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u268 ( .A(oc8051_alu1_n50), .B(oc8051_alu1_n36), .S0(src1[1]), .Y(oc8051_alu1_n260) );
  AOI21_X0P5M_A12TS oc8051_alu1_u267 ( .A0(oc8051_alu1_dec[1]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_n260), .Y(oc8051_alu1_n257) );
  XOR2_X0P5M_A12TS oc8051_alu1_u266 ( .A(src2[1]), .B(src1[1]), .Y(
        oc8051_alu1_n253) );
  INV_X0P5B_A12TS oc8051_alu1_u265 ( .A(src1[1]), .Y(oc8051_alu1_n8) );
  INV_X0P5B_A12TS oc8051_alu1_u264 ( .A(src2[1]), .Y(oc8051_alu1_n239) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u263 ( .A0(oc8051_alu1_n8), .A1(
        oc8051_alu1_n44), .B0(oc8051_alu1_n221), .C0(oc8051_alu1_n239), .Y(
        oc8051_alu1_n259) );
  AOI221_X0P5M_A12TS oc8051_alu1_u262 ( .A0(oc8051_alu1_inc[1]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_n46), .B1(oc8051_alu1_n253), .C0(
        oc8051_alu1_n259), .Y(oc8051_alu1_n258) );
  AND2_X0P5M_A12TS oc8051_alu1_u261 ( .A(oc8051_alu1_n257), .B(
        oc8051_alu1_n258), .Y(oc8051_alu1_n7) );
  NOR2_X0P5A_A12TS oc8051_alu1_u260 ( .A(src1[0]), .B(oc8051_alu1_n256), .Y(
        oc8051_alu1_n255) );
  OAI22_X0P5M_A12TS oc8051_alu1_u259 ( .A0(src2[0]), .A1(oc8051_alu1_n27), 
        .B0(alu_cy), .B1(oc8051_alu1_n255), .Y(oc8051_alu1_n246) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u258 ( .A(oc8051_alu1_n246), .B(
        oc8051_alu1_n253), .Y(sub_result[1]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u257 ( .A0(oc8051_alu1_divsrc1[1]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n24), .B1(sub_result[1]), .Y(
        oc8051_alu1_n249) );
  NOR2_X0P5A_A12TS oc8051_alu1_u256 ( .A(oc8051_alu1_n51), .B(oc8051_alu1_n254), .Y(oc8051_alu1_n126) );
  CGENI_X1M_A12TS oc8051_alu1_u255 ( .A(src1[0]), .B(alu_cy), .CI(src2[0]), 
        .CON(oc8051_alu1_n237) );
  XOR2_X0P5M_A12TS oc8051_alu1_u254 ( .A(oc8051_alu1_n237), .B(
        oc8051_alu1_n253), .Y(oc8051_alu1_n252) );
  OAI22_X0P5M_A12TS oc8051_alu1_u253 ( .A0(oc8051_alu1_n126), .A1(
        oc8051_alu1_n27), .B0(oc8051_alu1_n111), .B1(oc8051_alu1_n252), .Y(
        oc8051_alu1_n251) );
  AOI221_X0P5M_A12TS oc8051_alu1_u252 ( .A0(src1[2]), .A1(oc8051_alu1_n124), 
        .B0(oc8051_alu1_mulsrc1[1]), .B1(oc8051_alu1_n290), .C0(
        oc8051_alu1_n251), .Y(oc8051_alu1_n250) );
  NAND4_X0P5A_A12TS oc8051_alu1_u251 ( .A(oc8051_alu1_n248), .B(oc8051_alu1_n7), .C(oc8051_alu1_n249), .D(oc8051_alu1_n250), .Y(oc8051_alu1_n2140) );
  NAND2B_X0P5M_A12TS oc8051_alu1_u250 ( .AN(oc8051_alu1_n246), .B(
        oc8051_alu1_n8), .Y(oc8051_alu1_n247) );
  AOI22_X0P5M_A12TS oc8051_alu1_u249 ( .A0(oc8051_alu1_n246), .A1(src1[1]), 
        .B0(oc8051_alu1_n239), .B1(oc8051_alu1_n247), .Y(oc8051_alu1_n216) );
  XOR2_X0P5M_A12TS oc8051_alu1_u248 ( .A(src2[2]), .B(src1[2]), .Y(
        oc8051_alu1_n236) );
  XOR2_X0P5M_A12TS oc8051_alu1_u247 ( .A(oc8051_alu1_n216), .B(
        oc8051_alu1_n236), .Y(sub_result[2]) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u246 ( .A(oc8051_alu1_n50), .B(oc8051_alu1_n36), .S0(src1[2]), .Y(oc8051_alu1_n245) );
  AOI21_X0P5M_A12TS oc8051_alu1_u245 ( .A0(oc8051_alu1_dec[2]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_n245), .Y(oc8051_alu1_n241) );
  INV_X0P5B_A12TS oc8051_alu1_u244 ( .A(src1[2]), .Y(oc8051_alu1_n211) );
  INV_X0P5B_A12TS oc8051_alu1_u243 ( .A(src2[2]), .Y(oc8051_alu1_n244) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u242 ( .A0(oc8051_alu1_n211), .A1(
        oc8051_alu1_n44), .B0(oc8051_alu1_n221), .C0(oc8051_alu1_n244), .Y(
        oc8051_alu1_n243) );
  AOI221_X0P5M_A12TS oc8051_alu1_u241 ( .A0(oc8051_alu1_inc[2]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_n46), .B1(oc8051_alu1_n236), .C0(
        oc8051_alu1_n243), .Y(oc8051_alu1_n242) );
  NAND2_X0P5A_A12TS oc8051_alu1_u240 ( .A(oc8051_alu1_n241), .B(
        oc8051_alu1_n242), .Y(oc8051_alu1_n5) );
  AOI21_X0P5M_A12TS oc8051_alu1_u239 ( .A0(oc8051_alu1_n24), .A1(sub_result[2]), .B0(oc8051_alu1_n5), .Y(oc8051_alu1_n228) );
  AOI22_X0P5M_A12TS oc8051_alu1_u238 ( .A0(oc8051_alu1_mulsrc1[2]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc1[2]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n229) );
  INV_X0P5B_A12TS oc8051_alu1_u237 ( .A(oc8051_alu1_n126), .Y(oc8051_alu1_n165) );
  AOI22_X0P5M_A12TS oc8051_alu1_u236 ( .A0(src1[1]), .A1(oc8051_alu1_n165), 
        .B0(src1[3]), .B1(oc8051_alu1_n124), .Y(oc8051_alu1_n230) );
  INV_X0P5B_A12TS oc8051_alu1_u235 ( .A(oc8051_alu1_n237), .Y(oc8051_alu1_n240) );
  NOR2_X0P5A_A12TS oc8051_alu1_u234 ( .A(src1[1]), .B(oc8051_alu1_n240), .Y(
        oc8051_alu1_n238) );
  OAI22_X0P5M_A12TS oc8051_alu1_u233 ( .A0(oc8051_alu1_n237), .A1(
        oc8051_alu1_n8), .B0(oc8051_alu1_n238), .B1(oc8051_alu1_n239), .Y(
        oc8051_alu1_n214) );
  XOR2_X0P5M_A12TS oc8051_alu1_u232 ( .A(oc8051_alu1_n214), .B(
        oc8051_alu1_n236), .Y(oc8051_alu1_n232) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u231 ( .A0(oc8051_alu1_n8), .A1(
        oc8051_alu1_n30), .B0(oc8051_alu1_n225), .C0(oc8051_alu1_n211), .Y(
        oc8051_alu1_n233) );
  NAND2_X0P5A_A12TS oc8051_alu1_u230 ( .A(oc8051_alu1_n227), .B(
        oc8051_alu1_n235), .Y(oc8051_alu1_n226) );
  INV_X0P5B_A12TS oc8051_alu1_u229 ( .A(oc8051_alu1_n226), .Y(oc8051_alu1_n234) );
  AOI211_X0P5M_A12TS oc8051_alu1_u228 ( .A0(oc8051_alu1_n232), .A1(
        oc8051_alu1_n289), .B0(oc8051_alu1_n233), .C0(oc8051_alu1_n234), .Y(
        oc8051_alu1_n231) );
  NAND4_X0P5A_A12TS oc8051_alu1_u227 ( .A(oc8051_alu1_n228), .B(
        oc8051_alu1_n229), .C(oc8051_alu1_n230), .D(oc8051_alu1_n231), .Y(
        oc8051_alu1_n2150) );
  NOR2_X0P5A_A12TS oc8051_alu1_u226 ( .A(oc8051_alu1_n227), .B(oc8051_alu1_n30), .Y(oc8051_alu1_n223) );
  NAND2_X0P5A_A12TS oc8051_alu1_u225 ( .A(oc8051_alu1_n225), .B(
        oc8051_alu1_n226), .Y(oc8051_alu1_n224) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u224 ( .A(oc8051_alu1_n223), .B(
        oc8051_alu1_n224), .S0(src1[3]), .Y(oc8051_alu1_n207) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u223 ( .A(oc8051_alu1_n50), .B(oc8051_alu1_n36), .S0(src1[3]), .Y(oc8051_alu1_n222) );
  AOI21_X0P5M_A12TS oc8051_alu1_u222 ( .A0(oc8051_alu1_dec[3]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_n222), .Y(oc8051_alu1_n218) );
  INV_X0P5B_A12TS oc8051_alu1_u221 ( .A(src2[3]), .Y(oc8051_alu1_n197) );
  XOR2_X0P5M_A12TS oc8051_alu1_u220 ( .A(oc8051_alu1_n197), .B(oc8051_alu1_n4), 
        .Y(oc8051_alu1_n213) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u219 ( .A0(oc8051_alu1_n4), .A1(
        oc8051_alu1_n44), .B0(oc8051_alu1_n221), .C0(oc8051_alu1_n197), .Y(
        oc8051_alu1_n220) );
  AOI221_X0P5M_A12TS oc8051_alu1_u218 ( .A0(oc8051_alu1_inc[3]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_n46), .B1(oc8051_alu1_n213), .C0(
        oc8051_alu1_n220), .Y(oc8051_alu1_n219) );
  AND2_X0P5M_A12TS oc8051_alu1_u217 ( .A(oc8051_alu1_n218), .B(
        oc8051_alu1_n219), .Y(oc8051_alu1_n2) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u216 ( .AN(oc8051_alu1_n216), .B(src1[2]), .Y(
        oc8051_alu1_n217) );
  OAI22_X0P5M_A12TS oc8051_alu1_u215 ( .A0(oc8051_alu1_n216), .A1(
        oc8051_alu1_n211), .B0(src2[2]), .B1(oc8051_alu1_n217), .Y(
        oc8051_alu1_n198) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u214 ( .A(oc8051_alu1_n198), .B(
        oc8051_alu1_n213), .Y(sub_result[3]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u213 ( .A0(oc8051_alu1_divsrc1[3]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n24), .B1(sub_result[3]), .Y(
        oc8051_alu1_n208) );
  NAND2B_X0P5M_A12TS oc8051_alu1_u212 ( .AN(oc8051_alu1_n214), .B(
        oc8051_alu1_n211), .Y(oc8051_alu1_n215) );
  AOI22_X0P5M_A12TS oc8051_alu1_u211 ( .A0(oc8051_alu1_n214), .A1(src1[2]), 
        .B0(oc8051_alu1_n215), .B1(src2[2]), .Y(oc8051_alu1_n195) );
  XOR2_X0P5M_A12TS oc8051_alu1_u210 ( .A(oc8051_alu1_n195), .B(
        oc8051_alu1_n213), .Y(oc8051_alu1_n212) );
  OAI22_X0P5M_A12TS oc8051_alu1_u209 ( .A0(oc8051_alu1_n126), .A1(
        oc8051_alu1_n211), .B0(oc8051_alu1_n111), .B1(oc8051_alu1_n212), .Y(
        oc8051_alu1_n210) );
  AOI221_X0P5M_A12TS oc8051_alu1_u208 ( .A0(src1[4]), .A1(oc8051_alu1_n124), 
        .B0(oc8051_alu1_mulsrc1[3]), .B1(oc8051_alu1_n290), .C0(
        oc8051_alu1_n210), .Y(oc8051_alu1_n209) );
  NAND4_X0P5A_A12TS oc8051_alu1_u207 ( .A(oc8051_alu1_n207), .B(oc8051_alu1_n2), .C(oc8051_alu1_n208), .D(oc8051_alu1_n209), .Y(oc8051_alu1_n2160) );
  NOR2_X0P5A_A12TS oc8051_alu1_u206 ( .A(oc8051_alu1_n47), .B(oc8051_alu1_n29), 
        .Y(oc8051_alu1_n205) );
  NAND2_X0P5A_A12TS oc8051_alu1_u205 ( .A(oc8051_alu1_n92), .B(
        oc8051_alu1_n133), .Y(oc8051_alu1_n123) );
  NAND2_X0P5A_A12TS oc8051_alu1_u204 ( .A(oc8051_alu1_n35), .B(
        oc8051_alu1_n123), .Y(oc8051_alu1_n62) );
  NAND2B_X0P5M_A12TS oc8051_alu1_u203 ( .AN(oc8051_alu1_n62), .B(
        oc8051_alu1_n36), .Y(oc8051_alu1_n148) );
  OAI21B_X0P5M_A12TS oc8051_alu1_u202 ( .A0(oc8051_alu1_n180), .A1(
        oc8051_alu1_n47), .B0N(oc8051_alu1_n148), .Y(oc8051_alu1_n206) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u201 ( .A(oc8051_alu1_n205), .B(
        oc8051_alu1_n206), .S0(src1[4]), .Y(oc8051_alu1_n189) );
  INV_X0P5B_A12TS oc8051_alu1_u200 ( .A(src2[4]), .Y(oc8051_alu1_n188) );
  INV_X0P5B_A12TS oc8051_alu1_u199 ( .A(src1[4]), .Y(oc8051_alu1_n122) );
  NAND2_X0P5A_A12TS oc8051_alu1_u198 ( .A(src2[4]), .B(src1[4]), .Y(
        oc8051_alu1_n203) );
  INV_X0P5B_A12TS oc8051_alu1_u197 ( .A(oc8051_alu1_n203), .Y(oc8051_alu1_n183) );
  AOI21_X0P5M_A12TS oc8051_alu1_u196 ( .A0(oc8051_alu1_n188), .A1(
        oc8051_alu1_n122), .B0(oc8051_alu1_n183), .Y(oc8051_alu1_n194) );
  NOR2_X0P5A_A12TS oc8051_alu1_u195 ( .A(oc8051_alu1_n204), .B(
        oc8051_alu1_n133), .Y(oc8051_alu1_n65) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u194 ( .AN(oc8051_alu1_n36), .B(
        oc8051_alu1_n65), .Y(oc8051_alu1_n143) );
  OAI22_X0P5M_A12TS oc8051_alu1_u193 ( .A0(oc8051_alu1_n203), .A1(
        oc8051_alu1_n44), .B0(oc8051_alu1_n188), .B1(oc8051_alu1_n143), .Y(
        oc8051_alu1_n200) );
  INV_X0P5B_A12TS oc8051_alu1_u192 ( .A(oc8051_alu1_n50), .Y(oc8051_alu1_n170)
         );
  AOI222_X0P5M_A12TS oc8051_alu1_u191 ( .A0(oc8051_alu1_dec[4]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_inc[4]), .B1(oc8051_alu1_n66), .C0(
        oc8051_alu1_n170), .C1(oc8051_alu1_n122), .Y(oc8051_alu1_n202) );
  INV_X0P5B_A12TS oc8051_alu1_u190 ( .A(oc8051_alu1_n202), .Y(oc8051_alu1_n201) );
  AOI211_X0P5M_A12TS oc8051_alu1_u189 ( .A0(oc8051_alu1_n194), .A1(
        oc8051_alu1_n46), .B0(oc8051_alu1_n200), .C0(oc8051_alu1_n201), .Y(
        oc8051_alu1_n121) );
  NAND2B_X0P5M_A12TS oc8051_alu1_u188 ( .AN(oc8051_alu1_n198), .B(
        oc8051_alu1_n4), .Y(oc8051_alu1_n199) );
  AOI22_X0P5M_A12TS oc8051_alu1_u187 ( .A0(oc8051_alu1_n198), .A1(src1[3]), 
        .B0(oc8051_alu1_n197), .B1(oc8051_alu1_n199), .Y(oc8051_alu1_n55) );
  XOR2_X0P5M_A12TS oc8051_alu1_u186 ( .A(oc8051_alu1_n55), .B(oc8051_alu1_n194), .Y(sub_result[4]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u185 ( .A0(oc8051_alu1_divsrc1[4]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n24), .B1(sub_result[4]), .Y(
        oc8051_alu1_n190) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u184 ( .AN(oc8051_alu1_n195), .B(src1[3]), .Y(
        oc8051_alu1_n196) );
  OAI22_X0P5M_A12TS oc8051_alu1_u183 ( .A0(oc8051_alu1_n195), .A1(
        oc8051_alu1_n4), .B0(oc8051_alu1_n196), .B1(oc8051_alu1_n197), .Y(
        oc8051_alu1_n54) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u182 ( .A(oc8051_alu1_n194), .B(
        oc8051_alu1_n54), .Y(oc8051_alu1_n193) );
  OAI22_X0P5M_A12TS oc8051_alu1_u181 ( .A0(oc8051_alu1_n126), .A1(
        oc8051_alu1_n4), .B0(oc8051_alu1_n111), .B1(oc8051_alu1_n193), .Y(
        oc8051_alu1_n192) );
  AOI221_X0P5M_A12TS oc8051_alu1_u180 ( .A0(src1[5]), .A1(oc8051_alu1_n124), 
        .B0(oc8051_alu1_mulsrc1[4]), .B1(oc8051_alu1_n290), .C0(
        oc8051_alu1_n192), .Y(oc8051_alu1_n191) );
  NAND4_X0P5A_A12TS oc8051_alu1_u179 ( .A(oc8051_alu1_n189), .B(
        oc8051_alu1_n121), .C(oc8051_alu1_n190), .D(oc8051_alu1_n191), .Y(
        oc8051_alu1_n2170) );
  INV_X0P5B_A12TS oc8051_alu1_u178 ( .A(oc8051_alu1_n55), .Y(oc8051_alu1_n173)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_u177 ( .A(oc8051_alu1_n55), .B(oc8051_alu1_n122), .Y(oc8051_alu1_n187) );
  OAI22_X0P5M_A12TS oc8051_alu1_u176 ( .A0(src1[4]), .A1(oc8051_alu1_n173), 
        .B0(oc8051_alu1_n187), .B1(oc8051_alu1_n188), .Y(oc8051_alu1_n186) );
  INV_X0P5B_A12TS oc8051_alu1_u175 ( .A(src2[5]), .Y(oc8051_alu1_n161) );
  INV_X0P5B_A12TS oc8051_alu1_u174 ( .A(src1[5]), .Y(oc8051_alu1_n119) );
  NOR2_X0P5A_A12TS oc8051_alu1_u173 ( .A(oc8051_alu1_n161), .B(
        oc8051_alu1_n119), .Y(oc8051_alu1_n164) );
  AOI21_X0P5M_A12TS oc8051_alu1_u172 ( .A0(oc8051_alu1_n161), .A1(
        oc8051_alu1_n119), .B0(oc8051_alu1_n164), .Y(oc8051_alu1_n182) );
  XOR2_X0P5M_A12TS oc8051_alu1_u171 ( .A(oc8051_alu1_n186), .B(
        oc8051_alu1_n182), .Y(sub_result[5]) );
  INV_X0P5B_A12TS oc8051_alu1_u170 ( .A(oc8051_alu1_n44), .Y(oc8051_alu1_n144)
         );
  AOI22_X0P5M_A12TS oc8051_alu1_u169 ( .A0(oc8051_alu1_n164), .A1(
        oc8051_alu1_n144), .B0(oc8051_alu1_n46), .B1(oc8051_alu1_n182), .Y(
        oc8051_alu1_n184) );
  AOI222_X0P5M_A12TS oc8051_alu1_u168 ( .A0(oc8051_alu1_dec[5]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_inc[5]), .B1(oc8051_alu1_n66), .C0(
        oc8051_alu1_n170), .C1(oc8051_alu1_n119), .Y(oc8051_alu1_n185) );
  OAI211_X0P5M_A12TS oc8051_alu1_u167 ( .A0(oc8051_alu1_n143), .A1(
        oc8051_alu1_n161), .B0(oc8051_alu1_n184), .C0(oc8051_alu1_n185), .Y(
        oc8051_alu1_n120) );
  AOI21_X0P5M_A12TS oc8051_alu1_u166 ( .A0(sub_result[5]), .A1(oc8051_alu1_n24), .B0(oc8051_alu1_n120), .Y(oc8051_alu1_n174) );
  AOI22_X0P5M_A12TS oc8051_alu1_u165 ( .A0(oc8051_alu1_mulsrc1[5]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc1[5]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n175) );
  AOI22_X0P5M_A12TS oc8051_alu1_u164 ( .A0(src1[4]), .A1(oc8051_alu1_n165), 
        .B0(src1[6]), .B1(oc8051_alu1_n124), .Y(oc8051_alu1_n176) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u163 ( .A0(src2[4]), .A1(src1[4]), .B0(
        oc8051_alu1_n54), .C0(oc8051_alu1_n183), .Y(oc8051_alu1_n162) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u162 ( .A(oc8051_alu1_n162), .B(
        oc8051_alu1_n182), .Y(oc8051_alu1_n178) );
  OAI21_X0P5M_A12TS oc8051_alu1_u161 ( .A0(src1[5]), .A1(src1[6]), .B0(src1[7]), .Y(oc8051_alu1_n181) );
  NAND3_X0P5A_A12TS oc8051_alu1_u160 ( .A(oc8051_alu1_n29), .B(
        oc8051_alu1_n133), .C(oc8051_alu1_n181), .Y(oc8051_alu1_n151) );
  NAND2_X0P5A_A12TS oc8051_alu1_u159 ( .A(oc8051_alu1_n180), .B(src1[4]), .Y(
        oc8051_alu1_n159) );
  XNOR3_X0P5M_A12TS oc8051_alu1_u158 ( .A(oc8051_alu1_n151), .B(src1[5]), .C(
        oc8051_alu1_n159), .Y(oc8051_alu1_n179) );
  AOI222_X0P5M_A12TS oc8051_alu1_u157 ( .A0(src1[5]), .A1(oc8051_alu1_n148), 
        .B0(oc8051_alu1_n178), .B1(oc8051_alu1_n289), .C0(oc8051_alu1_n179), 
        .C1(oc8051_alu1_n41), .Y(oc8051_alu1_n177) );
  NAND4_X0P5A_A12TS oc8051_alu1_u156 ( .A(oc8051_alu1_n174), .B(
        oc8051_alu1_n175), .C(oc8051_alu1_n176), .D(oc8051_alu1_n177), .Y(
        oc8051_alu1_n2180) );
  XOR2_X0P5M_A12TS oc8051_alu1_u155 ( .A(src2[6]), .B(src1[6]), .Y(
        oc8051_alu1_n160) );
  NOR2_X0P5A_A12TS oc8051_alu1_u154 ( .A(src1[4]), .B(oc8051_alu1_n173), .Y(
        oc8051_alu1_n172) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u153 ( .A0(oc8051_alu1_n55), .A1(
        oc8051_alu1_n122), .B0(src2[4]), .C0(oc8051_alu1_n172), .Y(
        oc8051_alu1_n171) );
  CGENI_X1M_A12TS oc8051_alu1_u152 ( .A(src1[5]), .B(oc8051_alu1_n161), .CI(
        oc8051_alu1_n171), .CON(oc8051_alu1_n136) );
  XOR2_X0P5M_A12TS oc8051_alu1_u151 ( .A(oc8051_alu1_n160), .B(
        oc8051_alu1_n136), .Y(sub_result[6]) );
  INV_X0P5B_A12TS oc8051_alu1_u150 ( .A(src1[6]), .Y(oc8051_alu1_n116) );
  AOI22_X0P5M_A12TS oc8051_alu1_u149 ( .A0(oc8051_alu1_n170), .A1(
        oc8051_alu1_n116), .B0(oc8051_alu1_dec[6]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n166) );
  INV_X0P5B_A12TS oc8051_alu1_u148 ( .A(src2[6]), .Y(oc8051_alu1_n169) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u147 ( .A0(oc8051_alu1_n116), .A1(
        oc8051_alu1_n44), .B0(oc8051_alu1_n143), .C0(oc8051_alu1_n169), .Y(
        oc8051_alu1_n168) );
  AOI221_X0P5M_A12TS oc8051_alu1_u146 ( .A0(oc8051_alu1_inc[6]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_n46), .B1(oc8051_alu1_n160), .C0(
        oc8051_alu1_n168), .Y(oc8051_alu1_n167) );
  NAND2_X0P5A_A12TS oc8051_alu1_u145 ( .A(oc8051_alu1_n166), .B(
        oc8051_alu1_n167), .Y(oc8051_alu1_n117) );
  AOI21_X0P5M_A12TS oc8051_alu1_u144 ( .A0(oc8051_alu1_n24), .A1(sub_result[6]), .B0(oc8051_alu1_n117), .Y(oc8051_alu1_n153) );
  AOI22_X0P5M_A12TS oc8051_alu1_u143 ( .A0(oc8051_alu1_mulsrc1[6]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc1[6]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n154) );
  AOI22_X0P5M_A12TS oc8051_alu1_u142 ( .A0(src1[5]), .A1(oc8051_alu1_n165), 
        .B0(src1[7]), .B1(oc8051_alu1_n124), .Y(oc8051_alu1_n155) );
  INV_X0P5B_A12TS oc8051_alu1_u141 ( .A(oc8051_alu1_n164), .Y(oc8051_alu1_n163) );
  AO21A1AI2_X0P5M_A12TS oc8051_alu1_u140 ( .A0(oc8051_alu1_n161), .A1(
        oc8051_alu1_n119), .B0(oc8051_alu1_n162), .C0(oc8051_alu1_n163), .Y(
        oc8051_alu1_n149) );
  XOR2_X0P5M_A12TS oc8051_alu1_u139 ( .A(oc8051_alu1_n149), .B(
        oc8051_alu1_n160), .Y(oc8051_alu1_n157) );
  AO1B2_X0P5M_A12TS oc8051_alu1_u138 ( .B0(oc8051_alu1_n151), .B1(src1[5]), 
        .A0N(oc8051_alu1_n159), .Y(oc8051_alu1_n152) );
  XNOR3_X0P5M_A12TS oc8051_alu1_u137 ( .A(oc8051_alu1_n116), .B(
        oc8051_alu1_n151), .C(oc8051_alu1_n152), .Y(oc8051_alu1_n158) );
  AOI222_X0P5M_A12TS oc8051_alu1_u136 ( .A0(src1[6]), .A1(oc8051_alu1_n148), 
        .B0(oc8051_alu1_n157), .B1(oc8051_alu1_n289), .C0(oc8051_alu1_n41), 
        .C1(oc8051_alu1_n158), .Y(oc8051_alu1_n156) );
  NAND4_X0P5A_A12TS oc8051_alu1_u135 ( .A(oc8051_alu1_n153), .B(
        oc8051_alu1_n154), .C(oc8051_alu1_n155), .D(oc8051_alu1_n156), .Y(
        oc8051_alu1_n2190) );
  AOI21_X0P5M_A12TS oc8051_alu1_u134 ( .A0(oc8051_alu1_n151), .A1(src1[6]), 
        .B0(oc8051_alu1_n152), .Y(oc8051_alu1_n39) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u133 ( .AN(oc8051_alu1_n149), .B(
        oc8051_alu1_n116), .Y(oc8051_alu1_n150) );
  OAI22_X0P5M_A12TS oc8051_alu1_u132 ( .A0(src1[6]), .A1(oc8051_alu1_n149), 
        .B0(src2[6]), .B1(oc8051_alu1_n150), .Y(oc8051_alu1_n18) );
  XOR2_X0P5M_A12TS oc8051_alu1_u131 ( .A(src2[7]), .B(oc8051_alu1_n18), .Y(
        oc8051_alu1_n112) );
  OAI22_X0P5M_A12TS oc8051_alu1_u130 ( .A0(oc8051_alu1_n39), .A1(
        oc8051_alu1_n47), .B0(oc8051_alu1_n112), .B1(oc8051_alu1_n111), .Y(
        oc8051_alu1_n145) );
  AOI221_X0P5M_A12TS oc8051_alu1_u129 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n112), .B0(oc8051_alu1_n41), .B1(oc8051_alu1_n39), .C0(
        oc8051_alu1_n148), .Y(oc8051_alu1_n147) );
  INV_X0P5B_A12TS oc8051_alu1_u128 ( .A(oc8051_alu1_n147), .Y(oc8051_alu1_n146) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u127 ( .A(oc8051_alu1_n145), .B(
        oc8051_alu1_n146), .S0(src1[7]), .Y(oc8051_alu1_n129) );
  INV_X0P5B_A12TS oc8051_alu1_u126 ( .A(src1[7]), .Y(oc8051_alu1_n40) );
  NOR2_X0P5A_A12TS oc8051_alu1_u125 ( .A(oc8051_alu1_n40), .B(oc8051_alu1_n48), 
        .Y(oc8051_alu1_n140) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u124 ( .A(oc8051_alu1_n46), .B(
        oc8051_alu1_n144), .S0(src1[7]), .Y(oc8051_alu1_n142) );
  NAND2_X0P5A_A12TS oc8051_alu1_u123 ( .A(oc8051_alu1_n142), .B(
        oc8051_alu1_n143), .Y(oc8051_alu1_n141) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u122 ( .A(oc8051_alu1_n140), .B(
        oc8051_alu1_n141), .S0(src2[7]), .Y(oc8051_alu1_n138) );
  AOI22_X0P5M_A12TS oc8051_alu1_u121 ( .A0(oc8051_alu1_inc[7]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[7]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n139) );
  OA211_X0P5M_A12TS oc8051_alu1_u120 ( .A0(src1[7]), .A1(oc8051_alu1_n50), 
        .B0(oc8051_alu1_n138), .C0(oc8051_alu1_n139), .Y(oc8051_alu1_n113) );
  NAND2B_X0P5M_A12TS oc8051_alu1_u119 ( .AN(oc8051_alu1_n136), .B(src1[6]), 
        .Y(oc8051_alu1_n137) );
  AOI22_X0P5M_A12TS oc8051_alu1_u118 ( .A0(oc8051_alu1_n116), .A1(
        oc8051_alu1_n136), .B0(oc8051_alu1_n137), .B1(src2[6]), .Y(
        oc8051_alu1_n20) );
  INV_X0P5B_A12TS oc8051_alu1_u117 ( .A(src2[7]), .Y(oc8051_alu1_n31) );
  XOR2_X0P5M_A12TS oc8051_alu1_u116 ( .A(oc8051_alu1_n20), .B(oc8051_alu1_n31), 
        .Y(oc8051_alu1_n135) );
  NAND2_X0P5A_A12TS oc8051_alu1_u115 ( .A(oc8051_alu1_n135), .B(
        oc8051_alu1_n40), .Y(oc8051_alu1_n32) );
  OAI21_X0P5M_A12TS oc8051_alu1_u114 ( .A0(oc8051_alu1_n135), .A1(
        oc8051_alu1_n40), .B0(oc8051_alu1_n32), .Y(sub_result[7]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u113 ( .A0(oc8051_alu1_divsrc1[7]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n24), .B1(sub_result[7]), .Y(
        oc8051_alu1_n130) );
  INV_X0P5B_A12TS oc8051_alu1_u112 ( .A(oc8051_alu1_n134), .Y(oc8051_alu1_n45)
         );
  OAI22_X0P5M_A12TS oc8051_alu1_u111 ( .A0(oc8051_alu1_n133), .A1(
        oc8051_alu1_n28), .B0(oc8051_alu1_n126), .B1(oc8051_alu1_n116), .Y(
        oc8051_alu1_n132) );
  AOI221_X0P5M_A12TS oc8051_alu1_u110 ( .A0(oc8051_alu1_n45), .A1(src1[0]), 
        .B0(oc8051_alu1_mulsrc1[7]), .B1(oc8051_alu1_n290), .C0(
        oc8051_alu1_n132), .Y(oc8051_alu1_n131) );
  NAND4_X0P5A_A12TS oc8051_alu1_u109 ( .A(oc8051_alu1_n129), .B(
        oc8051_alu1_n113), .C(oc8051_alu1_n130), .D(oc8051_alu1_n131), .Y(
        oc8051_alu1_n2200) );
  NAND2_X0P5A_A12TS oc8051_alu1_u108 ( .A(oc8051_alu1_malicious1), .B(
        oc8051_alu1_n46), .Y(oc8051_alu1_n2400) );
  INV_X0P5B_A12TS oc8051_alu1_u107 ( .A(oc8051_alu1_n2400), .Y(oc8051_alu1_n1)
         );
  AND4_X0P5M_A12TS oc8051_alu1_u106 ( .A(oc8051_alu1_n47), .B(oc8051_alu1_n127), .C(oc8051_alu1_n128), .D(oc8051_alu1_n111), .Y(oc8051_alu1_n125) );
  NAND4B_X0P5M_A12TS oc8051_alu1_u105 ( .AN(oc8051_alu1_n124), .B(
        oc8051_alu1_n125), .C(oc8051_alu1_n35), .D(oc8051_alu1_n126), .Y(
        oc8051_alu1_n6) );
  INV_X0P5B_A12TS oc8051_alu1_u104 ( .A(oc8051_alu1_n6), .Y(oc8051_alu1_n3) );
  AND3_X0P5M_A12TS oc8051_alu1_u103 ( .A(oc8051_alu1_n36), .B(oc8051_alu1_n3), 
        .C(oc8051_alu1_n123), .Y(oc8051_alu1_n114) );
  INV_X0P5B_A12TS oc8051_alu1_u102 ( .A(oc8051_alu1_n120), .Y(oc8051_alu1_n118) );
  INV_X0P5B_A12TS oc8051_alu1_u101 ( .A(oc8051_alu1_n117), .Y(oc8051_alu1_n115) );
  OAI22_X0P5M_A12TS oc8051_alu1_u100 ( .A0(oc8051_alu1_n31), .A1(
        oc8051_alu1_n18), .B0(oc8051_alu1_n112), .B1(oc8051_alu1_n40), .Y(
        oc8051_alu1_n104) );
  INV_X0P5B_A12TS oc8051_alu1_u99 ( .A(oc8051_alu1_n104), .Y(oc8051_alu1_n110)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_u98 ( .A(oc8051_alu1_n111), .B(oc8051_alu1_n110), .Y(oc8051_alu1_n26) );
  INV_X0P5B_A12TS oc8051_alu1_u97 ( .A(oc8051_alu1_n26), .Y(oc8051_alu1_n17)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_u96 ( .A(oc8051_alu1_n289), .B(
        oc8051_alu1_n110), .Y(oc8051_alu1_n16) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u95 ( .A(oc8051_alu1_n17), .B(oc8051_alu1_n16), 
        .S0(src3[0]), .Y(oc8051_alu1_n109) );
  AOI21_X0P5M_A12TS oc8051_alu1_u94 ( .A0(oc8051_alu1_dec[8]), .A1(
        oc8051_alu1_n67), .B0(oc8051_alu1_n109), .Y(oc8051_alu1_n105) );
  AOI22_X0P5M_A12TS oc8051_alu1_u93 ( .A0(oc8051_alu1_n92), .A1(src1[0]), .B0(
        oc8051_alu1_inc[8]), .B1(oc8051_alu1_n66), .Y(oc8051_alu1_n106) );
  AOI22_X0P5M_A12TS oc8051_alu1_u92 ( .A0(oc8051_alu1_mulsrc2[0]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc2[0]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n107) );
  INV_X0P5B_A12TS oc8051_alu1_u91 ( .A(oc8051_alu1_n35), .Y(oc8051_alu1_n56)
         );
  AOI22_X0P5M_A12TS oc8051_alu1_u90 ( .A0(oc8051_alu1_n56), .A1(src2[0]), .B0(
        oc8051_alu1_n51), .B1(src1[4]), .Y(oc8051_alu1_n108) );
  NAND4_X0P5A_A12TS oc8051_alu1_u89 ( .A(oc8051_alu1_n105), .B(
        oc8051_alu1_n106), .C(oc8051_alu1_n107), .D(oc8051_alu1_n108), .Y(
        des2[0]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u88 ( .A0(oc8051_alu1_inc[9]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[9]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n99) );
  AOI22_X0P5M_A12TS oc8051_alu1_u87 ( .A0(oc8051_alu1_divsrc2[1]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n92), .B1(src1[1]), .Y(
        oc8051_alu1_n100) );
  AOI22_X0P5M_A12TS oc8051_alu1_u86 ( .A0(oc8051_alu1_n51), .A1(src1[5]), .B0(
        oc8051_alu1_mulsrc2[1]), .B1(oc8051_alu1_n290), .Y(oc8051_alu1_n101)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_u85 ( .A(oc8051_alu1_n104), .B(src3[0]), .Y(
        oc8051_alu1_n98) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u84 ( .A(src3[1]), .B(oc8051_alu1_n98), .Y(
        oc8051_alu1_n103) );
  AOI22_X0P5M_A12TS oc8051_alu1_u83 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n103), .B0(oc8051_alu1_n56), .B1(src2[1]), .Y(
        oc8051_alu1_n102) );
  NAND4_X0P5A_A12TS oc8051_alu1_u82 ( .A(oc8051_alu1_n99), .B(oc8051_alu1_n100), .C(oc8051_alu1_n101), .D(oc8051_alu1_n102), .Y(des2[1]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u81 ( .A0(oc8051_alu1_inc[10]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[10]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n93) );
  AOI22_X0P5M_A12TS oc8051_alu1_u80 ( .A0(oc8051_alu1_divsrc2[2]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n92), .B1(src1[2]), .Y(
        oc8051_alu1_n94) );
  AOI22_X0P5M_A12TS oc8051_alu1_u79 ( .A0(oc8051_alu1_n51), .A1(src1[6]), .B0(
        oc8051_alu1_mulsrc2[2]), .B1(oc8051_alu1_n290), .Y(oc8051_alu1_n95) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u78 ( .AN(src3[1]), .B(oc8051_alu1_n98), .Y(
        oc8051_alu1_n91) );
  XOR2_X0P5M_A12TS oc8051_alu1_u77 ( .A(src3[2]), .B(oc8051_alu1_n91), .Y(
        oc8051_alu1_n97) );
  AOI22_X0P5M_A12TS oc8051_alu1_u76 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n97), .B0(oc8051_alu1_n56), .B1(src2[2]), .Y(
        oc8051_alu1_n96) );
  NAND4_X0P5A_A12TS oc8051_alu1_u75 ( .A(oc8051_alu1_n93), .B(oc8051_alu1_n94), 
        .C(oc8051_alu1_n95), .D(oc8051_alu1_n96), .Y(des2[2]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u74 ( .A0(oc8051_alu1_inc[11]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[11]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n86) );
  AOI22_X0P5M_A12TS oc8051_alu1_u73 ( .A0(oc8051_alu1_divsrc2[3]), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n92), .B1(src1[3]), .Y(
        oc8051_alu1_n87) );
  AOI22_X0P5M_A12TS oc8051_alu1_u72 ( .A0(oc8051_alu1_n51), .A1(src1[7]), .B0(
        oc8051_alu1_mulsrc2[3]), .B1(oc8051_alu1_n290), .Y(oc8051_alu1_n88) );
  NAND2_X0P5A_A12TS oc8051_alu1_u71 ( .A(src3[2]), .B(oc8051_alu1_n91), .Y(
        oc8051_alu1_n85) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u70 ( .A(src3[3]), .B(oc8051_alu1_n85), .Y(
        oc8051_alu1_n90) );
  AOI22_X0P5M_A12TS oc8051_alu1_u69 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n90), .B0(oc8051_alu1_n56), .B1(src2[3]), .Y(
        oc8051_alu1_n89) );
  NAND4_X0P5A_A12TS oc8051_alu1_u68 ( .A(oc8051_alu1_n86), .B(oc8051_alu1_n87), 
        .C(oc8051_alu1_n88), .D(oc8051_alu1_n89), .Y(des2[3]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u67 ( .A0(oc8051_alu1_inc[12]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[12]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n80) );
  AOI22_X0P5M_A12TS oc8051_alu1_u66 ( .A0(oc8051_alu1_mulsrc2[4]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc2[4]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n81) );
  AOI22_X0P5M_A12TS oc8051_alu1_u65 ( .A0(oc8051_alu1_n65), .A1(src1[4]), .B0(
        oc8051_alu1_n51), .B1(src1[0]), .Y(oc8051_alu1_n82) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u64 ( .AN(src3[3]), .B(oc8051_alu1_n85), .Y(
        oc8051_alu1_n79) );
  XOR2_X0P5M_A12TS oc8051_alu1_u63 ( .A(src3[4]), .B(oc8051_alu1_n79), .Y(
        oc8051_alu1_n84) );
  AOI22_X0P5M_A12TS oc8051_alu1_u62 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n84), .B0(src2[4]), .B1(oc8051_alu1_n62), .Y(
        oc8051_alu1_n83) );
  NAND4_X0P5A_A12TS oc8051_alu1_u61 ( .A(oc8051_alu1_n80), .B(oc8051_alu1_n81), 
        .C(oc8051_alu1_n82), .D(oc8051_alu1_n83), .Y(des2[4]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u60 ( .A0(oc8051_alu1_inc[13]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[13]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n74) );
  AOI22_X0P5M_A12TS oc8051_alu1_u59 ( .A0(oc8051_alu1_mulsrc2[5]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc2[5]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n75) );
  AOI22_X0P5M_A12TS oc8051_alu1_u58 ( .A0(oc8051_alu1_n65), .A1(src1[5]), .B0(
        oc8051_alu1_n51), .B1(src1[1]), .Y(oc8051_alu1_n76) );
  NAND2_X0P5A_A12TS oc8051_alu1_u57 ( .A(src3[4]), .B(oc8051_alu1_n79), .Y(
        oc8051_alu1_n73) );
  XNOR2_X0P5M_A12TS oc8051_alu1_u56 ( .A(src3[5]), .B(oc8051_alu1_n73), .Y(
        oc8051_alu1_n78) );
  AOI22_X0P5M_A12TS oc8051_alu1_u55 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n78), .B0(src2[5]), .B1(oc8051_alu1_n62), .Y(
        oc8051_alu1_n77) );
  NAND4_X0P5A_A12TS oc8051_alu1_u54 ( .A(oc8051_alu1_n74), .B(oc8051_alu1_n75), 
        .C(oc8051_alu1_n76), .D(oc8051_alu1_n77), .Y(des2[5]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u53 ( .A0(oc8051_alu1_inc[14]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[14]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n68) );
  AOI22_X0P5M_A12TS oc8051_alu1_u52 ( .A0(oc8051_alu1_mulsrc2[6]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc2[6]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n69) );
  AOI22_X0P5M_A12TS oc8051_alu1_u51 ( .A0(oc8051_alu1_n65), .A1(src1[6]), .B0(
        oc8051_alu1_n51), .B1(src1[2]), .Y(oc8051_alu1_n70) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u50 ( .AN(src3[5]), .B(oc8051_alu1_n73), .Y(
        oc8051_alu1_n64) );
  XOR2_X0P5M_A12TS oc8051_alu1_u49 ( .A(src3[6]), .B(oc8051_alu1_n64), .Y(
        oc8051_alu1_n72) );
  AOI22_X0P5M_A12TS oc8051_alu1_u48 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n72), .B0(src2[6]), .B1(oc8051_alu1_n62), .Y(
        oc8051_alu1_n71) );
  NAND4_X0P5A_A12TS oc8051_alu1_u47 ( .A(oc8051_alu1_n68), .B(oc8051_alu1_n69), 
        .C(oc8051_alu1_n70), .D(oc8051_alu1_n71), .Y(des2[6]) );
  AOI22_X0P5M_A12TS oc8051_alu1_u46 ( .A0(oc8051_alu1_inc[15]), .A1(
        oc8051_alu1_n66), .B0(oc8051_alu1_dec[15]), .B1(oc8051_alu1_n67), .Y(
        oc8051_alu1_n57) );
  AOI22_X0P5M_A12TS oc8051_alu1_u45 ( .A0(oc8051_alu1_mulsrc2[7]), .A1(
        oc8051_alu1_n290), .B0(oc8051_alu1_divsrc2[7]), .B1(oc8051_alu1_n288), 
        .Y(oc8051_alu1_n58) );
  AOI22_X0P5M_A12TS oc8051_alu1_u44 ( .A0(oc8051_alu1_n65), .A1(src1[7]), .B0(
        oc8051_alu1_n51), .B1(src1[3]), .Y(oc8051_alu1_n59) );
  AND2_X0P5M_A12TS oc8051_alu1_u43 ( .A(oc8051_alu1_n64), .B(src3[6]), .Y(
        oc8051_alu1_n63) );
  XOR2_X0P5M_A12TS oc8051_alu1_u42 ( .A(src3[7]), .B(oc8051_alu1_n63), .Y(
        oc8051_alu1_n61) );
  AOI22_X0P5M_A12TS oc8051_alu1_u41 ( .A0(oc8051_alu1_n289), .A1(
        oc8051_alu1_n61), .B0(src2[7]), .B1(oc8051_alu1_n62), .Y(
        oc8051_alu1_n60) );
  NAND4_X0P5A_A12TS oc8051_alu1_u40 ( .A(oc8051_alu1_n57), .B(oc8051_alu1_n58), 
        .C(oc8051_alu1_n59), .D(oc8051_alu1_n60), .Y(des2[7]) );
  AOI222_X0P5M_A12TS oc8051_alu1_u39 ( .A0(oc8051_alu1_n54), .A1(
        oc8051_alu1_n289), .B0(oc8051_alu1_n55), .B1(oc8051_alu1_n24), .C0(
        oc8051_alu1_n56), .C1(srcac), .Y(oc8051_alu1_n53) );
  INV_X0P5B_A12TS oc8051_alu1_u38 ( .A(oc8051_alu1_n53), .Y(desac) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u37 ( .A(oc8051_alu1_n37), .B(oc8051_alu1_n36), 
        .S0(bit_out), .Y(oc8051_alu1_n52) );
  AOI21_X0P5M_A12TS oc8051_alu1_u36 ( .A0(oc8051_alu1_n51), .A1(src1[7]), .B0(
        oc8051_alu1_n52), .Y(oc8051_alu1_n21) );
  INV_X0P5B_A12TS oc8051_alu1_u35 ( .A(bit_out), .Y(oc8051_alu1_n49) );
  OAI221_X0P5M_A12TS oc8051_alu1_u34 ( .A0(oc8051_alu1_n39), .A1(
        oc8051_alu1_n47), .B0(oc8051_alu1_n48), .B1(oc8051_alu1_n49), .C0(
        oc8051_alu1_n50), .Y(oc8051_alu1_n33) );
  NOR2_X0P5A_A12TS oc8051_alu1_u33 ( .A(oc8051_alu1_n45), .B(oc8051_alu1_n46), 
        .Y(oc8051_alu1_n43) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u32 ( .A(oc8051_alu1_n43), .B(oc8051_alu1_n44), 
        .S0(bit_out), .Y(oc8051_alu1_n42) );
  OA21A1OI2_X0P5M_A12TS oc8051_alu1_u31 ( .A0(oc8051_alu1_n39), .A1(
        oc8051_alu1_n40), .B0(oc8051_alu1_n41), .C0(oc8051_alu1_n42), .Y(
        oc8051_alu1_n38) );
  NAND4_X0P5A_A12TS oc8051_alu1_u30 ( .A(oc8051_alu1_n35), .B(oc8051_alu1_n36), 
        .C(oc8051_alu1_n37), .D(oc8051_alu1_n38), .Y(oc8051_alu1_n34) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u29 ( .A(oc8051_alu1_n33), .B(oc8051_alu1_n34), 
        .S0(alu_cy), .Y(oc8051_alu1_n22) );
  OAI21_X0P5M_A12TS oc8051_alu1_u28 ( .A0(oc8051_alu1_n20), .A1(
        oc8051_alu1_n31), .B0(oc8051_alu1_n32), .Y(oc8051_alu1_n19) );
  OAI22_X0P5M_A12TS oc8051_alu1_u27 ( .A0(oc8051_alu1_n27), .A1(
        oc8051_alu1_n28), .B0(oc8051_alu1_n29), .B1(oc8051_alu1_n30), .Y(
        oc8051_alu1_n25) );
  AOI211_X0P5M_A12TS oc8051_alu1_u26 ( .A0(oc8051_alu1_n24), .A1(
        oc8051_alu1_n19), .B0(oc8051_alu1_n25), .C0(oc8051_alu1_n26), .Y(
        oc8051_alu1_n23) );
  AOI31_X0P5M_A12TS oc8051_alu1_u25 ( .A0(oc8051_alu1_n21), .A1(
        oc8051_alu1_n22), .A2(oc8051_alu1_n23), .B0(oc8051_alu1_n1), .Y(descy)
         );
  XOR2_X0P5M_A12TS oc8051_alu1_u24 ( .A(oc8051_alu1_n19), .B(oc8051_alu1_n20), 
        .Y(oc8051_alu1_n10) );
  NAND2_X0P5A_A12TS oc8051_alu1_u23 ( .A(oc8051_alu1_mulov), .B(
        oc8051_alu1_n290), .Y(oc8051_alu1_n12) );
  MXIT2_X0P5M_A12TS oc8051_alu1_u22 ( .A(oc8051_alu1_n16), .B(oc8051_alu1_n17), 
        .S0(oc8051_alu1_n18), .Y(oc8051_alu1_n15) );
  AOI21_X0P5M_A12TS oc8051_alu1_u21 ( .A0(oc8051_alu1_divov), .A1(
        oc8051_alu1_n288), .B0(oc8051_alu1_n15), .Y(oc8051_alu1_n13) );
  OAI211_X0P5M_A12TS oc8051_alu1_u20 ( .A0(oc8051_alu1_n10), .A1(
        oc8051_alu1_n11), .B0(oc8051_alu1_n12), .C0(oc8051_alu1_n13), .Y(desov) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u19 ( .AN(oc8051_alu1_des_acc_1[0]), .B(
        oc8051_alu1_n1), .Y(des_acc[0]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u18 ( .AN(oc8051_alu1_des_acc_1[1]), .B(
        oc8051_alu1_n1), .Y(des_acc[1]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u17 ( .AN(oc8051_alu1_des_acc_1[2]), .B(
        oc8051_alu1_n1), .Y(des_acc[2]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u16 ( .AN(oc8051_alu1_des_acc_1[3]), .B(
        oc8051_alu1_n1), .Y(des_acc[3]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u15 ( .AN(oc8051_alu1_des_acc_1[4]), .B(
        oc8051_alu1_n1), .Y(des_acc[4]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u14 ( .AN(oc8051_alu1_des_acc_1[5]), .B(
        oc8051_alu1_n1), .Y(des_acc[5]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u13 ( .AN(oc8051_alu1_des_acc_1[6]), .B(
        oc8051_alu1_n1), .Y(des_acc[6]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_u12 ( .AN(oc8051_alu1_des_acc_1[7]), .B(
        oc8051_alu1_n1), .Y(des_acc[7]) );
  AO22_X0P5M_A12TS oc8051_alu1_u11 ( .A0(oc8051_alu1_n2400), .A1(
        oc8051_alu1_n9), .B0(oc8051_alu1_n6), .B1(src1[0]), .Y(wr_dat[0]) );
  AO22_X0P5M_A12TS oc8051_alu1_u10 ( .A0(oc8051_alu1_n2400), .A1(
        oc8051_alu1_n5), .B0(oc8051_alu1_n6), .B1(src1[2]), .Y(wr_dat[2]) );
  TIEHI_X1M_A12TS oc8051_alu1_u9 ( .Y(oc8051_alu1_n14) );
  OAI22_X1M_A12TS oc8051_alu1_u8 ( .A0(oc8051_alu1_n1), .A1(oc8051_alu1_n115), 
        .B0(oc8051_alu1_n114), .B1(oc8051_alu1_n116), .Y(wr_dat[6]) );
  OAI22_X1M_A12TS oc8051_alu1_u7 ( .A0(oc8051_alu1_n1), .A1(oc8051_alu1_n113), 
        .B0(oc8051_alu1_n114), .B1(oc8051_alu1_n40), .Y(wr_dat[7]) );
  OAI22_X1M_A12TS oc8051_alu1_u6 ( .A0(oc8051_alu1_n1), .A1(oc8051_alu1_n118), 
        .B0(oc8051_alu1_n114), .B1(oc8051_alu1_n119), .Y(wr_dat[5]) );
  OAI22_X1M_A12TS oc8051_alu1_u5 ( .A0(oc8051_alu1_n1), .A1(oc8051_alu1_n121), 
        .B0(oc8051_alu1_n114), .B1(oc8051_alu1_n122), .Y(wr_dat[4]) );
  OAI22_X1M_A12TS oc8051_alu1_u4 ( .A0(oc8051_alu1_n1), .A1(oc8051_alu1_n2), 
        .B0(oc8051_alu1_n3), .B1(oc8051_alu1_n4), .Y(wr_dat[3]) );
  OAI22_X1M_A12TS oc8051_alu1_u3 ( .A0(oc8051_alu1_n1), .A1(oc8051_alu1_n7), 
        .B0(oc8051_alu1_n3), .B1(oc8051_alu1_n8), .Y(wr_dat[1]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_0_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2130), .Q(oc8051_alu1_des_acc_1[0]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_1_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2140), .Q(oc8051_alu1_des_acc_1[1]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_2_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2150), .Q(oc8051_alu1_des_acc_1[2]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_3_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2160), .Q(oc8051_alu1_des_acc_1[3]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_4_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2170), .Q(oc8051_alu1_des_acc_1[4]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_5_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2180), .Q(oc8051_alu1_des_acc_1[5]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_6_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2190), .Q(oc8051_alu1_des_acc_1[6]) );
  LATQ_X1M_A12TS oc8051_alu1_des_acc_1_reg_7_ ( .G(oc8051_alu1_n2400), .D(
        oc8051_alu1_n2200), .Q(oc8051_alu1_des_acc_1[7]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_alu_malicious_u12 ( .AN(oc8051_alu1_n289), .B(
        wb_rst_i), .Y(oc8051_alu1_alu_malicious_n5) );
  INV_X0P5B_A12TS oc8051_alu1_alu_malicious_u11 ( .A(
        oc8051_alu1_alu_malicious_state_0_), .Y(oc8051_alu1_alu_malicious_n2)
         );
  NAND2_X0P5A_A12TS oc8051_alu1_alu_malicious_u10 ( .A(
        oc8051_alu1_alu_malicious_n5), .B(oc8051_alu1_alu_malicious_n2), .Y(
        oc8051_alu1_alu_malicious_n7) );
  INV_X0P5B_A12TS oc8051_alu1_alu_malicious_u9 ( .A(
        oc8051_alu1_alu_malicious_n7), .Y(oc8051_alu1_alu_malicious_n70) );
  NAND2_X0P5A_A12TS oc8051_alu1_alu_malicious_u8 ( .A(
        oc8051_alu1_alu_malicious_n5), .B(oc8051_alu1_alu_malicious_state_0_), 
        .Y(oc8051_alu1_alu_malicious_n6) );
  MXIT2_X0P5M_A12TS oc8051_alu1_alu_malicious_u7 ( .A(
        oc8051_alu1_alu_malicious_n6), .B(oc8051_alu1_alu_malicious_n7), .S0(
        oc8051_alu1_alu_malicious_state_1_), .Y(oc8051_alu1_alu_malicious_n8)
         );
  AOI2XB1_X0P5M_A12TS oc8051_alu1_alu_malicious_u6 ( .A1N(
        oc8051_alu1_alu_malicious_state_1_), .A0(oc8051_alu1_alu_malicious_n5), 
        .B0(oc8051_alu1_alu_malicious_n70), .Y(oc8051_alu1_alu_malicious_n3)
         );
  NAND3_X0P5A_A12TS oc8051_alu1_alu_malicious_u5 ( .A(
        oc8051_alu1_alu_malicious_n5), .B(oc8051_alu1_alu_malicious_state_0_), 
        .C(oc8051_alu1_alu_malicious_state_1_), .Y(
        oc8051_alu1_alu_malicious_n4) );
  MXIT2_X0P5M_A12TS oc8051_alu1_alu_malicious_u4 ( .A(
        oc8051_alu1_alu_malicious_n3), .B(oc8051_alu1_alu_malicious_n4), .S0(
        oc8051_alu1_alu_malicious_n1), .Y(oc8051_alu1_alu_malicious_n9) );
  NOR3_X0P5A_A12TS oc8051_alu1_alu_malicious_u3 ( .A(
        oc8051_alu1_alu_malicious_n2), .B(oc8051_alu1_alu_malicious_state_1_), 
        .C(oc8051_alu1_alu_malicious_n1), .Y(oc8051_alu1_malicious1) );
  DFFQN_X1M_A12TS oc8051_alu1_alu_malicious_state_reg_2_ ( .D(
        oc8051_alu1_alu_malicious_n9), .CK(wb_clk_i), .QN(
        oc8051_alu1_alu_malicious_n1) );
  DFFQ_X1M_A12TS oc8051_alu1_alu_malicious_state_reg_1_ ( .D(
        oc8051_alu1_alu_malicious_n8), .CK(wb_clk_i), .Q(
        oc8051_alu1_alu_malicious_state_1_) );
  DFFQ_X1M_A12TS oc8051_alu1_alu_malicious_state_reg_0_ ( .D(
        oc8051_alu1_alu_malicious_n70), .CK(wb_clk_i), .Q(
        oc8051_alu1_alu_malicious_state_0_) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u74 ( .AN(
        oc8051_alu1_oc8051_mul1_cycle_1_), .B(oc8051_alu1_oc8051_mul1_cycle_0_), .Y(oc8051_alu1_oc8051_mul1_n1) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u73 ( .A(
        oc8051_alu1_oc8051_mul1_cycle_0_), .B(oc8051_alu1_oc8051_mul1_cycle_1_), .Y(oc8051_alu1_oc8051_mul1_n20) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u72 ( .A0(src2[2]), .A1(
        oc8051_alu1_oc8051_mul1_n1), .B0(src2[6]), .B1(
        oc8051_alu1_oc8051_mul1_n20), .Y(oc8051_alu1_oc8051_mul1_n53) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u71 ( .AN(
        oc8051_alu1_oc8051_mul1_cycle_0_), .B(oc8051_alu1_oc8051_mul1_cycle_1_), .Y(oc8051_alu1_oc8051_mul1_n3) );
  AOI32_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u70 ( .A0(
        oc8051_alu1_oc8051_mul1_cycle_0_), .A1(
        oc8051_alu1_oc8051_mul1_cycle_1_), .A2(src2[0]), .B0(src2[4]), .B1(
        oc8051_alu1_oc8051_mul1_n3), .Y(oc8051_alu1_oc8051_mul1_n54) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u69 ( .A(
        oc8051_alu1_oc8051_mul1_n53), .B(oc8051_alu1_oc8051_mul1_n54), .Y(
        oc8051_alu1_oc8051_mul1_n70) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u68 ( .A0(src2[3]), .A1(
        oc8051_alu1_oc8051_mul1_n1), .B0(src2[7]), .B1(
        oc8051_alu1_oc8051_mul1_n20), .Y(oc8051_alu1_oc8051_mul1_n51) );
  AOI32_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u67 ( .A0(
        oc8051_alu1_oc8051_mul1_cycle_0_), .A1(
        oc8051_alu1_oc8051_mul1_cycle_1_), .A2(src2[1]), .B0(src2[5]), .B1(
        oc8051_alu1_oc8051_mul1_n3), .Y(oc8051_alu1_oc8051_mul1_n52) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u66 ( .A(
        oc8051_alu1_oc8051_mul1_n51), .B(oc8051_alu1_oc8051_mul1_n52), .Y(
        oc8051_alu1_oc8051_mul1_n80) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u65 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul_1_), .B(oc8051_alu1_oc8051_mul1_n20), 
        .Y(oc8051_alu1_oc8051_mul1_n16) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u64 ( .A(oc8051_alu1_oc8051_mul1_n20), .Y(oc8051_alu1_oc8051_mul1_n25) );
  AND3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u63 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1_2_), .B(
        oc8051_alu1_oc8051_mul1_n25), .C(oc8051_alu1_oc8051_mul1_tmp_mul_0_), 
        .Y(oc8051_alu1_oc8051_mul1_n18) );
  CGENI_X1M_A12TS oc8051_alu1_oc8051_mul1_u62 ( .A(oc8051_alu1_oc8051_mul1_n16), .B(oc8051_alu1_oc8051_mul1_mul_result1_3_), .CI(oc8051_alu1_oc8051_mul1_n18), 
        .CON(oc8051_alu1_oc8051_mul1_n15) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u61 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_2_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n14) );
  AND2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u60 ( .A(
        oc8051_alu1_oc8051_mul1_n14), .B(oc8051_alu1_oc8051_mul1_n15), .Y(
        oc8051_alu1_oc8051_mul1_n50) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u59 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1_4_), .Y(
        oc8051_alu1_oc8051_mul1_n13) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u58 ( .A0(
        oc8051_alu1_oc8051_mul1_n15), .A1(oc8051_alu1_oc8051_mul1_n14), .B0(
        oc8051_alu1_oc8051_mul1_n50), .B1(oc8051_alu1_oc8051_mul1_n13), .Y(
        oc8051_alu1_oc8051_mul1_n11) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u57 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_3_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n12) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u56 ( .A(oc8051_alu1_oc8051_mul1_n12), .Y(oc8051_alu1_oc8051_mul1_n48) );
  OR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u55 ( .A(oc8051_alu1_oc8051_mul1_n11), .B(oc8051_alu1_oc8051_mul1_n48), .Y(oc8051_alu1_oc8051_mul1_n49) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u54 ( .A0(
        oc8051_alu1_oc8051_mul1_n11), .A1(oc8051_alu1_oc8051_mul1_n48), .B0(
        oc8051_alu1_oc8051_mul1_n49), .B1(
        oc8051_alu1_oc8051_mul1_mul_result1_5_), .Y(oc8051_alu1_oc8051_mul1_n8) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u53 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_4_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n10) );
  AND2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u52 ( .A(
        oc8051_alu1_oc8051_mul1_n10), .B(oc8051_alu1_oc8051_mul1_n8), .Y(
        oc8051_alu1_oc8051_mul1_n47) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u51 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1_6_), .Y(oc8051_alu1_oc8051_mul1_n9) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u50 ( .A0(
        oc8051_alu1_oc8051_mul1_n8), .A1(oc8051_alu1_oc8051_mul1_n10), .B0(
        oc8051_alu1_oc8051_mul1_n47), .B1(oc8051_alu1_oc8051_mul1_n9), .Y(
        oc8051_alu1_oc8051_mul1_n6) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u49 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_5_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n7) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u48 ( .A(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_oc8051_mul1_n45) );
  OR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u47 ( .A(oc8051_alu1_oc8051_mul1_n6), 
        .B(oc8051_alu1_oc8051_mul1_n45), .Y(oc8051_alu1_oc8051_mul1_n46) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u46 ( .A0(
        oc8051_alu1_oc8051_mul1_n6), .A1(oc8051_alu1_oc8051_mul1_n45), .B0(
        oc8051_alu1_oc8051_mul1_n46), .B1(
        oc8051_alu1_oc8051_mul1_mul_result1_7_), .Y(
        oc8051_alu1_oc8051_mul1_n41) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u45 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1_8_), .Y(
        oc8051_alu1_oc8051_mul1_n44) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u44 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_6_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n42) );
  XNOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u43 ( .A(
        oc8051_alu1_oc8051_mul1_n41), .B(oc8051_alu1_oc8051_mul1_n44), .C(
        oc8051_alu1_oc8051_mul1_n42), .Y(oc8051_alu1_mulsrc1[0]) );
  AND2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u42 ( .A(
        oc8051_alu1_oc8051_mul1_n42), .B(oc8051_alu1_oc8051_mul1_n41), .Y(
        oc8051_alu1_oc8051_mul1_n43) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u41 ( .A0(
        oc8051_alu1_oc8051_mul1_n41), .A1(oc8051_alu1_oc8051_mul1_n42), .B0(
        oc8051_alu1_oc8051_mul1_n43), .B1(oc8051_alu1_oc8051_mul1_n44), .Y(
        oc8051_alu1_oc8051_mul1_n40) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u40 ( .A(oc8051_alu1_oc8051_mul1_n40), .Y(oc8051_alu1_oc8051_mul1_n36) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u39 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1_9_), .Y(
        oc8051_alu1_oc8051_mul1_n39) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u38 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_7_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n37) );
  XNOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u37 ( .A(
        oc8051_alu1_oc8051_mul1_n36), .B(oc8051_alu1_oc8051_mul1_n39), .C(
        oc8051_alu1_oc8051_mul1_n37), .Y(oc8051_alu1_mulsrc1[1]) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u36 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_8_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n35) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u35 ( .AN(
        oc8051_alu1_oc8051_mul1_n37), .B(oc8051_alu1_oc8051_mul1_n40), .Y(
        oc8051_alu1_oc8051_mul1_n38) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u34 ( .A0(
        oc8051_alu1_oc8051_mul1_n36), .A1(oc8051_alu1_oc8051_mul1_n37), .B0(
        oc8051_alu1_oc8051_mul1_n38), .B1(oc8051_alu1_oc8051_mul1_n39), .Y(
        oc8051_alu1_oc8051_mul1_n34) );
  XNOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u33 ( .A(
        oc8051_alu1_oc8051_mul1_n35), .B(oc8051_alu1_oc8051_mul1_n34), .Y(
        oc8051_alu1_mulsrc1[2]) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u32 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_9_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n33) );
  AND2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u31 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_8_), .B(oc8051_alu1_oc8051_mul1_n34), 
        .Y(oc8051_alu1_oc8051_mul1_n32) );
  XNOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u30 ( .A(
        oc8051_alu1_oc8051_mul1_n33), .B(oc8051_alu1_oc8051_mul1_n32), .Y(
        oc8051_alu1_mulsrc1[3]) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u29 ( .A(
        oc8051_alu1_oc8051_mul1_n32), .B(oc8051_alu1_oc8051_mul1_tmp_mul_9_), 
        .Y(oc8051_alu1_oc8051_mul1_n29) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u28 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_10_), .Y(oc8051_alu1_oc8051_mul1_n30)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u27 ( .A(
        oc8051_alu1_oc8051_mul1_n20), .B(oc8051_alu1_oc8051_mul1_n30), .Y(
        oc8051_alu1_oc8051_mul1_n31) );
  XNOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u26 ( .A(
        oc8051_alu1_oc8051_mul1_n29), .B(oc8051_alu1_oc8051_mul1_n31), .Y(
        oc8051_alu1_mulsrc1[4]) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u25 ( .A(
        oc8051_alu1_oc8051_mul1_n29), .B(oc8051_alu1_oc8051_mul1_n30), .Y(
        oc8051_alu1_oc8051_mul1_n27) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u24 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul_11_), .B(oc8051_alu1_oc8051_mul1_n20), 
        .Y(oc8051_alu1_oc8051_mul1_n28) );
  XOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u23 ( .A(
        oc8051_alu1_oc8051_mul1_n27), .B(oc8051_alu1_oc8051_mul1_n28), .Y(
        oc8051_alu1_mulsrc1[5]) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u22 ( .A(
        oc8051_alu1_oc8051_mul1_n27), .B(oc8051_alu1_oc8051_mul1_tmp_mul_11_), 
        .Y(oc8051_alu1_oc8051_mul1_n24) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_mul1_u21 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_12_), .Y(oc8051_alu1_oc8051_mul1_n23)
         );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u20 ( .A(
        oc8051_alu1_oc8051_mul1_n20), .B(oc8051_alu1_oc8051_mul1_n23), .Y(
        oc8051_alu1_oc8051_mul1_n26) );
  XNOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u19 ( .A(
        oc8051_alu1_oc8051_mul1_n24), .B(oc8051_alu1_oc8051_mul1_n26), .Y(
        oc8051_alu1_mulsrc1[6]) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u18 ( .A(
        oc8051_alu1_oc8051_mul1_tmp_mul_13_), .B(oc8051_alu1_oc8051_mul1_n25), 
        .Y(oc8051_alu1_oc8051_mul1_n21) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_mul1_u17 ( .A(
        oc8051_alu1_oc8051_mul1_n23), .B(oc8051_alu1_oc8051_mul1_n24), .Y(
        oc8051_alu1_oc8051_mul1_n22) );
  XNOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u16 ( .A(
        oc8051_alu1_oc8051_mul1_n21), .B(oc8051_alu1_oc8051_mul1_n22), .Y(
        oc8051_alu1_mulsrc1[7]) );
  NOR2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u15 ( .AN(
        oc8051_alu1_oc8051_mul1_tmp_mul_0_), .B(oc8051_alu1_oc8051_mul1_n20), 
        .Y(oc8051_alu1_oc8051_mul1_n19) );
  XOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u14 ( .A(
        oc8051_alu1_oc8051_mul1_mul_result1_2_), .B(
        oc8051_alu1_oc8051_mul1_n19), .Y(oc8051_alu1_mulsrc2[2]) );
  XOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u13 ( .A(
        oc8051_alu1_oc8051_mul1_n16), .B(oc8051_alu1_oc8051_mul1_n18), .C(
        oc8051_alu1_oc8051_mul1_mul_result1_3_), .Y(oc8051_alu1_mulsrc2[3]) );
  XNOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u12 ( .A(
        oc8051_alu1_oc8051_mul1_n13), .B(oc8051_alu1_oc8051_mul1_n14), .C(
        oc8051_alu1_oc8051_mul1_n15), .Y(oc8051_alu1_mulsrc2[4]) );
  XNOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u11 ( .A(
        oc8051_alu1_oc8051_mul1_n11), .B(
        oc8051_alu1_oc8051_mul1_mul_result1_5_), .C(
        oc8051_alu1_oc8051_mul1_n12), .Y(oc8051_alu1_mulsrc2[5]) );
  XNOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u10 ( .A(
        oc8051_alu1_oc8051_mul1_n8), .B(oc8051_alu1_oc8051_mul1_n9), .C(
        oc8051_alu1_oc8051_mul1_n10), .Y(oc8051_alu1_mulsrc2[6]) );
  XNOR3_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u9 ( .A(oc8051_alu1_oc8051_mul1_n6), .B(oc8051_alu1_oc8051_mul1_mul_result1_7_), .C(oc8051_alu1_oc8051_mul1_n7), 
        .Y(oc8051_alu1_mulsrc2[7]) );
  OR4_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u8 ( .A(oc8051_alu1_mulsrc1[6]), .B(
        oc8051_alu1_mulsrc1[5]), .C(oc8051_alu1_mulsrc1[4]), .D(
        oc8051_alu1_mulsrc1[3]), .Y(oc8051_alu1_oc8051_mul1_n4) );
  OR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u7 ( .A(oc8051_alu1_mulsrc1[1]), .B(
        oc8051_alu1_mulsrc1[2]), .Y(oc8051_alu1_oc8051_mul1_n5) );
  OR4_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u6 ( .A(oc8051_alu1_oc8051_mul1_n4), 
        .B(oc8051_alu1_mulsrc1[7]), .C(oc8051_alu1_mulsrc1[0]), .D(
        oc8051_alu1_oc8051_mul1_n5), .Y(oc8051_alu1_mulov) );
  XOR2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u5 ( .A(oc8051_alu1_n290), .B(
        oc8051_alu1_oc8051_mul1_cycle_0_), .Y(oc8051_alu1_oc8051_mul1_n17) );
  MXIT2_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u4 ( .A(
        oc8051_alu1_oc8051_mul1_cycle_1_), .B(oc8051_alu1_oc8051_mul1_n3), 
        .S0(oc8051_alu1_n290), .Y(oc8051_alu1_oc8051_mul1_n2) );
  NAND2B_X0P5M_A12TS oc8051_alu1_oc8051_mul1_u3 ( .AN(
        oc8051_alu1_oc8051_mul1_n1), .B(oc8051_alu1_oc8051_mul1_n2), .Y(
        oc8051_alu1_oc8051_mul1_n55) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_cycle_reg_0_ ( .D(
        oc8051_alu1_oc8051_mul1_n17), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_cycle_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_cycle_reg_1_ ( .D(
        oc8051_alu1_oc8051_mul1_n55), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_cycle_1_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_9_ ( .D(
        oc8051_alu1_mulsrc1[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_9_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_11_ ( .D(
        oc8051_alu1_mulsrc1[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_11_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_8_ ( .D(
        oc8051_alu1_mulsrc1[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_8_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_0_ ( .D(
        oc8051_alu1_mulsrc2[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_13_ ( .D(
        oc8051_alu1_mulsrc1[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_13_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_7_ ( .D(
        oc8051_alu1_mulsrc2[7]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_7_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_6_ ( .D(
        oc8051_alu1_mulsrc2[6]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_6_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_5_ ( .D(
        oc8051_alu1_mulsrc2[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_5_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_4_ ( .D(
        oc8051_alu1_mulsrc2[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_4_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_3_ ( .D(
        oc8051_alu1_mulsrc2[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_3_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_2_ ( .D(
        oc8051_alu1_mulsrc2[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_2_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_12_ ( .D(
        oc8051_alu1_mulsrc1[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_12_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_10_ ( .D(
        oc8051_alu1_mulsrc1[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_10_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_mul1_tmp_mul_reg_1_ ( .D(
        oc8051_alu1_mulsrc2[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_mul1_tmp_mul_1_) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u47 ( .A(
        oc8051_alu1_oc8051_mul1_n80), .Y(oc8051_alu1_oc8051_mul1_mult_90_n32)
         );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u46 ( .A(
        oc8051_alu1_oc8051_mul1_n70), .Y(oc8051_alu1_oc8051_mul1_mult_90_n33)
         );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u45 ( .A(src1[3]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n28) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u44 ( .A(src1[6]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n25) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u43 ( .A(src1[2]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n29) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u42 ( .A(src1[7]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n24) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u41 ( .A(src1[4]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n27) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u40 ( .A(src1[5]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n26) );
  INV_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u39 ( .A(src1[1]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n30) );
  INV_X0P5M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u38 ( .A(src1[0]), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n31) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u25 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n31), .Y(oc8051_alu1_mulsrc2[0]) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u24 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n30), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n23) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u23 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n29), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n22) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u22 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n28), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n21) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u21 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n27), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n20) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u20 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n26), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n19) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u19 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n25), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n18) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u18 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n33), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n24), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n17) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u17 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n31), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n16) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u16 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n30), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n15) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u15 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n29), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n14) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u14 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n28), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n13) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u13 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n27), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n12) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u12 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n26), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n11) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u11 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n25), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n10) );
  NOR2_X1A_A12TS oc8051_alu1_oc8051_mul1_mult_90_u10 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n32), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n24), .Y(
        oc8051_alu1_oc8051_mul1_mult_90_n9) );
  ADDH_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u9 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n23), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n16), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n8), .S(oc8051_alu1_mulsrc2[1]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u8 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n22), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n15), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n8), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n7), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_2_) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u7 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n21), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n14), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n7), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n6), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_3_) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u6 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n20), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n13), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n6), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n5), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_4_) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u5 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n19), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n12), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n5), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n4), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_5_) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u4 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n18), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n11), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n4), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n3), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_6_) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u3 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n17), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n10), .CI(
        oc8051_alu1_oc8051_mul1_mult_90_n3), .CO(
        oc8051_alu1_oc8051_mul1_mult_90_n2), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_7_) );
  ADDH_X1M_A12TS oc8051_alu1_oc8051_mul1_mult_90_u2 ( .A(
        oc8051_alu1_oc8051_mul1_mult_90_n2), .B(
        oc8051_alu1_oc8051_mul1_mult_90_n9), .CO(
        oc8051_alu1_oc8051_mul1_mul_result1_9_), .S(
        oc8051_alu1_oc8051_mul1_mul_result1_8_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u67 ( .A(src2[0]), .Y(
        oc8051_alu1_oc8051_div1_n7) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u66 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .B(oc8051_alu1_oc8051_div1_cycle_0_), .Y(oc8051_alu1_oc8051_div1_n18) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u65 ( .A(oc8051_alu1_oc8051_div1_n7), .B(oc8051_alu1_oc8051_div1_n18), .Y(oc8051_alu1_oc8051_div1_cmp1_1_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u64 ( .A(src2[1]), .Y(
        oc8051_alu1_oc8051_div1_n8) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u63 ( .A(
        oc8051_alu1_oc8051_div1_n18), .B(oc8051_alu1_oc8051_div1_n8), .Y(
        oc8051_alu1_oc8051_div1_cmp1_2_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u62 ( .A(src2[2]), .Y(
        oc8051_alu1_oc8051_div1_n9) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u61 ( .A(
        oc8051_alu1_oc8051_div1_cycle_0_), .Y(oc8051_alu1_oc8051_div1_n23) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u60 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .B(oc8051_alu1_oc8051_div1_n23), 
        .Y(oc8051_alu1_oc8051_div1_n3) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u59 ( .A0(
        oc8051_alu1_oc8051_div1_n9), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n3), .B1(oc8051_alu1_oc8051_div1_n7), .Y(
        oc8051_alu1_oc8051_div1_cmp1_3_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u58 ( .A(src2[3]), .Y(
        oc8051_alu1_oc8051_div1_n10) );
  OAI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u57 ( .A0(
        oc8051_alu1_oc8051_div1_n10), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n8), .B1(oc8051_alu1_oc8051_div1_n3), .Y(
        oc8051_alu1_oc8051_div1_cmp1_4_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u56 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .Y(oc8051_alu1_oc8051_div1_n24) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u55 ( .A(
        oc8051_alu1_oc8051_div1_cycle_0_), .B(oc8051_alu1_oc8051_div1_n24), 
        .Y(oc8051_alu1_oc8051_div1_n30) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u54 ( .A(src2[4]), .Y(
        oc8051_alu1_oc8051_div1_n11) );
  OAI222_X0P5M_A12TS oc8051_alu1_oc8051_div1_u53 ( .A0(
        oc8051_alu1_oc8051_div1_n9), .A1(oc8051_alu1_oc8051_div1_n3), .B0(
        oc8051_alu1_oc8051_div1_n30), .B1(oc8051_alu1_oc8051_div1_n7), .C0(
        oc8051_alu1_oc8051_div1_n11), .C1(oc8051_alu1_oc8051_div1_n18), .Y(
        oc8051_alu1_oc8051_div1_cmp1_5_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u52 ( .A(src2[5]), .Y(
        oc8051_alu1_oc8051_div1_n12) );
  OAI222_X0P5M_A12TS oc8051_alu1_oc8051_div1_u51 ( .A0(
        oc8051_alu1_oc8051_div1_n10), .A1(oc8051_alu1_oc8051_div1_n3), .B0(
        oc8051_alu1_oc8051_div1_n8), .B1(oc8051_alu1_oc8051_div1_n30), .C0(
        oc8051_alu1_oc8051_div1_n12), .C1(oc8051_alu1_oc8051_div1_n18), .Y(
        oc8051_alu1_oc8051_div1_cmp1_6_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u50 ( .A(src2[6]), .Y(
        oc8051_alu1_oc8051_div1_n13) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u49 ( .A(
        oc8051_alu1_oc8051_div1_n23), .B(oc8051_alu1_oc8051_div1_n24), .Y(
        oc8051_alu1_oc8051_div1_n15) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u48 ( .A(oc8051_alu1_oc8051_div1_n30), .Y(oc8051_alu1_oc8051_div1_n4) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u47 ( .A(oc8051_alu1_oc8051_div1_n3), 
        .Y(oc8051_alu1_oc8051_div1_n28) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u46 ( .A0(
        oc8051_alu1_oc8051_div1_n4), .A1(src2[2]), .B0(src2[4]), .B1(
        oc8051_alu1_oc8051_div1_n28), .Y(oc8051_alu1_oc8051_div1_n29) );
  OAI221_X0P5M_A12TS oc8051_alu1_oc8051_div1_u45 ( .A0(
        oc8051_alu1_oc8051_div1_n13), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n15), .B1(oc8051_alu1_oc8051_div1_n7), .C0(
        oc8051_alu1_oc8051_div1_n29), .Y(oc8051_alu1_oc8051_div1_cmp1_7_) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u44 ( .A(src2[7]), .Y(
        oc8051_alu1_oc8051_div1_n14) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u43 ( .A0(
        oc8051_alu1_oc8051_div1_n4), .A1(src2[3]), .B0(
        oc8051_alu1_oc8051_div1_n28), .B1(src2[5]), .Y(
        oc8051_alu1_oc8051_div1_n27) );
  OAI221_X0P5M_A12TS oc8051_alu1_oc8051_div1_u42 ( .A0(
        oc8051_alu1_oc8051_div1_n14), .A1(oc8051_alu1_oc8051_div1_n18), .B0(
        oc8051_alu1_oc8051_div1_n15), .B1(oc8051_alu1_oc8051_div1_n8), .C0(
        oc8051_alu1_oc8051_div1_n27), .Y(oc8051_alu1_oc8051_div1_cmp0_7_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u41 ( .A(src1[0]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[0]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_sub1[0]) );
  AOI22_X0P5M_A12TS oc8051_alu1_oc8051_div1_u40 ( .A0(src2[5]), .A1(
        oc8051_alu1_oc8051_div1_n23), .B0(src2[3]), .B1(
        oc8051_alu1_oc8051_div1_n24), .Y(oc8051_alu1_oc8051_div1_n19) );
  INV_X0P5B_A12TS oc8051_alu1_oc8051_div1_u39 ( .A(oc8051_alu1_oc8051_div1_n15), .Y(oc8051_alu1_oc8051_div1_n21) );
  AOI21_X0P5M_A12TS oc8051_alu1_oc8051_div1_u38 ( .A0(
        oc8051_alu1_oc8051_div1_n11), .A1(oc8051_alu1_oc8051_div1_n12), .B0(
        oc8051_alu1_oc8051_div1_cycle_1_), .Y(oc8051_alu1_oc8051_div1_n22) );
  AOI221_X0P5M_A12TS oc8051_alu1_oc8051_div1_u37 ( .A0(
        oc8051_alu1_oc8051_div1_n18), .A1(src2[6]), .B0(
        oc8051_alu1_oc8051_div1_n21), .B1(src2[2]), .C0(
        oc8051_alu1_oc8051_div1_n22), .Y(oc8051_alu1_oc8051_div1_n16) );
  AOI211_X0P5M_A12TS oc8051_alu1_oc8051_div1_u36 ( .A0(src2[1]), .A1(
        oc8051_alu1_oc8051_div1_n21), .B0(oc8051_alu1_oc8051_div1_sub1[8]), 
        .C0(src2[7]), .Y(oc8051_alu1_oc8051_div1_n20) );
  AND3_X0P5M_A12TS oc8051_alu1_oc8051_div1_u35 ( .A(
        oc8051_alu1_oc8051_div1_n19), .B(oc8051_alu1_oc8051_div1_n16), .C(
        oc8051_alu1_oc8051_div1_n20), .Y(oc8051_alu1_divsrc2[1]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u34 ( .A(
        oc8051_alu1_oc8051_div1_sub1[0]), .B(oc8051_alu1_oc8051_div1_sub1[0]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_0_) );
  AOI21_X0P5M_A12TS oc8051_alu1_oc8051_div1_u33 ( .A0(src2[7]), .A1(
        oc8051_alu1_oc8051_div1_n18), .B0(oc8051_alu1_oc8051_div1_sub0[8]), 
        .Y(oc8051_alu1_oc8051_div1_n17) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u32 ( .A(
        oc8051_alu1_oc8051_div1_rem1_0_), .B(oc8051_alu1_oc8051_div1_sub0[0]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[0]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u31 ( .A(src1[1]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[1]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_1_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u30 ( .A(
        oc8051_alu1_oc8051_div1_rem2_1_), .B(oc8051_alu1_oc8051_div1_sub1[1]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_1_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u29 ( .A(
        oc8051_alu1_oc8051_div1_rem1_1_), .B(oc8051_alu1_oc8051_div1_sub0[1]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[1]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u28 ( .A(src1[2]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[2]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_2_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u27 ( .A(
        oc8051_alu1_oc8051_div1_rem2_2_), .B(oc8051_alu1_oc8051_div1_sub1[2]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_2_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u26 ( .A(
        oc8051_alu1_oc8051_div1_rem1_2_), .B(oc8051_alu1_oc8051_div1_sub0[2]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[2]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u25 ( .A(src1[3]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[3]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_3_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u24 ( .A(
        oc8051_alu1_oc8051_div1_rem2_3_), .B(oc8051_alu1_oc8051_div1_sub1[3]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_3_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u23 ( .A(
        oc8051_alu1_oc8051_div1_rem1_3_), .B(oc8051_alu1_oc8051_div1_sub0[3]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[3]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u22 ( .A(src1[4]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[4]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_4_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u21 ( .A(
        oc8051_alu1_oc8051_div1_rem2_4_), .B(oc8051_alu1_oc8051_div1_sub1[4]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_4_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u20 ( .A(
        oc8051_alu1_oc8051_div1_rem1_4_), .B(oc8051_alu1_oc8051_div1_sub0[4]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[4]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u19 ( .A(src1[5]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[5]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_5_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u18 ( .A(
        oc8051_alu1_oc8051_div1_rem2_5_), .B(oc8051_alu1_oc8051_div1_sub1[5]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_5_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u17 ( .A(
        oc8051_alu1_oc8051_div1_rem1_5_), .B(oc8051_alu1_oc8051_div1_sub0[5]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[5]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u16 ( .A(src1[6]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[6]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_6_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u15 ( .A(
        oc8051_alu1_oc8051_div1_rem2_6_), .B(oc8051_alu1_oc8051_div1_sub1[6]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_6_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u14 ( .A(
        oc8051_alu1_oc8051_div1_rem1_6_), .B(oc8051_alu1_oc8051_div1_sub0[6]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[6]) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u13 ( .A(src1[7]), .B(
        oc8051_alu1_oc8051_div1_tmp_rem[7]), .S0(oc8051_alu1_oc8051_div1_n15), 
        .Y(oc8051_alu1_oc8051_div1_rem2_7_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u12 ( .A(
        oc8051_alu1_oc8051_div1_rem2_7_), .B(oc8051_alu1_oc8051_div1_sub1[7]), 
        .S0(oc8051_alu1_divsrc2[1]), .Y(oc8051_alu1_oc8051_div1_rem1_7_) );
  MXT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u11 ( .A(
        oc8051_alu1_oc8051_div1_rem1_7_), .B(oc8051_alu1_oc8051_div1_sub0[7]), 
        .S0(oc8051_alu1_divsrc2[0]), .Y(oc8051_alu1_divsrc1[7]) );
  NAND4_X0P5A_A12TS oc8051_alu1_oc8051_div1_u10 ( .A(
        oc8051_alu1_oc8051_div1_n11), .B(oc8051_alu1_oc8051_div1_n12), .C(
        oc8051_alu1_oc8051_div1_n13), .D(oc8051_alu1_oc8051_div1_n14), .Y(
        oc8051_alu1_oc8051_div1_n5) );
  NAND4_X0P5A_A12TS oc8051_alu1_oc8051_div1_u9 ( .A(oc8051_alu1_oc8051_div1_n7), .B(oc8051_alu1_oc8051_div1_n8), .C(oc8051_alu1_oc8051_div1_n9), .D(
        oc8051_alu1_oc8051_div1_n10), .Y(oc8051_alu1_oc8051_div1_n6) );
  NOR2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u8 ( .A(oc8051_alu1_oc8051_div1_n5), 
        .B(oc8051_alu1_oc8051_div1_n6), .Y(oc8051_alu1_divov) );
  MXIT2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u7 ( .A(
        oc8051_alu1_oc8051_div1_cycle_1_), .B(oc8051_alu1_oc8051_div1_n4), 
        .S0(oc8051_alu1_n288), .Y(oc8051_alu1_oc8051_div1_n2) );
  NAND2_X0P5A_A12TS oc8051_alu1_oc8051_div1_u6 ( .A(oc8051_alu1_oc8051_div1_n2), .B(oc8051_alu1_oc8051_div1_n3), .Y(oc8051_alu1_oc8051_div1_n25) );
  XOR2_X0P5M_A12TS oc8051_alu1_oc8051_div1_u5 ( .A(oc8051_alu1_n288), .B(
        oc8051_alu1_oc8051_div1_cycle_0_), .Y(oc8051_alu1_oc8051_div1_n26) );
  TIELO_X1M_A12TS oc8051_alu1_oc8051_div1_u4 ( .Y(
        oc8051_alu1_oc8051_div1_cmp1_0_) );
  OA211_X1M_A12TS oc8051_alu1_oc8051_div1_u3 ( .A0(oc8051_alu1_oc8051_div1_n15), .A1(oc8051_alu1_oc8051_div1_n10), .B0(oc8051_alu1_oc8051_div1_n16), .C0(
        oc8051_alu1_oc8051_div1_n17), .Y(oc8051_alu1_divsrc2[0]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_cycle_reg_1_ ( .D(
        oc8051_alu1_oc8051_div1_n25), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_cycle_1_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_cycle_reg_0_ ( .D(
        oc8051_alu1_oc8051_div1_n26), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_cycle_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_1_ ( .D(
        oc8051_alu1_divsrc2[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_0_ ( .D(
        oc8051_alu1_divsrc2[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_3_ ( .D(
        oc8051_alu1_divsrc2[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_2_ ( .D(
        oc8051_alu1_divsrc2[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_5_ ( .D(
        oc8051_alu1_divsrc2[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_div_reg_4_ ( .D(
        oc8051_alu1_divsrc2[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_divsrc2[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_2_ ( .D(
        oc8051_alu1_divsrc1[2]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_3_ ( .D(
        oc8051_alu1_divsrc1[3]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_4_ ( .D(
        oc8051_alu1_divsrc1[4]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_5_ ( .D(
        oc8051_alu1_divsrc1[5]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_6_ ( .D(
        oc8051_alu1_divsrc1[6]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_7_ ( .D(
        oc8051_alu1_divsrc1[7]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_1_ ( .D(
        oc8051_alu1_divsrc1[1]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu1_oc8051_div1_tmp_rem_reg_0_ ( .D(
        oc8051_alu1_divsrc1[0]), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_alu1_oc8051_div1_tmp_rem[0]) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u11 ( .A(
        oc8051_alu1_oc8051_div1_cmp0_7_), .Y(oc8051_alu1_oc8051_div1_sub_98_n3) );
  OR2_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u10 ( .A(
        oc8051_alu1_oc8051_div1_rem1_0_), .B(
        oc8051_alu1_oc8051_div1_sub_98_n10), .Y(
        oc8051_alu1_oc8051_div1_sub_98_n1) );
  XNOR2_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u9 ( .A(
        oc8051_alu1_oc8051_div1_sub_98_n10), .B(
        oc8051_alu1_oc8051_div1_rem1_0_), .Y(oc8051_alu1_oc8051_div1_sub0[0])
         );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u8 ( .A(
        oc8051_alu1_oc8051_div1_sub_98_carry[8]), .Y(
        oc8051_alu1_oc8051_div1_sub0[8]) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u7 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_7_), .Y(oc8051_alu1_oc8051_div1_sub_98_n4) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u6 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_6_), .Y(oc8051_alu1_oc8051_div1_sub_98_n5) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u5 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_5_), .Y(oc8051_alu1_oc8051_div1_sub_98_n6) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u4 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_4_), .Y(oc8051_alu1_oc8051_div1_sub_98_n7) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u3 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_3_), .Y(oc8051_alu1_oc8051_div1_sub_98_n8) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_1_), .Y(
        oc8051_alu1_oc8051_div1_sub_98_n10) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u1 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_2_), .Y(oc8051_alu1_oc8051_div1_sub_98_n9) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_1 ( .A(
        oc8051_alu1_oc8051_div1_rem1_1_), .B(oc8051_alu1_oc8051_div1_sub_98_n9), .CI(oc8051_alu1_oc8051_div1_sub_98_n1), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[2]), .S(
        oc8051_alu1_oc8051_div1_sub0[1]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_2 ( .A(
        oc8051_alu1_oc8051_div1_rem1_2_), .B(oc8051_alu1_oc8051_div1_sub_98_n8), .CI(oc8051_alu1_oc8051_div1_sub_98_carry[2]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[3]), .S(
        oc8051_alu1_oc8051_div1_sub0[2]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_3 ( .A(
        oc8051_alu1_oc8051_div1_rem1_3_), .B(oc8051_alu1_oc8051_div1_sub_98_n7), .CI(oc8051_alu1_oc8051_div1_sub_98_carry[3]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[4]), .S(
        oc8051_alu1_oc8051_div1_sub0[3]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_4 ( .A(
        oc8051_alu1_oc8051_div1_rem1_4_), .B(oc8051_alu1_oc8051_div1_sub_98_n6), .CI(oc8051_alu1_oc8051_div1_sub_98_carry[4]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[5]), .S(
        oc8051_alu1_oc8051_div1_sub0[4]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_5 ( .A(
        oc8051_alu1_oc8051_div1_rem1_5_), .B(oc8051_alu1_oc8051_div1_sub_98_n5), .CI(oc8051_alu1_oc8051_div1_sub_98_carry[5]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[6]), .S(
        oc8051_alu1_oc8051_div1_sub0[5]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_6 ( .A(
        oc8051_alu1_oc8051_div1_rem1_6_), .B(oc8051_alu1_oc8051_div1_sub_98_n4), .CI(oc8051_alu1_oc8051_div1_sub_98_carry[6]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[7]), .S(
        oc8051_alu1_oc8051_div1_sub0[6]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_98_u2_7 ( .A(
        oc8051_alu1_oc8051_div1_rem1_7_), .B(oc8051_alu1_oc8051_div1_sub_98_n3), .CI(oc8051_alu1_oc8051_div1_sub_98_carry[7]), .CO(
        oc8051_alu1_oc8051_div1_sub_98_carry[8]), .S(
        oc8051_alu1_oc8051_div1_sub0[7]) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u10 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_7_), .Y(oc8051_alu1_oc8051_div1_sub_94_n3) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u9 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_3_), .Y(oc8051_alu1_oc8051_div1_sub_94_n7) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u8 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_6_), .Y(oc8051_alu1_oc8051_div1_sub_94_n4) );
  OR2_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u7 ( .A(
        oc8051_alu1_oc8051_div1_rem2_1_), .B(oc8051_alu1_oc8051_div1_sub_94_n9), .Y(oc8051_alu1_oc8051_div1_sub_94_n1) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u6 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_4_), .Y(oc8051_alu1_oc8051_div1_sub_94_n6) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u5 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_5_), .Y(oc8051_alu1_oc8051_div1_sub_94_n5) );
  XNOR2_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u4 ( .A(
        oc8051_alu1_oc8051_div1_sub_94_n9), .B(oc8051_alu1_oc8051_div1_rem2_1_), .Y(oc8051_alu1_oc8051_div1_sub1[1]) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u3 ( .A(
        oc8051_alu1_oc8051_div1_sub_94_carry[8]), .Y(
        oc8051_alu1_oc8051_div1_sub1[8]) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_1_), .Y(oc8051_alu1_oc8051_div1_sub_94_n9) );
  INV_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u1 ( .A(
        oc8051_alu1_oc8051_div1_cmp1_2_), .Y(oc8051_alu1_oc8051_div1_sub_94_n8) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_2 ( .A(
        oc8051_alu1_oc8051_div1_rem2_2_), .B(oc8051_alu1_oc8051_div1_sub_94_n8), .CI(oc8051_alu1_oc8051_div1_sub_94_n1), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[3]), .S(
        oc8051_alu1_oc8051_div1_sub1[2]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_3 ( .A(
        oc8051_alu1_oc8051_div1_rem2_3_), .B(oc8051_alu1_oc8051_div1_sub_94_n7), .CI(oc8051_alu1_oc8051_div1_sub_94_carry[3]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[4]), .S(
        oc8051_alu1_oc8051_div1_sub1[3]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_4 ( .A(
        oc8051_alu1_oc8051_div1_rem2_4_), .B(oc8051_alu1_oc8051_div1_sub_94_n6), .CI(oc8051_alu1_oc8051_div1_sub_94_carry[4]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[5]), .S(
        oc8051_alu1_oc8051_div1_sub1[4]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_5 ( .A(
        oc8051_alu1_oc8051_div1_rem2_5_), .B(oc8051_alu1_oc8051_div1_sub_94_n5), .CI(oc8051_alu1_oc8051_div1_sub_94_carry[5]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[6]), .S(
        oc8051_alu1_oc8051_div1_sub1[5]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_6 ( .A(
        oc8051_alu1_oc8051_div1_rem2_6_), .B(oc8051_alu1_oc8051_div1_sub_94_n4), .CI(oc8051_alu1_oc8051_div1_sub_94_carry[6]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[7]), .S(
        oc8051_alu1_oc8051_div1_sub1[6]) );
  ADDF_X1M_A12TS oc8051_alu1_oc8051_div1_sub_94_u2_7 ( .A(
        oc8051_alu1_oc8051_div1_rem2_7_), .B(oc8051_alu1_oc8051_div1_sub_94_n3), .CI(oc8051_alu1_oc8051_div1_sub_94_carry[7]), .CO(
        oc8051_alu1_oc8051_div1_sub_94_carry[8]), .S(
        oc8051_alu1_oc8051_div1_sub1[7]) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u30 ( .A(src1[3]), .B(
        oc8051_alu1_sub_205_n5), .Y(oc8051_alu1_dec[3]) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u29 ( .A(oc8051_alu1_sub_205_n10), .B(
        src2[5]), .Y(oc8051_alu1_sub_205_n13) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u28 ( .A(oc8051_alu1_sub_205_n8), .B(
        src2[3]), .Y(oc8051_alu1_sub_205_n12) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u27 ( .A(oc8051_alu1_sub_205_n9), .B(
        src2[1]), .Y(oc8051_alu1_sub_205_n11) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u26 ( .A(oc8051_alu1_sub_205_n12), .B(
        src2[4]), .Y(oc8051_alu1_sub_205_n10) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u25 ( .A(oc8051_alu1_sub_205_n4), .B(
        src2[0]), .Y(oc8051_alu1_sub_205_n9) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u24 ( .A(oc8051_alu1_sub_205_n11), .B(
        src2[2]), .Y(oc8051_alu1_sub_205_n8) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u23 ( .A(oc8051_alu1_sub_205_n5), .B(
        src1[3]), .Y(oc8051_alu1_sub_205_n7) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u22 ( .A(oc8051_alu1_sub_205_n2), .B(
        src1[6]), .Y(oc8051_alu1_sub_205_n6) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u21 ( .A(oc8051_alu1_sub_205_n1), .B(
        src1[2]), .Y(oc8051_alu1_sub_205_n5) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u20 ( .A(oc8051_alu1_sub_205_n6), .B(
        src1[7]), .Y(oc8051_alu1_sub_205_n4) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u19 ( .A(oc8051_alu1_sub_205_n7), .B(
        src1[4]), .Y(oc8051_alu1_sub_205_n3) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u18 ( .A(oc8051_alu1_sub_205_n3), .B(
        src1[5]), .Y(oc8051_alu1_sub_205_n2) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u17 ( .A(src1[2]), .B(
        oc8051_alu1_sub_205_n1), .Y(oc8051_alu1_dec[2]) );
  INV_X0P5M_A12TS oc8051_alu1_sub_205_u16 ( .A(src1[0]), .Y(oc8051_alu1_dec[0]) );
  OR2_X1M_A12TS oc8051_alu1_sub_205_u15 ( .A(src1[0]), .B(src1[1]), .Y(
        oc8051_alu1_sub_205_n1) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u14 ( .A(src1[6]), .B(
        oc8051_alu1_sub_205_n2), .Y(oc8051_alu1_dec[6]) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u13 ( .A(src1[7]), .B(
        oc8051_alu1_sub_205_n6), .Y(oc8051_alu1_dec[7]) );
  NOR2_X1A_A12TS oc8051_alu1_sub_205_u12 ( .A(oc8051_alu1_sub_205_n13), .B(
        src2[6]), .Y(oc8051_alu1_sub_205_n14) );
  XOR2_X1M_A12TS oc8051_alu1_sub_205_u11 ( .A(src2[7]), .B(
        oc8051_alu1_sub_205_n14), .Y(oc8051_alu1_dec[15]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u10 ( .A(src2[5]), .B(
        oc8051_alu1_sub_205_n10), .Y(oc8051_alu1_dec[13]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u9 ( .A(src2[3]), .B(
        oc8051_alu1_sub_205_n8), .Y(oc8051_alu1_dec[11]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u8 ( .A(src2[1]), .B(
        oc8051_alu1_sub_205_n9), .Y(oc8051_alu1_dec[9]) );
  XNOR2_X0P5M_A12TS oc8051_alu1_sub_205_u7 ( .A(src1[5]), .B(
        oc8051_alu1_sub_205_n3), .Y(oc8051_alu1_dec[5]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u6 ( .A(src2[4]), .B(
        oc8051_alu1_sub_205_n12), .Y(oc8051_alu1_dec[12]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u5 ( .A(src2[0]), .B(
        oc8051_alu1_sub_205_n4), .Y(oc8051_alu1_dec[8]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u4 ( .A(src2[6]), .B(
        oc8051_alu1_sub_205_n13), .Y(oc8051_alu1_dec[14]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u3 ( .A(src2[2]), .B(
        oc8051_alu1_sub_205_n11), .Y(oc8051_alu1_dec[10]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u2 ( .A(src1[4]), .B(
        oc8051_alu1_sub_205_n7), .Y(oc8051_alu1_dec[4]) );
  XNOR2_X1M_A12TS oc8051_alu1_sub_205_u1 ( .A(src1[1]), .B(src1[0]), .Y(
        oc8051_alu1_dec[1]) );
  XOR2_X0P5M_A12TS oc8051_alu1_add_204_u2 ( .A(oc8051_alu1_add_204_carry[15]), 
        .B(src2[7]), .Y(oc8051_alu1_inc[15]) );
  INV_X1M_A12TS oc8051_alu1_add_204_u1 ( .A(src1[0]), .Y(oc8051_alu1_inc[0])
         );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_1 ( .A(src1[1]), .B(src1[0]), .CO(
        oc8051_alu1_add_204_carry[2]), .S(oc8051_alu1_inc[1]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_5 ( .A(src1[5]), .B(
        oc8051_alu1_add_204_carry[5]), .CO(oc8051_alu1_add_204_carry[6]), .S(
        oc8051_alu1_inc[5]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_4 ( .A(src1[4]), .B(
        oc8051_alu1_add_204_carry[4]), .CO(oc8051_alu1_add_204_carry[5]), .S(
        oc8051_alu1_inc[4]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_7 ( .A(src1[7]), .B(
        oc8051_alu1_add_204_carry[7]), .CO(oc8051_alu1_add_204_carry[8]), .S(
        oc8051_alu1_inc[7]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_2 ( .A(src1[2]), .B(
        oc8051_alu1_add_204_carry[2]), .CO(oc8051_alu1_add_204_carry[3]), .S(
        oc8051_alu1_inc[2]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_6 ( .A(src1[6]), .B(
        oc8051_alu1_add_204_carry[6]), .CO(oc8051_alu1_add_204_carry[7]), .S(
        oc8051_alu1_inc[6]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_3 ( .A(src1[3]), .B(
        oc8051_alu1_add_204_carry[3]), .CO(oc8051_alu1_add_204_carry[4]), .S(
        oc8051_alu1_inc[3]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_10 ( .A(src2[2]), .B(
        oc8051_alu1_add_204_carry[10]), .CO(oc8051_alu1_add_204_carry[11]), 
        .S(oc8051_alu1_inc[10]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_8 ( .A(src2[0]), .B(
        oc8051_alu1_add_204_carry[8]), .CO(oc8051_alu1_add_204_carry[9]), .S(
        oc8051_alu1_inc[8]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_12 ( .A(src2[4]), .B(
        oc8051_alu1_add_204_carry[12]), .CO(oc8051_alu1_add_204_carry[13]), 
        .S(oc8051_alu1_inc[12]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_9 ( .A(src2[1]), .B(
        oc8051_alu1_add_204_carry[9]), .CO(oc8051_alu1_add_204_carry[10]), .S(
        oc8051_alu1_inc[9]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_11 ( .A(src2[3]), .B(
        oc8051_alu1_add_204_carry[11]), .CO(oc8051_alu1_add_204_carry[12]), 
        .S(oc8051_alu1_inc[11]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_13 ( .A(src2[5]), .B(
        oc8051_alu1_add_204_carry[13]), .CO(oc8051_alu1_add_204_carry[14]), 
        .S(oc8051_alu1_inc[13]) );
  ADDH_X1M_A12TS oc8051_alu1_add_204_u1_1_14 ( .A(src2[6]), .B(
        oc8051_alu1_add_204_carry[14]), .CO(oc8051_alu1_add_204_carry[15]), 
        .S(oc8051_alu1_inc[14]) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u110 ( .A(oc8051_ram_top1_rd_data_m[2]), 
        .B(oc8051_ram_top1_wr_data_r[2]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n56) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u109 ( .A(oc8051_ram_top1_rd_data_m[0]), 
        .B(oc8051_ram_top1_wr_data_r[0]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n58) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u108 ( .A(oc8051_ram_top1_rd_data_m[3]), 
        .B(oc8051_ram_top1_wr_data_r[3]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n55) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u107 ( .A(oc8051_ram_top1_rd_data_m[1]), 
        .B(oc8051_ram_top1_wr_data_r[1]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n57) );
  INV_X0P5B_A12TS oc8051_ram_top1_u106 ( .A(oc8051_ram_top1_n270), .Y(
        oc8051_ram_top1_n48) );
  MXT4_X0P5M_A12TS oc8051_ram_top1_u105 ( .A(oc8051_ram_top1_n56), .B(
        oc8051_ram_top1_n58), .C(oc8051_ram_top1_n55), .D(oc8051_ram_top1_n57), 
        .S0(oc8051_ram_top1_n48), .S1(oc8051_ram_top1_n260), .Y(
        oc8051_ram_top1_n74) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u104 ( .A(oc8051_ram_top1_rd_data_m[6]), 
        .B(oc8051_ram_top1_wr_data_r[6]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n51) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u103 ( .A(oc8051_ram_top1_rd_data_m[4]), 
        .B(oc8051_ram_top1_wr_data_r[4]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n54) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u102 ( .A(oc8051_ram_top1_rd_data_m[7]), 
        .B(oc8051_ram_top1_wr_data_r[7]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n50) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u101 ( .A(oc8051_ram_top1_rd_data_m[5]), 
        .B(oc8051_ram_top1_wr_data_r[5]), .S0(oc8051_ram_top1_rd_en_r), .Y(
        oc8051_ram_top1_n52) );
  MXT4_X0P5M_A12TS oc8051_ram_top1_u100 ( .A(oc8051_ram_top1_n51), .B(
        oc8051_ram_top1_n54), .C(oc8051_ram_top1_n50), .D(oc8051_ram_top1_n52), 
        .S0(oc8051_ram_top1_n48), .S1(oc8051_ram_top1_n260), .Y(
        oc8051_ram_top1_n75) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_u99 ( .A(oc8051_ram_top1_n74), .B(
        oc8051_ram_top1_n75), .S0(oc8051_ram_top1_n280), .Y(bit_data) );
  INV_X0P5B_A12TS oc8051_ram_top1_u98 ( .A(oc8051_ram_top1_bit_addr_r), .Y(
        oc8051_ram_top1_n13) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u97 ( .A(oc8051_ram_top1_n13), .B(
        wr_addr[7]), .Y(oc8051_ram_top1_n68) );
  AO22_X0P5M_A12TS oc8051_ram_top1_u96 ( .A0(wr_addr[1]), .A1(
        oc8051_ram_top1_n13), .B0(oc8051_ram_top1_n68), .B1(wr_addr[4]), .Y(
        oc8051_ram_top1_wr_addr_m_1_) );
  INV_X0P5B_A12TS oc8051_ram_top1_u95 ( .A(bit_addr_o), .Y(oc8051_ram_top1_n71) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u94 ( .A(oc8051_ram_top1_n71), .B(
        rd_addr[7]), .Y(oc8051_ram_top1_n67) );
  AO22_X0P5M_A12TS oc8051_ram_top1_u93 ( .A0(rd_addr[1]), .A1(
        oc8051_ram_top1_n71), .B0(oc8051_ram_top1_n67), .B1(rd_addr[4]), .Y(
        oc8051_ram_top1_rd_addr_m_1_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u92 ( .A(oc8051_ram_top1_wr_addr_m_1_), 
        .B(oc8051_ram_top1_rd_addr_m_1_), .Y(oc8051_ram_top1_n72) );
  AO22_X0P5M_A12TS oc8051_ram_top1_u91 ( .A0(wr_addr[0]), .A1(
        oc8051_ram_top1_n13), .B0(wr_addr[3]), .B1(oc8051_ram_top1_n68), .Y(
        oc8051_ram_top1_wr_addr_m_0_) );
  AO22_X0P5M_A12TS oc8051_ram_top1_u90 ( .A0(rd_addr[0]), .A1(
        oc8051_ram_top1_n71), .B0(rd_addr[3]), .B1(oc8051_ram_top1_n67), .Y(
        oc8051_ram_top1_rd_addr_m_0_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u89 ( .A(oc8051_ram_top1_wr_addr_m_0_), 
        .B(oc8051_ram_top1_rd_addr_m_0_), .Y(oc8051_ram_top1_n73) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u88 ( .A(oc8051_ram_top1_n72), .B(n_0_net_), .C(oc8051_ram_top1_n73), .Y(oc8051_ram_top1_n59) );
  AO22_X0P5M_A12TS oc8051_ram_top1_u87 ( .A0(wr_addr[2]), .A1(
        oc8051_ram_top1_n13), .B0(wr_addr[5]), .B1(oc8051_ram_top1_n68), .Y(
        oc8051_ram_top1_wr_addr_m_2_) );
  AO22_X0P5M_A12TS oc8051_ram_top1_u86 ( .A0(rd_addr[2]), .A1(
        oc8051_ram_top1_n71), .B0(rd_addr[5]), .B1(oc8051_ram_top1_n67), .Y(
        oc8051_ram_top1_rd_addr_m_2_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u85 ( .A(oc8051_ram_top1_wr_addr_m_2_), 
        .B(oc8051_ram_top1_rd_addr_m_2_), .Y(oc8051_ram_top1_n60) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u84 ( .A(rd_addr[7]), .B(wr_addr[7]), .Y(
        oc8051_ram_top1_n61) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_u83 ( .AN(wr_addr[6]), .B(
        oc8051_ram_top1_n68), .Y(oc8051_ram_top1_wr_addr_m_6_) );
  INV_X0P5B_A12TS oc8051_ram_top1_u82 ( .A(oc8051_ram_top1_n67), .Y(
        oc8051_ram_top1_n69) );
  AND2_X0P5M_A12TS oc8051_ram_top1_u81 ( .A(rd_addr[6]), .B(
        oc8051_ram_top1_n69), .Y(oc8051_ram_top1_rd_addr_m_6_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u80 ( .A(oc8051_ram_top1_wr_addr_m_6_), 
        .B(oc8051_ram_top1_rd_addr_m_6_), .Y(oc8051_ram_top1_n63) );
  INV_X0P5B_A12TS oc8051_ram_top1_u79 ( .A(oc8051_ram_top1_n68), .Y(
        oc8051_ram_top1_n70) );
  NAND2B_X0P5M_A12TS oc8051_ram_top1_u78 ( .AN(wr_addr[5]), .B(
        oc8051_ram_top1_n70), .Y(oc8051_ram_top1_wr_addr_m_5_) );
  OR2_X0P5M_A12TS oc8051_ram_top1_u77 ( .A(rd_addr[5]), .B(oc8051_ram_top1_n67), .Y(oc8051_ram_top1_rd_addr_m_5_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u76 ( .A(oc8051_ram_top1_wr_addr_m_5_), 
        .B(oc8051_ram_top1_rd_addr_m_5_), .Y(oc8051_ram_top1_n64) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_u75 ( .AN(wr_addr[4]), .B(
        oc8051_ram_top1_n68), .Y(oc8051_ram_top1_wr_addr_m_4_) );
  AND2_X0P5M_A12TS oc8051_ram_top1_u74 ( .A(rd_addr[4]), .B(
        oc8051_ram_top1_n69), .Y(oc8051_ram_top1_rd_addr_m_4_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u73 ( .A(oc8051_ram_top1_wr_addr_m_4_), 
        .B(oc8051_ram_top1_rd_addr_m_4_), .Y(oc8051_ram_top1_n65) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u72 ( .A(wr_addr[3]), .B(wr_addr[6]), .S0(
        oc8051_ram_top1_n68), .Y(oc8051_ram_top1_wr_addr_m_3_) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_u71 ( .A(rd_addr[3]), .B(rd_addr[6]), .S0(
        oc8051_ram_top1_n67), .Y(oc8051_ram_top1_rd_addr_m_3_) );
  XNOR2_X0P5M_A12TS oc8051_ram_top1_u70 ( .A(oc8051_ram_top1_wr_addr_m_3_), 
        .B(oc8051_ram_top1_rd_addr_m_3_), .Y(oc8051_ram_top1_n66) );
  AND4_X0P5M_A12TS oc8051_ram_top1_u69 ( .A(oc8051_ram_top1_n63), .B(
        oc8051_ram_top1_n64), .C(oc8051_ram_top1_n65), .D(oc8051_ram_top1_n66), 
        .Y(oc8051_ram_top1_n62) );
  NAND4B_X0P5M_A12TS oc8051_ram_top1_u68 ( .AN(oc8051_ram_top1_n59), .B(
        oc8051_ram_top1_n60), .C(oc8051_ram_top1_n61), .D(oc8051_ram_top1_n62), 
        .Y(oc8051_ram_top1_n53) );
  INV_X0P5B_A12TS oc8051_ram_top1_u67 ( .A(oc8051_ram_top1_n53), .Y(
        oc8051_ram_top1_n76) );
  INV_X0P5B_A12TS oc8051_ram_top1_u66 ( .A(oc8051_ram_top1_n58), .Y(
        ram_data[0]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u65 ( .A(oc8051_ram_top1_n57), .Y(
        ram_data[1]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u64 ( .A(oc8051_ram_top1_n56), .Y(
        ram_data[2]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u63 ( .A(oc8051_ram_top1_n55), .Y(
        ram_data[3]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u62 ( .A(oc8051_ram_top1_n54), .Y(
        ram_data[4]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u61 ( .A(oc8051_ram_top1_n52), .Y(
        ram_data[5]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u60 ( .A(oc8051_ram_top1_n51), .Y(
        ram_data[6]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u59 ( .A(oc8051_ram_top1_n50), .Y(
        ram_data[7]) );
  INV_X0P5B_A12TS oc8051_ram_top1_u58 ( .A(descy), .Y(oc8051_ram_top1_n10) );
  INV_X0P5B_A12TS oc8051_ram_top1_u57 ( .A(oc8051_ram_top1_n260), .Y(
        oc8051_ram_top1_n47) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u56 ( .A(oc8051_ram_top1_n13), .B(
        oc8051_ram_top1_n280), .Y(oc8051_ram_top1_n49) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u55 ( .A(oc8051_ram_top1_n47), .B(
        oc8051_ram_top1_n48), .C(oc8051_ram_top1_n49), .Y(oc8051_ram_top1_n28)
         );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u54 ( .A(oc8051_ram_top1_n49), .B(
        oc8051_ram_top1_n48), .C(oc8051_ram_top1_n260), .Y(oc8051_ram_top1_n26) );
  AND2_X0P5M_A12TS oc8051_ram_top1_u53 ( .A(oc8051_ram_top1_n280), .B(
        oc8051_ram_top1_bit_addr_r), .Y(oc8051_ram_top1_n46) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u52 ( .A(oc8051_ram_top1_n46), .B(
        oc8051_ram_top1_n48), .C(oc8051_ram_top1_n260), .Y(oc8051_ram_top1_n21) );
  INV_X0P5B_A12TS oc8051_ram_top1_u51 ( .A(oc8051_ram_top1_n21), .Y(
        oc8051_ram_top1_n19) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u50 ( .A(oc8051_ram_top1_n46), .B(
        oc8051_ram_top1_n47), .C(oc8051_ram_top1_n270), .Y(oc8051_ram_top1_n16) );
  INV_X0P5B_A12TS oc8051_ram_top1_u49 ( .A(oc8051_ram_top1_n16), .Y(
        oc8051_ram_top1_n24) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u48 ( .A(oc8051_ram_top1_n19), .B(
        oc8051_ram_top1_n24), .Y(oc8051_ram_top1_n14) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u47 ( .A(oc8051_ram_top1_n260), .B(
        oc8051_ram_top1_n49), .C(oc8051_ram_top1_n270), .Y(oc8051_ram_top1_n32) );
  INV_X0P5B_A12TS oc8051_ram_top1_u46 ( .A(oc8051_ram_top1_n32), .Y(
        oc8051_ram_top1_n40) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u45 ( .A(oc8051_ram_top1_n49), .B(
        oc8051_ram_top1_n47), .C(oc8051_ram_top1_n270), .Y(oc8051_ram_top1_n37) );
  INV_X0P5B_A12TS oc8051_ram_top1_u44 ( .A(oc8051_ram_top1_n37), .Y(
        oc8051_ram_top1_n35) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_u43 ( .A(oc8051_ram_top1_n40), .B(
        oc8051_ram_top1_n35), .Y(oc8051_ram_top1_n25) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u42 ( .A(oc8051_ram_top1_n47), .B(
        oc8051_ram_top1_n48), .C(oc8051_ram_top1_n46), .Y(oc8051_ram_top1_n27)
         );
  NAND3_X0P5A_A12TS oc8051_ram_top1_u41 ( .A(oc8051_ram_top1_n260), .B(
        oc8051_ram_top1_n46), .C(oc8051_ram_top1_n270), .Y(oc8051_ram_top1_n9)
         );
  NAND4_X0P5A_A12TS oc8051_ram_top1_u40 ( .A(oc8051_ram_top1_n14), .B(
        oc8051_ram_top1_n25), .C(oc8051_ram_top1_n27), .D(oc8051_ram_top1_n9), 
        .Y(oc8051_ram_top1_n43) );
  OAI2XB1_X0P5M_A12TS oc8051_ram_top1_u39 ( .A1N(oc8051_ram_top1_n26), .A0(
        oc8051_ram_top1_n43), .B0(ram_data[0]), .Y(oc8051_ram_top1_n44) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u38 ( .A(wr_dat[0]), .B(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n45) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u37 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n28), .B0(oc8051_ram_top1_n44), .C0(
        oc8051_ram_top1_n45), .Y(oc8051_ram_top1_wr_data_m[0]) );
  OAI2XB1_X0P5M_A12TS oc8051_ram_top1_u36 ( .A1N(oc8051_ram_top1_n28), .A0(
        oc8051_ram_top1_n43), .B0(ram_data[1]), .Y(oc8051_ram_top1_n41) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u35 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n26), .B0(oc8051_ram_top1_n41), .C0(
        oc8051_ram_top1_n42), .Y(oc8051_ram_top1_wr_data_m[1]) );
  AND4_X0P5M_A12TS oc8051_ram_top1_u34 ( .A(oc8051_ram_top1_n14), .B(
        oc8051_ram_top1_n26), .C(oc8051_ram_top1_n28), .D(oc8051_ram_top1_n9), 
        .Y(oc8051_ram_top1_n31) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u33 ( .A(oc8051_ram_top1_n31), .B(
        oc8051_ram_top1_n27), .Y(oc8051_ram_top1_n36) );
  OAI21_X0P5M_A12TS oc8051_ram_top1_u32 ( .A0(oc8051_ram_top1_n40), .A1(
        oc8051_ram_top1_n36), .B0(ram_data[2]), .Y(oc8051_ram_top1_n38) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u31 ( .A(wr_dat[2]), .B(
        oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n39) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u30 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n37), .B0(oc8051_ram_top1_n38), .C0(
        oc8051_ram_top1_n39), .Y(oc8051_ram_top1_wr_data_m[2]) );
  OAI21_X0P5M_A12TS oc8051_ram_top1_u29 ( .A0(oc8051_ram_top1_n35), .A1(
        oc8051_ram_top1_n36), .B0(ram_data[3]), .Y(oc8051_ram_top1_n33) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u28 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n32), .B0(oc8051_ram_top1_n33), .C0(
        oc8051_ram_top1_n34), .Y(oc8051_ram_top1_wr_data_m[3]) );
  AO1B2_X0P5M_A12TS oc8051_ram_top1_u27 ( .B0(oc8051_ram_top1_n25), .B1(
        oc8051_ram_top1_n31), .A0N(ram_data[4]), .Y(oc8051_ram_top1_n29) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u26 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n27), .B0(oc8051_ram_top1_n29), .C0(
        oc8051_ram_top1_n30), .Y(oc8051_ram_top1_wr_data_m[4]) );
  AND4_X0P5M_A12TS oc8051_ram_top1_u25 ( .A(oc8051_ram_top1_n25), .B(
        oc8051_ram_top1_n26), .C(oc8051_ram_top1_n27), .D(oc8051_ram_top1_n28), 
        .Y(oc8051_ram_top1_n15) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_u24 ( .A(oc8051_ram_top1_n15), .B(
        oc8051_ram_top1_n9), .Y(oc8051_ram_top1_n20) );
  OAI21_X0P5M_A12TS oc8051_ram_top1_u23 ( .A0(oc8051_ram_top1_n24), .A1(
        oc8051_ram_top1_n20), .B0(ram_data[5]), .Y(oc8051_ram_top1_n22) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u22 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n21), .B0(oc8051_ram_top1_n22), .C0(
        oc8051_ram_top1_n23), .Y(oc8051_ram_top1_wr_data_m[5]) );
  OAI21_X0P5M_A12TS oc8051_ram_top1_u21 ( .A0(oc8051_ram_top1_n19), .A1(
        oc8051_ram_top1_n20), .B0(ram_data[6]), .Y(oc8051_ram_top1_n17) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u20 ( .A0(oc8051_ram_top1_n10), .A1(
        oc8051_ram_top1_n16), .B0(oc8051_ram_top1_n17), .C0(
        oc8051_ram_top1_n18), .Y(oc8051_ram_top1_wr_data_m[6]) );
  AO1B2_X0P5M_A12TS oc8051_ram_top1_u19 ( .B0(oc8051_ram_top1_n14), .B1(
        oc8051_ram_top1_n15), .A0N(ram_data[7]), .Y(oc8051_ram_top1_n11) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_u18 ( .A0(oc8051_ram_top1_n9), .A1(
        oc8051_ram_top1_n10), .B0(oc8051_ram_top1_n11), .C0(
        oc8051_ram_top1_n12), .Y(oc8051_ram_top1_wr_data_m[7]) );
  TIEHI_X1M_A12TS oc8051_ram_top1_u17 ( .Y(oc8051_ram_top1__logic1_) );
  BUFH_X1M_A12TS oc8051_ram_top1_u16 ( .A(oc8051_ram_top1_wr_data_m[0]), .Y(
        oc8051_ram_top1_n1) );
  BUFH_X1M_A12TS oc8051_ram_top1_u15 ( .A(oc8051_ram_top1_wr_data_m[2]), .Y(
        oc8051_ram_top1_n3) );
  BUFH_X1M_A12TS oc8051_ram_top1_u14 ( .A(oc8051_ram_top1_wr_data_m[1]), .Y(
        oc8051_ram_top1_n2) );
  BUFH_X1M_A12TS oc8051_ram_top1_u13 ( .A(oc8051_ram_top1_wr_data_m[6]), .Y(
        oc8051_ram_top1_n7) );
  BUFH_X1M_A12TS oc8051_ram_top1_u12 ( .A(oc8051_ram_top1_wr_data_m[5]), .Y(
        oc8051_ram_top1_n6) );
  BUFH_X1M_A12TS oc8051_ram_top1_u11 ( .A(oc8051_ram_top1_wr_data_m[4]), .Y(
        oc8051_ram_top1_n5) );
  BUFH_X1M_A12TS oc8051_ram_top1_u10 ( .A(oc8051_ram_top1_wr_data_m[3]), .Y(
        oc8051_ram_top1_n4) );
  BUFH_X1M_A12TS oc8051_ram_top1_u9 ( .A(oc8051_ram_top1_wr_data_m[7]), .Y(
        oc8051_ram_top1_n8) );
  NAND2_X0P5M_A12TS oc8051_ram_top1_u8 ( .A(wr_dat[7]), .B(oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n12) );
  NAND2_X0P5M_A12TS oc8051_ram_top1_u7 ( .A(wr_dat[1]), .B(oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n42) );
  NAND2_X0P5M_A12TS oc8051_ram_top1_u6 ( .A(wr_dat[3]), .B(oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n34) );
  NAND2_X0P5M_A12TS oc8051_ram_top1_u5 ( .A(wr_dat[5]), .B(oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n23) );
  NAND2_X0P5M_A12TS oc8051_ram_top1_u4 ( .A(wr_dat[6]), .B(oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n18) );
  NAND2_X0P5M_A12TS oc8051_ram_top1_u3 ( .A(wr_dat[4]), .B(oc8051_ram_top1_n13), .Y(oc8051_ram_top1_n30) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_rd_en_r_reg ( .D(oc8051_ram_top1_n76), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_rd_en_r) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_select_reg_0_ ( .D(rd_addr[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_n260) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_select_reg_1_ ( .D(rd_addr[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_n270) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_select_reg_2_ ( .D(rd_addr[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_n280) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_bit_addr_r_reg ( .D(bit_addr_o), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_bit_addr_r) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_7_ ( .D(oc8051_ram_top1_n8), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_6_ ( .D(oc8051_ram_top1_n7), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_5_ ( .D(oc8051_ram_top1_n6), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_4_ ( .D(oc8051_ram_top1_n5), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_3_ ( .D(oc8051_ram_top1_n4), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_2_ ( .D(oc8051_ram_top1_n3), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_1_ ( .D(oc8051_ram_top1_n2), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_wr_data_r_reg_0_ ( .D(oc8051_ram_top1_n1), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_ram_top1_wr_data_r[0]) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4143 ( .A(
        oc8051_ram_top1_rd_addr_m_6_), .Y(oc8051_ram_top1_oc8051_idata_n2465)
         );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4142 ( .A(
        oc8051_ram_top1_oc8051_idata_n2465), .B(oc8051_ram_top1_wr_addr_m_6_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4644) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4141 ( .A(
        oc8051_ram_top1_rd_addr_m_5_), .Y(oc8051_ram_top1_oc8051_idata_n4639)
         );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4140 ( .A(
        oc8051_ram_top1_oc8051_idata_n4639), .B(oc8051_ram_top1_wr_addr_m_5_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4645) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4139 ( .A(
        oc8051_ram_top1_wr_addr_m_3_), .B(oc8051_ram_top1_rd_addr_m_3_), .Y(
        oc8051_ram_top1_oc8051_idata_n4652) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4138 ( .A(
        oc8051_ram_top1_wr_addr_m_4_), .B(oc8051_ram_top1_rd_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_n4653) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4137 ( .A(wr_addr[7]), .B(
        rd_addr[7]), .Y(oc8051_ram_top1_oc8051_idata_n4654) );
  NOR3_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4136 ( .A(
        oc8051_ram_top1_oc8051_idata_n4652), .B(
        oc8051_ram_top1_oc8051_idata_n4653), .C(
        oc8051_ram_top1_oc8051_idata_n4654), .Y(
        oc8051_ram_top1_oc8051_idata_n4646) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4135 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .Y(oc8051_ram_top1_oc8051_idata_n4643)
         );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4134 ( .A(
        oc8051_ram_top1_oc8051_idata_n4643), .B(oc8051_ram_top1_wr_addr_m_0_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4651) );
  NAND3_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4133 ( .A(
        oc8051_ram_top1_n53), .B(n_0_net_), .C(
        oc8051_ram_top1_oc8051_idata_n4651), .Y(
        oc8051_ram_top1_oc8051_idata_n4648) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4132 ( .A(
        oc8051_ram_top1_wr_addr_m_1_), .B(oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_n4649) );
  XOR2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4131 ( .A(
        oc8051_ram_top1_wr_addr_m_2_), .B(oc8051_ram_top1_rd_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_n4650) );
  NOR3_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4130 ( .A(
        oc8051_ram_top1_oc8051_idata_n4648), .B(
        oc8051_ram_top1_oc8051_idata_n4649), .C(
        oc8051_ram_top1_oc8051_idata_n4650), .Y(
        oc8051_ram_top1_oc8051_idata_n4647) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4129 ( .A(
        oc8051_ram_top1_oc8051_idata_n4644), .B(
        oc8051_ram_top1_oc8051_idata_n4645), .C(
        oc8051_ram_top1_oc8051_idata_n4646), .D(
        oc8051_ram_top1_oc8051_idata_n4647), .Y(
        oc8051_ram_top1_oc8051_idata_n1087) );
  NAND2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4128 ( .A(
        oc8051_ram_top1_n53), .B(oc8051_ram_top1_oc8051_idata_n1087), .Y(
        oc8051_ram_top1_oc8051_idata_n2466) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4127 ( .AN(rd_addr[7]), .B(
        oc8051_ram_top1_oc8051_idata_n2466), .Y(
        oc8051_ram_top1_oc8051_idata_n4565) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4126 ( .AN(
        oc8051_ram_top1_oc8051_idata_n4565), .B(
        oc8051_ram_top1_oc8051_idata_n2465), .Y(
        oc8051_ram_top1_oc8051_idata_n1286) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4125 ( .A(
        oc8051_ram_top1_oc8051_idata_n4639), .B(oc8051_ram_top1_rd_addr_m_4_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4616) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4124 ( .A(
        oc8051_ram_top1_rd_addr_m_3_), .Y(oc8051_ram_top1_oc8051_idata_n4640)
         );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4123 ( .A(
        oc8051_ram_top1_oc8051_idata_n4640), .B(oc8051_ram_top1_rd_addr_m_2_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4586) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4122 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4586), .Y(
        oc8051_ram_top1_oc8051_idata_n4641) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4121 ( .A(
        oc8051_ram_top1_rd_addr_m_0_), .B(oc8051_ram_top1_rd_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_n4587) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4120 ( .A(
        oc8051_ram_top1_oc8051_idata_n4641), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1200) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4119 ( .A(
        oc8051_ram_top1_oc8051_idata_n4643), .B(oc8051_ram_top1_rd_addr_m_1_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4589) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4118 ( .A(
        oc8051_ram_top1_oc8051_idata_n4641), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1201) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4117 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4635) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4116 ( .A(
        oc8051_ram_top1_rd_addr_m_1_), .Y(oc8051_ram_top1_oc8051_idata_n4642)
         );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4115 ( .A(
        oc8051_ram_top1_oc8051_idata_n4642), .B(oc8051_ram_top1_rd_addr_m_0_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4590) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4114 ( .A(
        oc8051_ram_top1_oc8051_idata_n4641), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1198) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4113 ( .A(
        oc8051_ram_top1_oc8051_idata_n4642), .B(
        oc8051_ram_top1_oc8051_idata_n4643), .Y(
        oc8051_ram_top1_oc8051_idata_n4591) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4112 ( .A(
        oc8051_ram_top1_oc8051_idata_n4641), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1199) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4111 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4636) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4110 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .Y(oc8051_ram_top1_oc8051_idata_n4628)
         );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4109 ( .A(
        oc8051_ram_top1_oc8051_idata_n4640), .B(
        oc8051_ram_top1_oc8051_idata_n4628), .Y(
        oc8051_ram_top1_oc8051_idata_n4634) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4108 ( .A(
        oc8051_ram_top1_oc8051_idata_n4634), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n4594) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4107 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4594), .Y(
        oc8051_ram_top1_oc8051_idata_n1196) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4106 ( .A(
        oc8051_ram_top1_rd_addr_m_4_), .Y(oc8051_ram_top1_oc8051_idata_n4609)
         );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4105 ( .A(
        oc8051_ram_top1_oc8051_idata_n4639), .B(
        oc8051_ram_top1_oc8051_idata_n4609), .Y(
        oc8051_ram_top1_oc8051_idata_n4623) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4104 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4586), .Y(
        oc8051_ram_top1_oc8051_idata_n4633) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4103 ( .A(
        oc8051_ram_top1_oc8051_idata_n4633), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1197) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4102 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4637) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4101 ( .A(
        oc8051_ram_top1_oc8051_idata_n4634), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n4593) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4100 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4593), .Y(
        oc8051_ram_top1_oc8051_idata_n1194) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4099 ( .A(
        oc8051_ram_top1_oc8051_idata_n4633), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1195) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4098 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4638) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4097 ( .A(
        oc8051_ram_top1_oc8051_idata_n4635), .B(
        oc8051_ram_top1_oc8051_idata_n4636), .C(
        oc8051_ram_top1_oc8051_idata_n4637), .D(
        oc8051_ram_top1_oc8051_idata_n4638), .Y(
        oc8051_ram_top1_oc8051_idata_n4567) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4096 ( .A(
        oc8051_ram_top1_oc8051_idata_n4634), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n4596) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4095 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4596), .Y(
        oc8051_ram_top1_oc8051_idata_n1188) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4094 ( .A(
        oc8051_ram_top1_oc8051_idata_n4633), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1189) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4093 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4629) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4092 ( .A(
        oc8051_ram_top1_oc8051_idata_n4634), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n4595) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4091 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4595), .Y(
        oc8051_ram_top1_oc8051_idata_n1186) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4090 ( .A(
        oc8051_ram_top1_oc8051_idata_n4633), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1187) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4089 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4630) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4088 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4594), .Y(
        oc8051_ram_top1_oc8051_idata_n1184) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4087 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4593), .Y(
        oc8051_ram_top1_oc8051_idata_n1185) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4086 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4631) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4085 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4596), .Y(
        oc8051_ram_top1_oc8051_idata_n1182) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4084 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4595), .Y(
        oc8051_ram_top1_oc8051_idata_n1183) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4083 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4632) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4082 ( .A(
        oc8051_ram_top1_oc8051_idata_n4629), .B(
        oc8051_ram_top1_oc8051_idata_n4630), .C(
        oc8051_ram_top1_oc8051_idata_n4631), .D(
        oc8051_ram_top1_oc8051_idata_n4632), .Y(
        oc8051_ram_top1_oc8051_idata_n4568) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4081 ( .A(
        oc8051_ram_top1_oc8051_idata_n4628), .B(oc8051_ram_top1_rd_addr_m_3_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4584) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4080 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4584), .Y(
        oc8051_ram_top1_oc8051_idata_n4627) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4079 ( .A(
        oc8051_ram_top1_oc8051_idata_n4627), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1171) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4078 ( .A(
        oc8051_ram_top1_oc8051_idata_n507), .Y(
        oc8051_ram_top1_oc8051_idata_n4624) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4077 ( .A(
        oc8051_ram_top1_oc8051_idata_n4627), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1173) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4076 ( .A(
        oc8051_ram_top1_oc8051_idata_n515), .Y(
        oc8051_ram_top1_oc8051_idata_n4625) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4075 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n1062) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4074 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n1072) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4073 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1062), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1072), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n4626) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4072 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n4624), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n4625), .C0(
        oc8051_ram_top1_oc8051_idata_n4626), .Y(
        oc8051_ram_top1_oc8051_idata_n4610) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4071 ( .A(
        oc8051_ram_top1_rd_addr_m_2_), .B(oc8051_ram_top1_rd_addr_m_3_), .Y(
        oc8051_ram_top1_oc8051_idata_n4578) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4070 ( .A(
        oc8051_ram_top1_oc8051_idata_n4623), .B(
        oc8051_ram_top1_oc8051_idata_n4578), .Y(
        oc8051_ram_top1_oc8051_idata_n4622) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4069 ( .A(
        oc8051_ram_top1_oc8051_idata_n4622), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1164) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4068 ( .A(
        oc8051_ram_top1_oc8051_idata_n491), .Y(
        oc8051_ram_top1_oc8051_idata_n4619) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4067 ( .A(
        oc8051_ram_top1_oc8051_idata_n4622), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1166) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4066 ( .A(
        oc8051_ram_top1_oc8051_idata_n499), .Y(
        oc8051_ram_top1_oc8051_idata_n4620) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4065 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n1036) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u4064 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n1048) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4063 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1036), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1048), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n4621) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4062 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n4619), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n4620), .C0(
        oc8051_ram_top1_oc8051_idata_n4621), .Y(
        oc8051_ram_top1_oc8051_idata_n4611) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4061 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4584), .Y(
        oc8051_ram_top1_oc8051_idata_n4618) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4060 ( .A(
        oc8051_ram_top1_oc8051_idata_n4618), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1159) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4059 ( .A(
        oc8051_ram_top1_oc8051_idata_n4618), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1160) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4058 ( .A0(
        oc8051_ram_top1_oc8051_idata_n483), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n475), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n4617) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4057 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4617), .Y(
        oc8051_ram_top1_oc8051_idata_n4612) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4056 ( .A(
        oc8051_ram_top1_oc8051_idata_n4616), .B(
        oc8051_ram_top1_oc8051_idata_n4578), .Y(
        oc8051_ram_top1_oc8051_idata_n4615) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4055 ( .A(
        oc8051_ram_top1_oc8051_idata_n4615), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1154) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4054 ( .A(
        oc8051_ram_top1_oc8051_idata_n4615), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1155) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4053 ( .A0(
        oc8051_ram_top1_oc8051_idata_n467), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n459), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n4614) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4052 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4614), .Y(
        oc8051_ram_top1_oc8051_idata_n4613) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4051 ( .A(
        oc8051_ram_top1_oc8051_idata_n4610), .B(
        oc8051_ram_top1_oc8051_idata_n4611), .C(
        oc8051_ram_top1_oc8051_idata_n4612), .D(
        oc8051_ram_top1_oc8051_idata_n4613), .Y(
        oc8051_ram_top1_oc8051_idata_n4569) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4050 ( .A(
        oc8051_ram_top1_oc8051_idata_n4609), .B(oc8051_ram_top1_rd_addr_m_5_), 
        .Y(oc8051_ram_top1_oc8051_idata_n4602) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4049 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4594), .Y(
        oc8051_ram_top1_oc8051_idata_n1148) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4048 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4593), .Y(
        oc8051_ram_top1_oc8051_idata_n1149) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4047 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4604) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4046 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4596), .Y(
        oc8051_ram_top1_oc8051_idata_n1146) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4045 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4595), .Y(
        oc8051_ram_top1_oc8051_idata_n1147) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4044 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4605) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4043 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4586), .Y(
        oc8051_ram_top1_oc8051_idata_n4608) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4042 ( .A(
        oc8051_ram_top1_oc8051_idata_n4608), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1144) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4041 ( .A(
        oc8051_ram_top1_oc8051_idata_n4608), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1145) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4040 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4606) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4039 ( .A(
        oc8051_ram_top1_oc8051_idata_n4608), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1142) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4038 ( .A(
        oc8051_ram_top1_oc8051_idata_n4608), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1143) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4037 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4607) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4036 ( .A(
        oc8051_ram_top1_oc8051_idata_n4604), .B(
        oc8051_ram_top1_oc8051_idata_n4605), .C(
        oc8051_ram_top1_oc8051_idata_n4606), .D(
        oc8051_ram_top1_oc8051_idata_n4607), .Y(
        oc8051_ram_top1_oc8051_idata_n4570) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4035 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4584), .Y(
        oc8051_ram_top1_oc8051_idata_n4603) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4034 ( .A(
        oc8051_ram_top1_oc8051_idata_n4603), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1136) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4033 ( .A(
        oc8051_ram_top1_oc8051_idata_n4603), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1137) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4032 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4597) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4031 ( .A(
        oc8051_ram_top1_oc8051_idata_n4603), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1134) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4030 ( .A(
        oc8051_ram_top1_oc8051_idata_n4603), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1135) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4029 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4598) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4028 ( .A(
        oc8051_ram_top1_oc8051_idata_n4602), .B(
        oc8051_ram_top1_oc8051_idata_n4578), .Y(
        oc8051_ram_top1_oc8051_idata_n4601) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4027 ( .A(
        oc8051_ram_top1_oc8051_idata_n4601), .B(
        oc8051_ram_top1_oc8051_idata_n4591), .Y(
        oc8051_ram_top1_oc8051_idata_n1132) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4026 ( .A(
        oc8051_ram_top1_oc8051_idata_n4601), .B(
        oc8051_ram_top1_oc8051_idata_n4590), .Y(
        oc8051_ram_top1_oc8051_idata_n1133) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4025 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4599) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4024 ( .A(
        oc8051_ram_top1_oc8051_idata_n4601), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1130) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4023 ( .A(
        oc8051_ram_top1_oc8051_idata_n4601), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1131) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4022 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4600) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4021 ( .A(
        oc8051_ram_top1_oc8051_idata_n4597), .B(
        oc8051_ram_top1_oc8051_idata_n4598), .C(
        oc8051_ram_top1_oc8051_idata_n4599), .D(
        oc8051_ram_top1_oc8051_idata_n4600), .Y(
        oc8051_ram_top1_oc8051_idata_n4571) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u4020 ( .A(
        oc8051_ram_top1_rd_addr_m_4_), .B(oc8051_ram_top1_rd_addr_m_5_), .Y(
        oc8051_ram_top1_oc8051_idata_n4588) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4019 ( .A(
        oc8051_ram_top1_oc8051_idata_n4596), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n1121) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4018 ( .A(
        oc8051_ram_top1_oc8051_idata_n4595), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n1122) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4017 ( .A0(
        oc8051_ram_top1_oc8051_idata_n451), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n443), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n4592) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4016 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4592), .Y(
        oc8051_ram_top1_oc8051_idata_n4573) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4015 ( .A(
        oc8051_ram_top1_oc8051_idata_n4591), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n4582) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4014 ( .A(
        oc8051_ram_top1_oc8051_idata_n4586), .B(
        oc8051_ram_top1_oc8051_idata_n4582), .Y(
        oc8051_ram_top1_oc8051_idata_n1116) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4013 ( .A(
        oc8051_ram_top1_oc8051_idata_n4590), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n4581) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4012 ( .A(
        oc8051_ram_top1_oc8051_idata_n4586), .B(
        oc8051_ram_top1_oc8051_idata_n4581), .Y(
        oc8051_ram_top1_oc8051_idata_n1117) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4011 ( .A(
        oc8051_ram_top1_oc8051_idata_n4589), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n4580) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4010 ( .A(
        oc8051_ram_top1_oc8051_idata_n4587), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n4579) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4009 ( .A0(
        oc8051_ram_top1_oc8051_idata_n435), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n427), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n4585) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4008 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4585), .Y(
        oc8051_ram_top1_oc8051_idata_n4574) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4007 ( .A(
        oc8051_ram_top1_oc8051_idata_n4584), .B(
        oc8051_ram_top1_oc8051_idata_n4582), .Y(
        oc8051_ram_top1_oc8051_idata_n1111) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4006 ( .A(
        oc8051_ram_top1_oc8051_idata_n4584), .B(
        oc8051_ram_top1_oc8051_idata_n4581), .Y(
        oc8051_ram_top1_oc8051_idata_n1112) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4005 ( .A0(
        oc8051_ram_top1_oc8051_idata_n419), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n411), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n4583) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4004 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4583), .Y(
        oc8051_ram_top1_oc8051_idata_n4575) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4003 ( .A(
        oc8051_ram_top1_oc8051_idata_n4582), .B(
        oc8051_ram_top1_oc8051_idata_n4578), .Y(
        oc8051_ram_top1_oc8051_idata_n1106) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4002 ( .A(
        oc8051_ram_top1_oc8051_idata_n4581), .B(
        oc8051_ram_top1_oc8051_idata_n4578), .Y(
        oc8051_ram_top1_oc8051_idata_n1107) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4001 ( .A0(
        oc8051_ram_top1_oc8051_idata_n403), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n395), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n4577) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u4000 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4577), .Y(
        oc8051_ram_top1_oc8051_idata_n4576) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3999 ( .A(
        oc8051_ram_top1_oc8051_idata_n4573), .B(
        oc8051_ram_top1_oc8051_idata_n4574), .C(
        oc8051_ram_top1_oc8051_idata_n4575), .D(
        oc8051_ram_top1_oc8051_idata_n4576), .Y(
        oc8051_ram_top1_oc8051_idata_n4572) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3998 ( .A(
        oc8051_ram_top1_oc8051_idata_n4567), .B(
        oc8051_ram_top1_oc8051_idata_n4568), .C(
        oc8051_ram_top1_oc8051_idata_n4569), .D(
        oc8051_ram_top1_oc8051_idata_n4570), .E(
        oc8051_ram_top1_oc8051_idata_n4571), .F(
        oc8051_ram_top1_oc8051_idata_n4572), .Y(
        oc8051_ram_top1_oc8051_idata_n4566) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3997 ( .A(
        oc8051_ram_top1_oc8051_idata_n2466), .B(
        oc8051_ram_top1_oc8051_idata_n1087), .Y(
        oc8051_ram_top1_oc8051_idata_n1288) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3996 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n4566), .B0(oc8051_ram_top1_rd_data_m[0]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n2375) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3995 ( .AN(
        oc8051_ram_top1_oc8051_idata_n4565), .B(oc8051_ram_top1_rd_addr_m_6_), 
        .Y(oc8051_ram_top1_oc8051_idata_n1090) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3994 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4561) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3993 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4562) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3992 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4563) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3991 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4564) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3990 ( .A(
        oc8051_ram_top1_oc8051_idata_n4561), .B(
        oc8051_ram_top1_oc8051_idata_n4562), .C(
        oc8051_ram_top1_oc8051_idata_n4563), .D(
        oc8051_ram_top1_oc8051_idata_n4564), .Y(
        oc8051_ram_top1_oc8051_idata_n2467) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3989 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4557) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3988 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4558) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3987 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4559) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3986 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4560) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3985 ( .A(
        oc8051_ram_top1_oc8051_idata_n4557), .B(
        oc8051_ram_top1_oc8051_idata_n4558), .C(
        oc8051_ram_top1_oc8051_idata_n4559), .D(
        oc8051_ram_top1_oc8051_idata_n4560), .Y(
        oc8051_ram_top1_oc8051_idata_n2468) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3984 ( .A(
        oc8051_ram_top1_oc8051_idata_n379), .Y(
        oc8051_ram_top1_oc8051_idata_n4554) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3983 ( .A(
        oc8051_ram_top1_oc8051_idata_n387), .Y(
        oc8051_ram_top1_oc8051_idata_n4555) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3982 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n954) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3981 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n963) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3980 ( .A0(
        oc8051_ram_top1_oc8051_idata_n954), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n963), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n4556) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3979 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n4554), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n4555), .C0(
        oc8051_ram_top1_oc8051_idata_n4556), .Y(
        oc8051_ram_top1_oc8051_idata_n4545) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3978 ( .A(
        oc8051_ram_top1_oc8051_idata_n363), .Y(
        oc8051_ram_top1_oc8051_idata_n4551) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3977 ( .A(
        oc8051_ram_top1_oc8051_idata_n371), .Y(
        oc8051_ram_top1_oc8051_idata_n4552) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3976 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n933) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3975 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n943) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3974 ( .A0(
        oc8051_ram_top1_oc8051_idata_n933), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n943), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n4553) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3973 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n4551), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n4552), .C0(
        oc8051_ram_top1_oc8051_idata_n4553), .Y(
        oc8051_ram_top1_oc8051_idata_n4546) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3972 ( .A0(
        oc8051_ram_top1_oc8051_idata_n355), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n347), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n4550) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3971 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4550), .Y(
        oc8051_ram_top1_oc8051_idata_n4547) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3970 ( .A0(
        oc8051_ram_top1_oc8051_idata_n339), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n331), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n4549) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3969 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4549), .Y(
        oc8051_ram_top1_oc8051_idata_n4548) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3968 ( .A(
        oc8051_ram_top1_oc8051_idata_n4545), .B(
        oc8051_ram_top1_oc8051_idata_n4546), .C(
        oc8051_ram_top1_oc8051_idata_n4547), .D(
        oc8051_ram_top1_oc8051_idata_n4548), .Y(
        oc8051_ram_top1_oc8051_idata_n2469) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3967 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4541) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3966 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4542) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3965 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4543) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3964 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4544) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3963 ( .A(
        oc8051_ram_top1_oc8051_idata_n4541), .B(
        oc8051_ram_top1_oc8051_idata_n4542), .C(
        oc8051_ram_top1_oc8051_idata_n4543), .D(
        oc8051_ram_top1_oc8051_idata_n4544), .Y(
        oc8051_ram_top1_oc8051_idata_n2470) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3962 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4537) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3961 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4538) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3960 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4539) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3959 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n4540) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3958 ( .A(
        oc8051_ram_top1_oc8051_idata_n4537), .B(
        oc8051_ram_top1_oc8051_idata_n4538), .C(
        oc8051_ram_top1_oc8051_idata_n4539), .D(
        oc8051_ram_top1_oc8051_idata_n4540), .Y(
        oc8051_ram_top1_oc8051_idata_n2471) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3957 ( .A0(
        oc8051_ram_top1_oc8051_idata_n323), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n315), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n4536) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3956 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4536), .Y(
        oc8051_ram_top1_oc8051_idata_n2473) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3955 ( .A0(
        oc8051_ram_top1_oc8051_idata_n307), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n299), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n4535) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3954 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4535), .Y(
        oc8051_ram_top1_oc8051_idata_n2474) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3953 ( .A0(
        oc8051_ram_top1_oc8051_idata_n291), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n283), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n4534) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3952 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4534), .Y(
        oc8051_ram_top1_oc8051_idata_n4531) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3951 ( .A0(
        oc8051_ram_top1_oc8051_idata_n275), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n267), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n4533) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3950 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n4533), .Y(
        oc8051_ram_top1_oc8051_idata_n4532) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3949 ( .A(
        oc8051_ram_top1_oc8051_idata_n2473), .B(
        oc8051_ram_top1_oc8051_idata_n2474), .C(
        oc8051_ram_top1_oc8051_idata_n4531), .D(
        oc8051_ram_top1_oc8051_idata_n4532), .Y(
        oc8051_ram_top1_oc8051_idata_n2472) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3948 ( .A(
        oc8051_ram_top1_oc8051_idata_n2467), .B(
        oc8051_ram_top1_oc8051_idata_n2468), .C(
        oc8051_ram_top1_oc8051_idata_n2469), .D(
        oc8051_ram_top1_oc8051_idata_n2470), .E(
        oc8051_ram_top1_oc8051_idata_n2471), .F(
        oc8051_ram_top1_oc8051_idata_n2472), .Y(
        oc8051_ram_top1_oc8051_idata_n2377) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3947 ( .A(
        oc8051_ram_top1_oc8051_idata_n2466), .B(rd_addr[7]), .Y(
        oc8051_ram_top1_oc8051_idata_n2422) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3946 ( .AN(
        oc8051_ram_top1_oc8051_idata_n2422), .B(
        oc8051_ram_top1_oc8051_idata_n2465), .Y(
        oc8051_ram_top1_oc8051_idata_n1092) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3945 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2461) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3944 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2462) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3943 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2463) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3942 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2464) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3941 ( .A(
        oc8051_ram_top1_oc8051_idata_n2461), .B(
        oc8051_ram_top1_oc8051_idata_n2462), .C(
        oc8051_ram_top1_oc8051_idata_n2463), .D(
        oc8051_ram_top1_oc8051_idata_n2464), .Y(
        oc8051_ram_top1_oc8051_idata_n2423) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3940 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2457) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3939 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2458) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3938 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2459) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3937 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2460) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3936 ( .A(
        oc8051_ram_top1_oc8051_idata_n2457), .B(
        oc8051_ram_top1_oc8051_idata_n2458), .C(
        oc8051_ram_top1_oc8051_idata_n2459), .D(
        oc8051_ram_top1_oc8051_idata_n2460), .Y(
        oc8051_ram_top1_oc8051_idata_n2424) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3935 ( .A(
        oc8051_ram_top1_oc8051_idata_n251), .Y(
        oc8051_ram_top1_oc8051_idata_n2454) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3934 ( .A(
        oc8051_ram_top1_oc8051_idata_n259), .Y(
        oc8051_ram_top1_oc8051_idata_n2455) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3933 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n852) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3932 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n861) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3931 ( .A0(
        oc8051_ram_top1_oc8051_idata_n852), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n861), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2456) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3930 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2454), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2455), .C0(
        oc8051_ram_top1_oc8051_idata_n2456), .Y(
        oc8051_ram_top1_oc8051_idata_n2445) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3929 ( .A(
        oc8051_ram_top1_oc8051_idata_n235), .Y(
        oc8051_ram_top1_oc8051_idata_n2451) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3928 ( .A(
        oc8051_ram_top1_oc8051_idata_n243), .Y(
        oc8051_ram_top1_oc8051_idata_n2452) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3927 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n831) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3926 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n841) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3925 ( .A0(
        oc8051_ram_top1_oc8051_idata_n831), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n841), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2453) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3924 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2451), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2452), .C0(
        oc8051_ram_top1_oc8051_idata_n2453), .Y(
        oc8051_ram_top1_oc8051_idata_n2446) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3923 ( .A0(
        oc8051_ram_top1_oc8051_idata_n227), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n219), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2450) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3922 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2450), .Y(
        oc8051_ram_top1_oc8051_idata_n2447) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3921 ( .A0(
        oc8051_ram_top1_oc8051_idata_n211), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n203), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2449) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3920 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2449), .Y(
        oc8051_ram_top1_oc8051_idata_n2448) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3919 ( .A(
        oc8051_ram_top1_oc8051_idata_n2445), .B(
        oc8051_ram_top1_oc8051_idata_n2446), .C(
        oc8051_ram_top1_oc8051_idata_n2447), .D(
        oc8051_ram_top1_oc8051_idata_n2448), .Y(
        oc8051_ram_top1_oc8051_idata_n2425) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3918 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2441) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3917 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2442) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3916 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2443) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3915 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2444) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3914 ( .A(
        oc8051_ram_top1_oc8051_idata_n2441), .B(
        oc8051_ram_top1_oc8051_idata_n2442), .C(
        oc8051_ram_top1_oc8051_idata_n2443), .D(
        oc8051_ram_top1_oc8051_idata_n2444), .Y(
        oc8051_ram_top1_oc8051_idata_n2426) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3913 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2437) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3912 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2438) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3911 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2439) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3910 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2440) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3909 ( .A(
        oc8051_ram_top1_oc8051_idata_n2437), .B(
        oc8051_ram_top1_oc8051_idata_n2438), .C(
        oc8051_ram_top1_oc8051_idata_n2439), .D(
        oc8051_ram_top1_oc8051_idata_n2440), .Y(
        oc8051_ram_top1_oc8051_idata_n2427) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3908 ( .A0(
        oc8051_ram_top1_oc8051_idata_n195), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n187), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2436) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3907 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2436), .Y(
        oc8051_ram_top1_oc8051_idata_n2429) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3906 ( .A0(
        oc8051_ram_top1_oc8051_idata_n179), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n171), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2435) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3905 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2435), .Y(
        oc8051_ram_top1_oc8051_idata_n2430) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3904 ( .A0(
        oc8051_ram_top1_oc8051_idata_n163), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n155), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2434) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3903 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2434), .Y(
        oc8051_ram_top1_oc8051_idata_n2431) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3902 ( .A0(
        oc8051_ram_top1_oc8051_idata_n147), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n139), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2433) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3901 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2433), .Y(
        oc8051_ram_top1_oc8051_idata_n2432) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3900 ( .A(
        oc8051_ram_top1_oc8051_idata_n2429), .B(
        oc8051_ram_top1_oc8051_idata_n2430), .C(
        oc8051_ram_top1_oc8051_idata_n2431), .D(
        oc8051_ram_top1_oc8051_idata_n2432), .Y(
        oc8051_ram_top1_oc8051_idata_n2428) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3899 ( .A(
        oc8051_ram_top1_oc8051_idata_n2423), .B(
        oc8051_ram_top1_oc8051_idata_n2424), .C(
        oc8051_ram_top1_oc8051_idata_n2425), .D(
        oc8051_ram_top1_oc8051_idata_n2426), .E(
        oc8051_ram_top1_oc8051_idata_n2427), .F(
        oc8051_ram_top1_oc8051_idata_n2428), .Y(
        oc8051_ram_top1_oc8051_idata_n2378) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3898 ( .AN(
        oc8051_ram_top1_oc8051_idata_n2422), .B(oc8051_ram_top1_rd_addr_m_6_), 
        .Y(oc8051_ram_top1_oc8051_idata_n1094) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3897 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2418) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3896 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2419) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3895 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2420) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3894 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2421) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3893 ( .A(
        oc8051_ram_top1_oc8051_idata_n2418), .B(
        oc8051_ram_top1_oc8051_idata_n2419), .C(
        oc8051_ram_top1_oc8051_idata_n2420), .D(
        oc8051_ram_top1_oc8051_idata_n2421), .Y(
        oc8051_ram_top1_oc8051_idata_n2380) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3892 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2414) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3891 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2415) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3890 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2416) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3889 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2417) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3888 ( .A(
        oc8051_ram_top1_oc8051_idata_n2414), .B(
        oc8051_ram_top1_oc8051_idata_n2415), .C(
        oc8051_ram_top1_oc8051_idata_n2416), .D(
        oc8051_ram_top1_oc8051_idata_n2417), .Y(
        oc8051_ram_top1_oc8051_idata_n2381) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3887 ( .A(
        oc8051_ram_top1_oc8051_idata_n123), .Y(
        oc8051_ram_top1_oc8051_idata_n2411) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3886 ( .A(
        oc8051_ram_top1_oc8051_idata_n131), .Y(
        oc8051_ram_top1_oc8051_idata_n2412) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3885 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n749) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3884 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n758) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3883 ( .A0(
        oc8051_ram_top1_oc8051_idata_n749), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n758), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2413) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3882 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2411), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2412), .C0(
        oc8051_ram_top1_oc8051_idata_n2413), .Y(
        oc8051_ram_top1_oc8051_idata_n2402) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3881 ( .A(
        oc8051_ram_top1_oc8051_idata_n107), .Y(
        oc8051_ram_top1_oc8051_idata_n2408) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3880 ( .A(
        oc8051_ram_top1_oc8051_idata_n115), .Y(
        oc8051_ram_top1_oc8051_idata_n2409) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3879 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n728) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3878 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n738) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3877 ( .A0(
        oc8051_ram_top1_oc8051_idata_n728), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n738), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2410) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3876 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2408), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2409), .C0(
        oc8051_ram_top1_oc8051_idata_n2410), .Y(
        oc8051_ram_top1_oc8051_idata_n2403) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3875 ( .A0(
        oc8051_ram_top1_oc8051_idata_n99), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n91), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2407) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3874 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2407), .Y(
        oc8051_ram_top1_oc8051_idata_n2404) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3873 ( .A0(
        oc8051_ram_top1_oc8051_idata_n83), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n75), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2406) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3872 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2406), .Y(
        oc8051_ram_top1_oc8051_idata_n2405) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3871 ( .A(
        oc8051_ram_top1_oc8051_idata_n2402), .B(
        oc8051_ram_top1_oc8051_idata_n2403), .C(
        oc8051_ram_top1_oc8051_idata_n2404), .D(
        oc8051_ram_top1_oc8051_idata_n2405), .Y(
        oc8051_ram_top1_oc8051_idata_n2382) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3870 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2398) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3869 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2399) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3868 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2400) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3867 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2401) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3866 ( .A(
        oc8051_ram_top1_oc8051_idata_n2398), .B(
        oc8051_ram_top1_oc8051_idata_n2399), .C(
        oc8051_ram_top1_oc8051_idata_n2400), .D(
        oc8051_ram_top1_oc8051_idata_n2401), .Y(
        oc8051_ram_top1_oc8051_idata_n2383) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3865 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2394) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3864 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2395) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3863 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2396) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3862 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__0_), .Y(
        oc8051_ram_top1_oc8051_idata_n2397) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3861 ( .A(
        oc8051_ram_top1_oc8051_idata_n2394), .B(
        oc8051_ram_top1_oc8051_idata_n2395), .C(
        oc8051_ram_top1_oc8051_idata_n2396), .D(
        oc8051_ram_top1_oc8051_idata_n2397), .Y(
        oc8051_ram_top1_oc8051_idata_n2384) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3860 ( .A0(
        oc8051_ram_top1_oc8051_idata_n67), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n59), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2393) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3859 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2393), .Y(
        oc8051_ram_top1_oc8051_idata_n2386) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3858 ( .A0(
        oc8051_ram_top1_oc8051_idata_n51), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n43), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2392) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3857 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2392), .Y(
        oc8051_ram_top1_oc8051_idata_n2387) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3856 ( .A0(
        oc8051_ram_top1_oc8051_idata_n35), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n27), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2391) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3855 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2391), .Y(
        oc8051_ram_top1_oc8051_idata_n2388) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3854 ( .A0(
        oc8051_ram_top1_oc8051_idata_n19), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n11), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2390) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3853 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__0_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__0_), .C0(
        oc8051_ram_top1_oc8051_idata_n2390), .Y(
        oc8051_ram_top1_oc8051_idata_n2389) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3852 ( .A(
        oc8051_ram_top1_oc8051_idata_n2386), .B(
        oc8051_ram_top1_oc8051_idata_n2387), .C(
        oc8051_ram_top1_oc8051_idata_n2388), .D(
        oc8051_ram_top1_oc8051_idata_n2389), .Y(
        oc8051_ram_top1_oc8051_idata_n2385) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3851 ( .A(
        oc8051_ram_top1_oc8051_idata_n2380), .B(
        oc8051_ram_top1_oc8051_idata_n2381), .C(
        oc8051_ram_top1_oc8051_idata_n2382), .D(
        oc8051_ram_top1_oc8051_idata_n2383), .E(
        oc8051_ram_top1_oc8051_idata_n2384), .F(
        oc8051_ram_top1_oc8051_idata_n2385), .Y(
        oc8051_ram_top1_oc8051_idata_n2379) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3850 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n2377), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n2378), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n2379), .Y(
        oc8051_ram_top1_oc8051_idata_n2376) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3849 ( .A0(
        oc8051_ram_top1_oc8051_idata_n528), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n2375), .C0(
        oc8051_ram_top1_oc8051_idata_n2376), .Y(
        oc8051_ram_top1_oc8051_idata_n2475) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3848 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2371) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3847 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2372) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3846 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2373) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3845 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2374) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3844 ( .A(
        oc8051_ram_top1_oc8051_idata_n2371), .B(
        oc8051_ram_top1_oc8051_idata_n2372), .C(
        oc8051_ram_top1_oc8051_idata_n2373), .D(
        oc8051_ram_top1_oc8051_idata_n2374), .Y(
        oc8051_ram_top1_oc8051_idata_n2333) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3843 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2367) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3842 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2368) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3841 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2369) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3840 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2370) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3839 ( .A(
        oc8051_ram_top1_oc8051_idata_n2367), .B(
        oc8051_ram_top1_oc8051_idata_n2368), .C(
        oc8051_ram_top1_oc8051_idata_n2369), .D(
        oc8051_ram_top1_oc8051_idata_n2370), .Y(
        oc8051_ram_top1_oc8051_idata_n2334) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3838 ( .A(
        oc8051_ram_top1_oc8051_idata_n506), .Y(
        oc8051_ram_top1_oc8051_idata_n2364) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3837 ( .A(
        oc8051_ram_top1_oc8051_idata_n514), .Y(
        oc8051_ram_top1_oc8051_idata_n2365) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3836 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n1061) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3835 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n1071) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3834 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1061), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1071), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2366) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3833 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2364), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2365), .C0(
        oc8051_ram_top1_oc8051_idata_n2366), .Y(
        oc8051_ram_top1_oc8051_idata_n2355) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3832 ( .A(
        oc8051_ram_top1_oc8051_idata_n490), .Y(
        oc8051_ram_top1_oc8051_idata_n2361) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3831 ( .A(
        oc8051_ram_top1_oc8051_idata_n498), .Y(
        oc8051_ram_top1_oc8051_idata_n2362) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3830 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n1035) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3829 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n1047) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3828 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1035), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1047), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2363) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3827 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2361), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2362), .C0(
        oc8051_ram_top1_oc8051_idata_n2363), .Y(
        oc8051_ram_top1_oc8051_idata_n2356) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3826 ( .A0(
        oc8051_ram_top1_oc8051_idata_n482), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n474), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2360) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3825 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2360), .Y(
        oc8051_ram_top1_oc8051_idata_n2357) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3824 ( .A0(
        oc8051_ram_top1_oc8051_idata_n466), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n458), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2359) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3823 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2359), .Y(
        oc8051_ram_top1_oc8051_idata_n2358) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3822 ( .A(
        oc8051_ram_top1_oc8051_idata_n2355), .B(
        oc8051_ram_top1_oc8051_idata_n2356), .C(
        oc8051_ram_top1_oc8051_idata_n2357), .D(
        oc8051_ram_top1_oc8051_idata_n2358), .Y(
        oc8051_ram_top1_oc8051_idata_n2335) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3821 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2351) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3820 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2352) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3819 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2353) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3818 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2354) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3817 ( .A(
        oc8051_ram_top1_oc8051_idata_n2351), .B(
        oc8051_ram_top1_oc8051_idata_n2352), .C(
        oc8051_ram_top1_oc8051_idata_n2353), .D(
        oc8051_ram_top1_oc8051_idata_n2354), .Y(
        oc8051_ram_top1_oc8051_idata_n2336) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3816 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2347) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3815 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2348) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3814 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2349) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3813 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2350) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3812 ( .A(
        oc8051_ram_top1_oc8051_idata_n2347), .B(
        oc8051_ram_top1_oc8051_idata_n2348), .C(
        oc8051_ram_top1_oc8051_idata_n2349), .D(
        oc8051_ram_top1_oc8051_idata_n2350), .Y(
        oc8051_ram_top1_oc8051_idata_n2337) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3811 ( .A0(
        oc8051_ram_top1_oc8051_idata_n450), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n442), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2346) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3810 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2346), .Y(
        oc8051_ram_top1_oc8051_idata_n2339) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3809 ( .A0(
        oc8051_ram_top1_oc8051_idata_n434), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n426), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2345) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3808 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2345), .Y(
        oc8051_ram_top1_oc8051_idata_n2340) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3807 ( .A0(
        oc8051_ram_top1_oc8051_idata_n418), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n410), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2344) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3806 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2344), .Y(
        oc8051_ram_top1_oc8051_idata_n2341) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3805 ( .A0(
        oc8051_ram_top1_oc8051_idata_n402), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n394), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2343) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3804 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2343), .Y(
        oc8051_ram_top1_oc8051_idata_n2342) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3803 ( .A(
        oc8051_ram_top1_oc8051_idata_n2339), .B(
        oc8051_ram_top1_oc8051_idata_n2340), .C(
        oc8051_ram_top1_oc8051_idata_n2341), .D(
        oc8051_ram_top1_oc8051_idata_n2342), .Y(
        oc8051_ram_top1_oc8051_idata_n2338) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3802 ( .A(
        oc8051_ram_top1_oc8051_idata_n2333), .B(
        oc8051_ram_top1_oc8051_idata_n2334), .C(
        oc8051_ram_top1_oc8051_idata_n2335), .D(
        oc8051_ram_top1_oc8051_idata_n2336), .E(
        oc8051_ram_top1_oc8051_idata_n2337), .F(
        oc8051_ram_top1_oc8051_idata_n2338), .Y(
        oc8051_ram_top1_oc8051_idata_n2332) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3801 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n2332), .B0(oc8051_ram_top1_rd_data_m[1]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n2201) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3800 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2328) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3799 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2329) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3798 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2330) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3797 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2331) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3796 ( .A(
        oc8051_ram_top1_oc8051_idata_n2328), .B(
        oc8051_ram_top1_oc8051_idata_n2329), .C(
        oc8051_ram_top1_oc8051_idata_n2330), .D(
        oc8051_ram_top1_oc8051_idata_n2331), .Y(
        oc8051_ram_top1_oc8051_idata_n2290) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3795 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2324) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3794 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2325) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3793 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2326) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3792 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2327) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3791 ( .A(
        oc8051_ram_top1_oc8051_idata_n2324), .B(
        oc8051_ram_top1_oc8051_idata_n2325), .C(
        oc8051_ram_top1_oc8051_idata_n2326), .D(
        oc8051_ram_top1_oc8051_idata_n2327), .Y(
        oc8051_ram_top1_oc8051_idata_n2291) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3790 ( .A(
        oc8051_ram_top1_oc8051_idata_n378), .Y(
        oc8051_ram_top1_oc8051_idata_n2321) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3789 ( .A(
        oc8051_ram_top1_oc8051_idata_n386), .Y(
        oc8051_ram_top1_oc8051_idata_n2322) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3788 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n953) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3787 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n962) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3786 ( .A0(
        oc8051_ram_top1_oc8051_idata_n953), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n962), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2323) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3785 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2321), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2322), .C0(
        oc8051_ram_top1_oc8051_idata_n2323), .Y(
        oc8051_ram_top1_oc8051_idata_n2312) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3784 ( .A(
        oc8051_ram_top1_oc8051_idata_n362), .Y(
        oc8051_ram_top1_oc8051_idata_n2318) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3783 ( .A(
        oc8051_ram_top1_oc8051_idata_n370), .Y(
        oc8051_ram_top1_oc8051_idata_n2319) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3782 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n932) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3781 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n942) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3780 ( .A0(
        oc8051_ram_top1_oc8051_idata_n932), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n942), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2320) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3779 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2318), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2319), .C0(
        oc8051_ram_top1_oc8051_idata_n2320), .Y(
        oc8051_ram_top1_oc8051_idata_n2313) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3778 ( .A0(
        oc8051_ram_top1_oc8051_idata_n354), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n346), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2317) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3777 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2317), .Y(
        oc8051_ram_top1_oc8051_idata_n2314) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3776 ( .A0(
        oc8051_ram_top1_oc8051_idata_n338), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n330), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2316) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3775 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2316), .Y(
        oc8051_ram_top1_oc8051_idata_n2315) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3774 ( .A(
        oc8051_ram_top1_oc8051_idata_n2312), .B(
        oc8051_ram_top1_oc8051_idata_n2313), .C(
        oc8051_ram_top1_oc8051_idata_n2314), .D(
        oc8051_ram_top1_oc8051_idata_n2315), .Y(
        oc8051_ram_top1_oc8051_idata_n2292) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3773 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2308) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3772 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2309) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3771 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2310) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3770 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2311) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3769 ( .A(
        oc8051_ram_top1_oc8051_idata_n2308), .B(
        oc8051_ram_top1_oc8051_idata_n2309), .C(
        oc8051_ram_top1_oc8051_idata_n2310), .D(
        oc8051_ram_top1_oc8051_idata_n2311), .Y(
        oc8051_ram_top1_oc8051_idata_n2293) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3768 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2304) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3767 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2305) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3766 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2306) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3765 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2307) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3764 ( .A(
        oc8051_ram_top1_oc8051_idata_n2304), .B(
        oc8051_ram_top1_oc8051_idata_n2305), .C(
        oc8051_ram_top1_oc8051_idata_n2306), .D(
        oc8051_ram_top1_oc8051_idata_n2307), .Y(
        oc8051_ram_top1_oc8051_idata_n2294) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3763 ( .A0(
        oc8051_ram_top1_oc8051_idata_n322), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n314), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2303) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3762 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2303), .Y(
        oc8051_ram_top1_oc8051_idata_n2296) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3761 ( .A0(
        oc8051_ram_top1_oc8051_idata_n306), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n298), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2302) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3760 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2302), .Y(
        oc8051_ram_top1_oc8051_idata_n2297) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3759 ( .A0(
        oc8051_ram_top1_oc8051_idata_n290), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n282), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2301) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3758 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2301), .Y(
        oc8051_ram_top1_oc8051_idata_n2298) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3757 ( .A0(
        oc8051_ram_top1_oc8051_idata_n274), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n266), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2300) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3756 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2300), .Y(
        oc8051_ram_top1_oc8051_idata_n2299) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3755 ( .A(
        oc8051_ram_top1_oc8051_idata_n2296), .B(
        oc8051_ram_top1_oc8051_idata_n2297), .C(
        oc8051_ram_top1_oc8051_idata_n2298), .D(
        oc8051_ram_top1_oc8051_idata_n2299), .Y(
        oc8051_ram_top1_oc8051_idata_n2295) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3754 ( .A(
        oc8051_ram_top1_oc8051_idata_n2290), .B(
        oc8051_ram_top1_oc8051_idata_n2291), .C(
        oc8051_ram_top1_oc8051_idata_n2292), .D(
        oc8051_ram_top1_oc8051_idata_n2293), .E(
        oc8051_ram_top1_oc8051_idata_n2294), .F(
        oc8051_ram_top1_oc8051_idata_n2295), .Y(
        oc8051_ram_top1_oc8051_idata_n2203) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3753 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2286) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3752 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2287) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3751 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2288) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3750 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2289) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3749 ( .A(
        oc8051_ram_top1_oc8051_idata_n2286), .B(
        oc8051_ram_top1_oc8051_idata_n2287), .C(
        oc8051_ram_top1_oc8051_idata_n2288), .D(
        oc8051_ram_top1_oc8051_idata_n2289), .Y(
        oc8051_ram_top1_oc8051_idata_n2248) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3748 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2282) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3747 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2283) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3746 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2284) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3745 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2285) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3744 ( .A(
        oc8051_ram_top1_oc8051_idata_n2282), .B(
        oc8051_ram_top1_oc8051_idata_n2283), .C(
        oc8051_ram_top1_oc8051_idata_n2284), .D(
        oc8051_ram_top1_oc8051_idata_n2285), .Y(
        oc8051_ram_top1_oc8051_idata_n2249) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3743 ( .A(
        oc8051_ram_top1_oc8051_idata_n250), .Y(
        oc8051_ram_top1_oc8051_idata_n2279) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3742 ( .A(
        oc8051_ram_top1_oc8051_idata_n258), .Y(
        oc8051_ram_top1_oc8051_idata_n2280) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3741 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n851) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3740 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n860) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3739 ( .A0(
        oc8051_ram_top1_oc8051_idata_n851), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n860), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2281) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3738 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2279), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2280), .C0(
        oc8051_ram_top1_oc8051_idata_n2281), .Y(
        oc8051_ram_top1_oc8051_idata_n2270) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3737 ( .A(
        oc8051_ram_top1_oc8051_idata_n234), .Y(
        oc8051_ram_top1_oc8051_idata_n2276) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3736 ( .A(
        oc8051_ram_top1_oc8051_idata_n242), .Y(
        oc8051_ram_top1_oc8051_idata_n2277) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3735 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n830) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3734 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n840) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3733 ( .A0(
        oc8051_ram_top1_oc8051_idata_n830), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n840), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2278) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3732 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2276), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2277), .C0(
        oc8051_ram_top1_oc8051_idata_n2278), .Y(
        oc8051_ram_top1_oc8051_idata_n2271) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3731 ( .A0(
        oc8051_ram_top1_oc8051_idata_n226), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n218), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2275) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3730 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2275), .Y(
        oc8051_ram_top1_oc8051_idata_n2272) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3729 ( .A0(
        oc8051_ram_top1_oc8051_idata_n210), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n202), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2274) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3728 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2274), .Y(
        oc8051_ram_top1_oc8051_idata_n2273) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3727 ( .A(
        oc8051_ram_top1_oc8051_idata_n2270), .B(
        oc8051_ram_top1_oc8051_idata_n2271), .C(
        oc8051_ram_top1_oc8051_idata_n2272), .D(
        oc8051_ram_top1_oc8051_idata_n2273), .Y(
        oc8051_ram_top1_oc8051_idata_n2250) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3726 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2266) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3725 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2267) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3724 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2268) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3723 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2269) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3722 ( .A(
        oc8051_ram_top1_oc8051_idata_n2266), .B(
        oc8051_ram_top1_oc8051_idata_n2267), .C(
        oc8051_ram_top1_oc8051_idata_n2268), .D(
        oc8051_ram_top1_oc8051_idata_n2269), .Y(
        oc8051_ram_top1_oc8051_idata_n2251) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3721 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2262) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3720 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2263) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3719 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2264) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3718 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2265) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3717 ( .A(
        oc8051_ram_top1_oc8051_idata_n2262), .B(
        oc8051_ram_top1_oc8051_idata_n2263), .C(
        oc8051_ram_top1_oc8051_idata_n2264), .D(
        oc8051_ram_top1_oc8051_idata_n2265), .Y(
        oc8051_ram_top1_oc8051_idata_n2252) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3716 ( .A0(
        oc8051_ram_top1_oc8051_idata_n194), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n186), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2261) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3715 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2261), .Y(
        oc8051_ram_top1_oc8051_idata_n2254) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3714 ( .A0(
        oc8051_ram_top1_oc8051_idata_n178), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n170), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2260) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3713 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2260), .Y(
        oc8051_ram_top1_oc8051_idata_n2255) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3712 ( .A0(
        oc8051_ram_top1_oc8051_idata_n162), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n154), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2259) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3711 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2259), .Y(
        oc8051_ram_top1_oc8051_idata_n2256) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3710 ( .A0(
        oc8051_ram_top1_oc8051_idata_n146), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n138), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2258) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3709 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2258), .Y(
        oc8051_ram_top1_oc8051_idata_n2257) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3708 ( .A(
        oc8051_ram_top1_oc8051_idata_n2254), .B(
        oc8051_ram_top1_oc8051_idata_n2255), .C(
        oc8051_ram_top1_oc8051_idata_n2256), .D(
        oc8051_ram_top1_oc8051_idata_n2257), .Y(
        oc8051_ram_top1_oc8051_idata_n2253) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3707 ( .A(
        oc8051_ram_top1_oc8051_idata_n2248), .B(
        oc8051_ram_top1_oc8051_idata_n2249), .C(
        oc8051_ram_top1_oc8051_idata_n2250), .D(
        oc8051_ram_top1_oc8051_idata_n2251), .E(
        oc8051_ram_top1_oc8051_idata_n2252), .F(
        oc8051_ram_top1_oc8051_idata_n2253), .Y(
        oc8051_ram_top1_oc8051_idata_n2204) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3706 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2244) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3705 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2245) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3704 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2246) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3703 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2247) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3702 ( .A(
        oc8051_ram_top1_oc8051_idata_n2244), .B(
        oc8051_ram_top1_oc8051_idata_n2245), .C(
        oc8051_ram_top1_oc8051_idata_n2246), .D(
        oc8051_ram_top1_oc8051_idata_n2247), .Y(
        oc8051_ram_top1_oc8051_idata_n2206) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3701 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2240) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3700 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2241) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3699 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2242) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3698 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2243) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3697 ( .A(
        oc8051_ram_top1_oc8051_idata_n2240), .B(
        oc8051_ram_top1_oc8051_idata_n2241), .C(
        oc8051_ram_top1_oc8051_idata_n2242), .D(
        oc8051_ram_top1_oc8051_idata_n2243), .Y(
        oc8051_ram_top1_oc8051_idata_n2207) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3696 ( .A(
        oc8051_ram_top1_oc8051_idata_n122), .Y(
        oc8051_ram_top1_oc8051_idata_n2237) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3695 ( .A(
        oc8051_ram_top1_oc8051_idata_n130), .Y(
        oc8051_ram_top1_oc8051_idata_n2238) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3694 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n748) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3693 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n757) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3692 ( .A0(
        oc8051_ram_top1_oc8051_idata_n748), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n757), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2239) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3691 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2237), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2238), .C0(
        oc8051_ram_top1_oc8051_idata_n2239), .Y(
        oc8051_ram_top1_oc8051_idata_n2228) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3690 ( .A(
        oc8051_ram_top1_oc8051_idata_n106), .Y(
        oc8051_ram_top1_oc8051_idata_n2234) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3689 ( .A(
        oc8051_ram_top1_oc8051_idata_n114), .Y(
        oc8051_ram_top1_oc8051_idata_n2235) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3688 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n727) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3687 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n737) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3686 ( .A0(
        oc8051_ram_top1_oc8051_idata_n727), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n737), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2236) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3685 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2234), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2235), .C0(
        oc8051_ram_top1_oc8051_idata_n2236), .Y(
        oc8051_ram_top1_oc8051_idata_n2229) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3684 ( .A0(
        oc8051_ram_top1_oc8051_idata_n98), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n90), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2233) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3683 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2233), .Y(
        oc8051_ram_top1_oc8051_idata_n2230) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3682 ( .A0(
        oc8051_ram_top1_oc8051_idata_n82), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n74), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2232) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3681 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2232), .Y(
        oc8051_ram_top1_oc8051_idata_n2231) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3680 ( .A(
        oc8051_ram_top1_oc8051_idata_n2228), .B(
        oc8051_ram_top1_oc8051_idata_n2229), .C(
        oc8051_ram_top1_oc8051_idata_n2230), .D(
        oc8051_ram_top1_oc8051_idata_n2231), .Y(
        oc8051_ram_top1_oc8051_idata_n2208) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3679 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2224) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3678 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2225) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3677 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2226) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3676 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2227) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3675 ( .A(
        oc8051_ram_top1_oc8051_idata_n2224), .B(
        oc8051_ram_top1_oc8051_idata_n2225), .C(
        oc8051_ram_top1_oc8051_idata_n2226), .D(
        oc8051_ram_top1_oc8051_idata_n2227), .Y(
        oc8051_ram_top1_oc8051_idata_n2209) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3674 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2220) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3673 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2221) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3672 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2222) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3671 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__1_), .Y(
        oc8051_ram_top1_oc8051_idata_n2223) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3670 ( .A(
        oc8051_ram_top1_oc8051_idata_n2220), .B(
        oc8051_ram_top1_oc8051_idata_n2221), .C(
        oc8051_ram_top1_oc8051_idata_n2222), .D(
        oc8051_ram_top1_oc8051_idata_n2223), .Y(
        oc8051_ram_top1_oc8051_idata_n2210) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3669 ( .A0(
        oc8051_ram_top1_oc8051_idata_n66), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n58), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2219) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3668 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2219), .Y(
        oc8051_ram_top1_oc8051_idata_n2212) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3667 ( .A0(
        oc8051_ram_top1_oc8051_idata_n50), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n42), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2218) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3666 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2218), .Y(
        oc8051_ram_top1_oc8051_idata_n2213) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3665 ( .A0(
        oc8051_ram_top1_oc8051_idata_n34), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n26), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2217) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3664 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2217), .Y(
        oc8051_ram_top1_oc8051_idata_n2214) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3663 ( .A0(
        oc8051_ram_top1_oc8051_idata_n18), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n10), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2216) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3662 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__1_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__1_), .C0(
        oc8051_ram_top1_oc8051_idata_n2216), .Y(
        oc8051_ram_top1_oc8051_idata_n2215) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3661 ( .A(
        oc8051_ram_top1_oc8051_idata_n2212), .B(
        oc8051_ram_top1_oc8051_idata_n2213), .C(
        oc8051_ram_top1_oc8051_idata_n2214), .D(
        oc8051_ram_top1_oc8051_idata_n2215), .Y(
        oc8051_ram_top1_oc8051_idata_n2211) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3660 ( .A(
        oc8051_ram_top1_oc8051_idata_n2206), .B(
        oc8051_ram_top1_oc8051_idata_n2207), .C(
        oc8051_ram_top1_oc8051_idata_n2208), .D(
        oc8051_ram_top1_oc8051_idata_n2209), .E(
        oc8051_ram_top1_oc8051_idata_n2210), .F(
        oc8051_ram_top1_oc8051_idata_n2211), .Y(
        oc8051_ram_top1_oc8051_idata_n2205) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3659 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n2203), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n2204), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n2205), .Y(
        oc8051_ram_top1_oc8051_idata_n2202) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3658 ( .A0(
        oc8051_ram_top1_oc8051_idata_n545), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n2201), .C0(
        oc8051_ram_top1_oc8051_idata_n2202), .Y(
        oc8051_ram_top1_oc8051_idata_n2476) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3657 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2197) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3656 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2198) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3655 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2199) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3654 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2200) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3653 ( .A(
        oc8051_ram_top1_oc8051_idata_n2197), .B(
        oc8051_ram_top1_oc8051_idata_n2198), .C(
        oc8051_ram_top1_oc8051_idata_n2199), .D(
        oc8051_ram_top1_oc8051_idata_n2200), .Y(
        oc8051_ram_top1_oc8051_idata_n2159) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3652 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2193) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3651 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2194) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3650 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2195) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3649 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2196) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3648 ( .A(
        oc8051_ram_top1_oc8051_idata_n2193), .B(
        oc8051_ram_top1_oc8051_idata_n2194), .C(
        oc8051_ram_top1_oc8051_idata_n2195), .D(
        oc8051_ram_top1_oc8051_idata_n2196), .Y(
        oc8051_ram_top1_oc8051_idata_n2160) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3647 ( .A(
        oc8051_ram_top1_oc8051_idata_n505), .Y(
        oc8051_ram_top1_oc8051_idata_n2190) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3646 ( .A(
        oc8051_ram_top1_oc8051_idata_n513), .Y(
        oc8051_ram_top1_oc8051_idata_n2191) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3645 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n1060) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3644 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n1070) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3643 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1060), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1070), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2192) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3642 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2190), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2191), .C0(
        oc8051_ram_top1_oc8051_idata_n2192), .Y(
        oc8051_ram_top1_oc8051_idata_n2181) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3641 ( .A(
        oc8051_ram_top1_oc8051_idata_n489), .Y(
        oc8051_ram_top1_oc8051_idata_n2187) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3640 ( .A(
        oc8051_ram_top1_oc8051_idata_n497), .Y(
        oc8051_ram_top1_oc8051_idata_n2188) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3639 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n1034) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3638 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n1046) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3637 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1034), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1046), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2189) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3636 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2187), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2188), .C0(
        oc8051_ram_top1_oc8051_idata_n2189), .Y(
        oc8051_ram_top1_oc8051_idata_n2182) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3635 ( .A0(
        oc8051_ram_top1_oc8051_idata_n481), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n473), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2186) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3634 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2186), .Y(
        oc8051_ram_top1_oc8051_idata_n2183) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3633 ( .A0(
        oc8051_ram_top1_oc8051_idata_n465), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n457), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2185) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3632 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2185), .Y(
        oc8051_ram_top1_oc8051_idata_n2184) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3631 ( .A(
        oc8051_ram_top1_oc8051_idata_n2181), .B(
        oc8051_ram_top1_oc8051_idata_n2182), .C(
        oc8051_ram_top1_oc8051_idata_n2183), .D(
        oc8051_ram_top1_oc8051_idata_n2184), .Y(
        oc8051_ram_top1_oc8051_idata_n2161) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3630 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2177) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3629 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2178) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3628 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2179) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3627 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2180) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3626 ( .A(
        oc8051_ram_top1_oc8051_idata_n2177), .B(
        oc8051_ram_top1_oc8051_idata_n2178), .C(
        oc8051_ram_top1_oc8051_idata_n2179), .D(
        oc8051_ram_top1_oc8051_idata_n2180), .Y(
        oc8051_ram_top1_oc8051_idata_n2162) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3625 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2173) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3624 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2174) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3623 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2175) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3622 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2176) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3621 ( .A(
        oc8051_ram_top1_oc8051_idata_n2173), .B(
        oc8051_ram_top1_oc8051_idata_n2174), .C(
        oc8051_ram_top1_oc8051_idata_n2175), .D(
        oc8051_ram_top1_oc8051_idata_n2176), .Y(
        oc8051_ram_top1_oc8051_idata_n2163) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3620 ( .A0(
        oc8051_ram_top1_oc8051_idata_n449), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n441), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2172) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3619 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2172), .Y(
        oc8051_ram_top1_oc8051_idata_n2165) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3618 ( .A0(
        oc8051_ram_top1_oc8051_idata_n433), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n425), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2171) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3617 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2171), .Y(
        oc8051_ram_top1_oc8051_idata_n2166) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3616 ( .A0(
        oc8051_ram_top1_oc8051_idata_n417), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n409), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2170) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3615 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2170), .Y(
        oc8051_ram_top1_oc8051_idata_n2167) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3614 ( .A0(
        oc8051_ram_top1_oc8051_idata_n401), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n393), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2169) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3613 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2169), .Y(
        oc8051_ram_top1_oc8051_idata_n2168) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3612 ( .A(
        oc8051_ram_top1_oc8051_idata_n2165), .B(
        oc8051_ram_top1_oc8051_idata_n2166), .C(
        oc8051_ram_top1_oc8051_idata_n2167), .D(
        oc8051_ram_top1_oc8051_idata_n2168), .Y(
        oc8051_ram_top1_oc8051_idata_n2164) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3611 ( .A(
        oc8051_ram_top1_oc8051_idata_n2159), .B(
        oc8051_ram_top1_oc8051_idata_n2160), .C(
        oc8051_ram_top1_oc8051_idata_n2161), .D(
        oc8051_ram_top1_oc8051_idata_n2162), .E(
        oc8051_ram_top1_oc8051_idata_n2163), .F(
        oc8051_ram_top1_oc8051_idata_n2164), .Y(
        oc8051_ram_top1_oc8051_idata_n2158) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3610 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n2158), .B0(oc8051_ram_top1_rd_data_m[2]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n2027) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3609 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2154) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3608 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2155) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3607 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2156) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3606 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2157) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3605 ( .A(
        oc8051_ram_top1_oc8051_idata_n2154), .B(
        oc8051_ram_top1_oc8051_idata_n2155), .C(
        oc8051_ram_top1_oc8051_idata_n2156), .D(
        oc8051_ram_top1_oc8051_idata_n2157), .Y(
        oc8051_ram_top1_oc8051_idata_n2116) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3604 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2150) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3603 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2151) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3602 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2152) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3601 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2153) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3600 ( .A(
        oc8051_ram_top1_oc8051_idata_n2150), .B(
        oc8051_ram_top1_oc8051_idata_n2151), .C(
        oc8051_ram_top1_oc8051_idata_n2152), .D(
        oc8051_ram_top1_oc8051_idata_n2153), .Y(
        oc8051_ram_top1_oc8051_idata_n2117) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3599 ( .A(
        oc8051_ram_top1_oc8051_idata_n377), .Y(
        oc8051_ram_top1_oc8051_idata_n2147) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3598 ( .A(
        oc8051_ram_top1_oc8051_idata_n385), .Y(
        oc8051_ram_top1_oc8051_idata_n2148) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3597 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n952) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3596 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n961) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3595 ( .A0(
        oc8051_ram_top1_oc8051_idata_n952), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n961), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2149) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3594 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2147), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2148), .C0(
        oc8051_ram_top1_oc8051_idata_n2149), .Y(
        oc8051_ram_top1_oc8051_idata_n2138) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3593 ( .A(
        oc8051_ram_top1_oc8051_idata_n361), .Y(
        oc8051_ram_top1_oc8051_idata_n2144) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3592 ( .A(
        oc8051_ram_top1_oc8051_idata_n369), .Y(
        oc8051_ram_top1_oc8051_idata_n2145) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3591 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n931) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3590 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n941) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3589 ( .A0(
        oc8051_ram_top1_oc8051_idata_n931), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n941), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2146) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3588 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2144), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2145), .C0(
        oc8051_ram_top1_oc8051_idata_n2146), .Y(
        oc8051_ram_top1_oc8051_idata_n2139) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3587 ( .A0(
        oc8051_ram_top1_oc8051_idata_n353), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n345), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2143) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3586 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2143), .Y(
        oc8051_ram_top1_oc8051_idata_n2140) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3585 ( .A0(
        oc8051_ram_top1_oc8051_idata_n337), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n329), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2142) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3584 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2142), .Y(
        oc8051_ram_top1_oc8051_idata_n2141) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3583 ( .A(
        oc8051_ram_top1_oc8051_idata_n2138), .B(
        oc8051_ram_top1_oc8051_idata_n2139), .C(
        oc8051_ram_top1_oc8051_idata_n2140), .D(
        oc8051_ram_top1_oc8051_idata_n2141), .Y(
        oc8051_ram_top1_oc8051_idata_n2118) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3582 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2134) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3581 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2135) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3580 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2136) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3579 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2137) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3578 ( .A(
        oc8051_ram_top1_oc8051_idata_n2134), .B(
        oc8051_ram_top1_oc8051_idata_n2135), .C(
        oc8051_ram_top1_oc8051_idata_n2136), .D(
        oc8051_ram_top1_oc8051_idata_n2137), .Y(
        oc8051_ram_top1_oc8051_idata_n2119) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3577 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2130) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3576 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2131) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3575 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2132) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3574 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2133) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3573 ( .A(
        oc8051_ram_top1_oc8051_idata_n2130), .B(
        oc8051_ram_top1_oc8051_idata_n2131), .C(
        oc8051_ram_top1_oc8051_idata_n2132), .D(
        oc8051_ram_top1_oc8051_idata_n2133), .Y(
        oc8051_ram_top1_oc8051_idata_n2120) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3572 ( .A0(
        oc8051_ram_top1_oc8051_idata_n321), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n313), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2129) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3571 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2129), .Y(
        oc8051_ram_top1_oc8051_idata_n2122) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3570 ( .A0(
        oc8051_ram_top1_oc8051_idata_n305), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n297), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2128) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3569 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2128), .Y(
        oc8051_ram_top1_oc8051_idata_n2123) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3568 ( .A0(
        oc8051_ram_top1_oc8051_idata_n289), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n281), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2127) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3567 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2127), .Y(
        oc8051_ram_top1_oc8051_idata_n2124) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3566 ( .A0(
        oc8051_ram_top1_oc8051_idata_n273), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n265), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2126) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3565 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2126), .Y(
        oc8051_ram_top1_oc8051_idata_n2125) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3564 ( .A(
        oc8051_ram_top1_oc8051_idata_n2122), .B(
        oc8051_ram_top1_oc8051_idata_n2123), .C(
        oc8051_ram_top1_oc8051_idata_n2124), .D(
        oc8051_ram_top1_oc8051_idata_n2125), .Y(
        oc8051_ram_top1_oc8051_idata_n2121) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3563 ( .A(
        oc8051_ram_top1_oc8051_idata_n2116), .B(
        oc8051_ram_top1_oc8051_idata_n2117), .C(
        oc8051_ram_top1_oc8051_idata_n2118), .D(
        oc8051_ram_top1_oc8051_idata_n2119), .E(
        oc8051_ram_top1_oc8051_idata_n2120), .F(
        oc8051_ram_top1_oc8051_idata_n2121), .Y(
        oc8051_ram_top1_oc8051_idata_n2029) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3562 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2112) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3561 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2113) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3560 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2114) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3559 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2115) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3558 ( .A(
        oc8051_ram_top1_oc8051_idata_n2112), .B(
        oc8051_ram_top1_oc8051_idata_n2113), .C(
        oc8051_ram_top1_oc8051_idata_n2114), .D(
        oc8051_ram_top1_oc8051_idata_n2115), .Y(
        oc8051_ram_top1_oc8051_idata_n2074) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3557 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2108) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3556 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2109) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3555 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2110) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3554 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2111) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3553 ( .A(
        oc8051_ram_top1_oc8051_idata_n2108), .B(
        oc8051_ram_top1_oc8051_idata_n2109), .C(
        oc8051_ram_top1_oc8051_idata_n2110), .D(
        oc8051_ram_top1_oc8051_idata_n2111), .Y(
        oc8051_ram_top1_oc8051_idata_n2075) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3552 ( .A(
        oc8051_ram_top1_oc8051_idata_n249), .Y(
        oc8051_ram_top1_oc8051_idata_n2105) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3551 ( .A(
        oc8051_ram_top1_oc8051_idata_n257), .Y(
        oc8051_ram_top1_oc8051_idata_n2106) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3550 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n850) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3549 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n859) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3548 ( .A0(
        oc8051_ram_top1_oc8051_idata_n850), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n859), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2107) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3547 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2105), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2106), .C0(
        oc8051_ram_top1_oc8051_idata_n2107), .Y(
        oc8051_ram_top1_oc8051_idata_n2096) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3546 ( .A(
        oc8051_ram_top1_oc8051_idata_n233), .Y(
        oc8051_ram_top1_oc8051_idata_n2102) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3545 ( .A(
        oc8051_ram_top1_oc8051_idata_n241), .Y(
        oc8051_ram_top1_oc8051_idata_n2103) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3544 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n829) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3543 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n839) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3542 ( .A0(
        oc8051_ram_top1_oc8051_idata_n829), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n839), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2104) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3541 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2102), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2103), .C0(
        oc8051_ram_top1_oc8051_idata_n2104), .Y(
        oc8051_ram_top1_oc8051_idata_n2097) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3540 ( .A0(
        oc8051_ram_top1_oc8051_idata_n225), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n217), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2101) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3539 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2101), .Y(
        oc8051_ram_top1_oc8051_idata_n2098) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3538 ( .A0(
        oc8051_ram_top1_oc8051_idata_n209), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n201), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2100) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3537 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2100), .Y(
        oc8051_ram_top1_oc8051_idata_n2099) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3536 ( .A(
        oc8051_ram_top1_oc8051_idata_n2096), .B(
        oc8051_ram_top1_oc8051_idata_n2097), .C(
        oc8051_ram_top1_oc8051_idata_n2098), .D(
        oc8051_ram_top1_oc8051_idata_n2099), .Y(
        oc8051_ram_top1_oc8051_idata_n2076) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3535 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2092) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3534 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2093) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3533 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2094) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3532 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2095) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3531 ( .A(
        oc8051_ram_top1_oc8051_idata_n2092), .B(
        oc8051_ram_top1_oc8051_idata_n2093), .C(
        oc8051_ram_top1_oc8051_idata_n2094), .D(
        oc8051_ram_top1_oc8051_idata_n2095), .Y(
        oc8051_ram_top1_oc8051_idata_n2077) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3530 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2088) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3529 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2089) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3528 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2090) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3527 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2091) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3526 ( .A(
        oc8051_ram_top1_oc8051_idata_n2088), .B(
        oc8051_ram_top1_oc8051_idata_n2089), .C(
        oc8051_ram_top1_oc8051_idata_n2090), .D(
        oc8051_ram_top1_oc8051_idata_n2091), .Y(
        oc8051_ram_top1_oc8051_idata_n2078) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3525 ( .A0(
        oc8051_ram_top1_oc8051_idata_n193), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n185), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2087) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3524 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2087), .Y(
        oc8051_ram_top1_oc8051_idata_n2080) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3523 ( .A0(
        oc8051_ram_top1_oc8051_idata_n177), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n169), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2086) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3522 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2086), .Y(
        oc8051_ram_top1_oc8051_idata_n2081) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3521 ( .A0(
        oc8051_ram_top1_oc8051_idata_n161), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n153), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2085) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3520 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2085), .Y(
        oc8051_ram_top1_oc8051_idata_n2082) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3519 ( .A0(
        oc8051_ram_top1_oc8051_idata_n145), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n137), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2084) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3518 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2084), .Y(
        oc8051_ram_top1_oc8051_idata_n2083) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3517 ( .A(
        oc8051_ram_top1_oc8051_idata_n2080), .B(
        oc8051_ram_top1_oc8051_idata_n2081), .C(
        oc8051_ram_top1_oc8051_idata_n2082), .D(
        oc8051_ram_top1_oc8051_idata_n2083), .Y(
        oc8051_ram_top1_oc8051_idata_n2079) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3516 ( .A(
        oc8051_ram_top1_oc8051_idata_n2074), .B(
        oc8051_ram_top1_oc8051_idata_n2075), .C(
        oc8051_ram_top1_oc8051_idata_n2076), .D(
        oc8051_ram_top1_oc8051_idata_n2077), .E(
        oc8051_ram_top1_oc8051_idata_n2078), .F(
        oc8051_ram_top1_oc8051_idata_n2079), .Y(
        oc8051_ram_top1_oc8051_idata_n2030) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3515 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2070) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3514 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2071) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3513 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2072) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3512 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2073) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3511 ( .A(
        oc8051_ram_top1_oc8051_idata_n2070), .B(
        oc8051_ram_top1_oc8051_idata_n2071), .C(
        oc8051_ram_top1_oc8051_idata_n2072), .D(
        oc8051_ram_top1_oc8051_idata_n2073), .Y(
        oc8051_ram_top1_oc8051_idata_n2032) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3510 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2066) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3509 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2067) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3508 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2068) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3507 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2069) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3506 ( .A(
        oc8051_ram_top1_oc8051_idata_n2066), .B(
        oc8051_ram_top1_oc8051_idata_n2067), .C(
        oc8051_ram_top1_oc8051_idata_n2068), .D(
        oc8051_ram_top1_oc8051_idata_n2069), .Y(
        oc8051_ram_top1_oc8051_idata_n2033) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3505 ( .A(
        oc8051_ram_top1_oc8051_idata_n121), .Y(
        oc8051_ram_top1_oc8051_idata_n2063) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3504 ( .A(
        oc8051_ram_top1_oc8051_idata_n129), .Y(
        oc8051_ram_top1_oc8051_idata_n2064) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3503 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n747) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3502 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n756) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3501 ( .A0(
        oc8051_ram_top1_oc8051_idata_n747), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n756), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2065) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3500 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2063), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2064), .C0(
        oc8051_ram_top1_oc8051_idata_n2065), .Y(
        oc8051_ram_top1_oc8051_idata_n2054) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3499 ( .A(
        oc8051_ram_top1_oc8051_idata_n105), .Y(
        oc8051_ram_top1_oc8051_idata_n2060) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3498 ( .A(
        oc8051_ram_top1_oc8051_idata_n113), .Y(
        oc8051_ram_top1_oc8051_idata_n2061) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3497 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n726) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3496 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n736) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3495 ( .A0(
        oc8051_ram_top1_oc8051_idata_n726), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n736), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2062) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3494 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2060), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2061), .C0(
        oc8051_ram_top1_oc8051_idata_n2062), .Y(
        oc8051_ram_top1_oc8051_idata_n2055) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3493 ( .A0(
        oc8051_ram_top1_oc8051_idata_n97), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n89), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2059) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3492 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2059), .Y(
        oc8051_ram_top1_oc8051_idata_n2056) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3491 ( .A0(
        oc8051_ram_top1_oc8051_idata_n81), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n73), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2058) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3490 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2058), .Y(
        oc8051_ram_top1_oc8051_idata_n2057) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3489 ( .A(
        oc8051_ram_top1_oc8051_idata_n2054), .B(
        oc8051_ram_top1_oc8051_idata_n2055), .C(
        oc8051_ram_top1_oc8051_idata_n2056), .D(
        oc8051_ram_top1_oc8051_idata_n2057), .Y(
        oc8051_ram_top1_oc8051_idata_n2034) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3488 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2050) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3487 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2051) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3486 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2052) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3485 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2053) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3484 ( .A(
        oc8051_ram_top1_oc8051_idata_n2050), .B(
        oc8051_ram_top1_oc8051_idata_n2051), .C(
        oc8051_ram_top1_oc8051_idata_n2052), .D(
        oc8051_ram_top1_oc8051_idata_n2053), .Y(
        oc8051_ram_top1_oc8051_idata_n2035) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3483 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2046) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3482 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2047) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3481 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2048) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3480 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__2_), .Y(
        oc8051_ram_top1_oc8051_idata_n2049) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3479 ( .A(
        oc8051_ram_top1_oc8051_idata_n2046), .B(
        oc8051_ram_top1_oc8051_idata_n2047), .C(
        oc8051_ram_top1_oc8051_idata_n2048), .D(
        oc8051_ram_top1_oc8051_idata_n2049), .Y(
        oc8051_ram_top1_oc8051_idata_n2036) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3478 ( .A0(
        oc8051_ram_top1_oc8051_idata_n65), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n57), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n2045) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3477 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2045), .Y(
        oc8051_ram_top1_oc8051_idata_n2038) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3476 ( .A0(
        oc8051_ram_top1_oc8051_idata_n49), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n41), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n2044) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3475 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2044), .Y(
        oc8051_ram_top1_oc8051_idata_n2039) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3474 ( .A0(
        oc8051_ram_top1_oc8051_idata_n33), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n25), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n2043) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3473 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2043), .Y(
        oc8051_ram_top1_oc8051_idata_n2040) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3472 ( .A0(
        oc8051_ram_top1_oc8051_idata_n17), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n9), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n2042) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3471 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__2_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__2_), .C0(
        oc8051_ram_top1_oc8051_idata_n2042), .Y(
        oc8051_ram_top1_oc8051_idata_n2041) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3470 ( .A(
        oc8051_ram_top1_oc8051_idata_n2038), .B(
        oc8051_ram_top1_oc8051_idata_n2039), .C(
        oc8051_ram_top1_oc8051_idata_n2040), .D(
        oc8051_ram_top1_oc8051_idata_n2041), .Y(
        oc8051_ram_top1_oc8051_idata_n2037) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3469 ( .A(
        oc8051_ram_top1_oc8051_idata_n2032), .B(
        oc8051_ram_top1_oc8051_idata_n2033), .C(
        oc8051_ram_top1_oc8051_idata_n2034), .D(
        oc8051_ram_top1_oc8051_idata_n2035), .E(
        oc8051_ram_top1_oc8051_idata_n2036), .F(
        oc8051_ram_top1_oc8051_idata_n2037), .Y(
        oc8051_ram_top1_oc8051_idata_n2031) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3468 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n2029), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n2030), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n2031), .Y(
        oc8051_ram_top1_oc8051_idata_n2028) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3467 ( .A0(
        oc8051_ram_top1_oc8051_idata_n562), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n2027), .C0(
        oc8051_ram_top1_oc8051_idata_n2028), .Y(
        oc8051_ram_top1_oc8051_idata_n2477) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3466 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2023) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3465 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2024) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3464 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2025) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3463 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2026) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3462 ( .A(
        oc8051_ram_top1_oc8051_idata_n2023), .B(
        oc8051_ram_top1_oc8051_idata_n2024), .C(
        oc8051_ram_top1_oc8051_idata_n2025), .D(
        oc8051_ram_top1_oc8051_idata_n2026), .Y(
        oc8051_ram_top1_oc8051_idata_n1985) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3461 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2019) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3460 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2020) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3459 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2021) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3458 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2022) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3457 ( .A(
        oc8051_ram_top1_oc8051_idata_n2019), .B(
        oc8051_ram_top1_oc8051_idata_n2020), .C(
        oc8051_ram_top1_oc8051_idata_n2021), .D(
        oc8051_ram_top1_oc8051_idata_n2022), .Y(
        oc8051_ram_top1_oc8051_idata_n1986) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3456 ( .A(
        oc8051_ram_top1_oc8051_idata_n504), .Y(
        oc8051_ram_top1_oc8051_idata_n2016) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3455 ( .A(
        oc8051_ram_top1_oc8051_idata_n512), .Y(
        oc8051_ram_top1_oc8051_idata_n2017) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3454 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1059) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3453 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1069) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3452 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1059), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1069), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n2018) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3451 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n2016), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n2017), .C0(
        oc8051_ram_top1_oc8051_idata_n2018), .Y(
        oc8051_ram_top1_oc8051_idata_n2007) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3450 ( .A(
        oc8051_ram_top1_oc8051_idata_n488), .Y(
        oc8051_ram_top1_oc8051_idata_n2013) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3449 ( .A(
        oc8051_ram_top1_oc8051_idata_n496), .Y(
        oc8051_ram_top1_oc8051_idata_n2014) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3448 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1033) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3447 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1045) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3446 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1033), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1045), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n2015) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3445 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n2013), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n2014), .C0(
        oc8051_ram_top1_oc8051_idata_n2015), .Y(
        oc8051_ram_top1_oc8051_idata_n2008) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3444 ( .A0(
        oc8051_ram_top1_oc8051_idata_n480), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n472), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n2012) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3443 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n2012), .Y(
        oc8051_ram_top1_oc8051_idata_n2009) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3442 ( .A0(
        oc8051_ram_top1_oc8051_idata_n464), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n456), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n2011) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3441 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n2011), .Y(
        oc8051_ram_top1_oc8051_idata_n2010) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3440 ( .A(
        oc8051_ram_top1_oc8051_idata_n2007), .B(
        oc8051_ram_top1_oc8051_idata_n2008), .C(
        oc8051_ram_top1_oc8051_idata_n2009), .D(
        oc8051_ram_top1_oc8051_idata_n2010), .Y(
        oc8051_ram_top1_oc8051_idata_n1987) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3439 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2003) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3438 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2004) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3437 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2005) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3436 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2006) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3435 ( .A(
        oc8051_ram_top1_oc8051_idata_n2003), .B(
        oc8051_ram_top1_oc8051_idata_n2004), .C(
        oc8051_ram_top1_oc8051_idata_n2005), .D(
        oc8051_ram_top1_oc8051_idata_n2006), .Y(
        oc8051_ram_top1_oc8051_idata_n1988) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3434 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1999) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3433 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2000) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3432 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2001) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3431 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n2002) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3430 ( .A(
        oc8051_ram_top1_oc8051_idata_n1999), .B(
        oc8051_ram_top1_oc8051_idata_n2000), .C(
        oc8051_ram_top1_oc8051_idata_n2001), .D(
        oc8051_ram_top1_oc8051_idata_n2002), .Y(
        oc8051_ram_top1_oc8051_idata_n1989) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3429 ( .A0(
        oc8051_ram_top1_oc8051_idata_n448), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n440), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1998) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3428 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1998), .Y(
        oc8051_ram_top1_oc8051_idata_n1991) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3427 ( .A0(
        oc8051_ram_top1_oc8051_idata_n432), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n424), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1997) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3426 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1997), .Y(
        oc8051_ram_top1_oc8051_idata_n1992) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3425 ( .A0(
        oc8051_ram_top1_oc8051_idata_n416), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n408), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1996) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3424 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1996), .Y(
        oc8051_ram_top1_oc8051_idata_n1993) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3423 ( .A0(
        oc8051_ram_top1_oc8051_idata_n400), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n392), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1995) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3422 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1995), .Y(
        oc8051_ram_top1_oc8051_idata_n1994) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3421 ( .A(
        oc8051_ram_top1_oc8051_idata_n1991), .B(
        oc8051_ram_top1_oc8051_idata_n1992), .C(
        oc8051_ram_top1_oc8051_idata_n1993), .D(
        oc8051_ram_top1_oc8051_idata_n1994), .Y(
        oc8051_ram_top1_oc8051_idata_n1990) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3420 ( .A(
        oc8051_ram_top1_oc8051_idata_n1985), .B(
        oc8051_ram_top1_oc8051_idata_n1986), .C(
        oc8051_ram_top1_oc8051_idata_n1987), .D(
        oc8051_ram_top1_oc8051_idata_n1988), .E(
        oc8051_ram_top1_oc8051_idata_n1989), .F(
        oc8051_ram_top1_oc8051_idata_n1990), .Y(
        oc8051_ram_top1_oc8051_idata_n1984) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3419 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n1984), .B0(oc8051_ram_top1_rd_data_m[3]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n1853) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3418 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1980) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3417 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1981) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3416 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1982) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3415 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1983) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3414 ( .A(
        oc8051_ram_top1_oc8051_idata_n1980), .B(
        oc8051_ram_top1_oc8051_idata_n1981), .C(
        oc8051_ram_top1_oc8051_idata_n1982), .D(
        oc8051_ram_top1_oc8051_idata_n1983), .Y(
        oc8051_ram_top1_oc8051_idata_n1942) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3413 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1976) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3412 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1977) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3411 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1978) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3410 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1979) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3409 ( .A(
        oc8051_ram_top1_oc8051_idata_n1976), .B(
        oc8051_ram_top1_oc8051_idata_n1977), .C(
        oc8051_ram_top1_oc8051_idata_n1978), .D(
        oc8051_ram_top1_oc8051_idata_n1979), .Y(
        oc8051_ram_top1_oc8051_idata_n1943) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3408 ( .A(
        oc8051_ram_top1_oc8051_idata_n376), .Y(
        oc8051_ram_top1_oc8051_idata_n1973) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3407 ( .A(
        oc8051_ram_top1_oc8051_idata_n384), .Y(
        oc8051_ram_top1_oc8051_idata_n1974) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3406 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n951) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3405 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n960) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3404 ( .A0(
        oc8051_ram_top1_oc8051_idata_n951), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n960), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1975) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3403 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1973), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1974), .C0(
        oc8051_ram_top1_oc8051_idata_n1975), .Y(
        oc8051_ram_top1_oc8051_idata_n1964) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3402 ( .A(
        oc8051_ram_top1_oc8051_idata_n360), .Y(
        oc8051_ram_top1_oc8051_idata_n1970) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3401 ( .A(
        oc8051_ram_top1_oc8051_idata_n368), .Y(
        oc8051_ram_top1_oc8051_idata_n1971) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3400 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n930) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3399 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n940) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3398 ( .A0(
        oc8051_ram_top1_oc8051_idata_n930), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n940), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1972) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3397 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1970), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1971), .C0(
        oc8051_ram_top1_oc8051_idata_n1972), .Y(
        oc8051_ram_top1_oc8051_idata_n1965) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3396 ( .A0(
        oc8051_ram_top1_oc8051_idata_n352), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n344), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1969) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3395 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1969), .Y(
        oc8051_ram_top1_oc8051_idata_n1966) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3394 ( .A0(
        oc8051_ram_top1_oc8051_idata_n336), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n328), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1968) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3393 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1968), .Y(
        oc8051_ram_top1_oc8051_idata_n1967) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3392 ( .A(
        oc8051_ram_top1_oc8051_idata_n1964), .B(
        oc8051_ram_top1_oc8051_idata_n1965), .C(
        oc8051_ram_top1_oc8051_idata_n1966), .D(
        oc8051_ram_top1_oc8051_idata_n1967), .Y(
        oc8051_ram_top1_oc8051_idata_n1944) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3391 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1960) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3390 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1961) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3389 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1962) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3388 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1963) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3387 ( .A(
        oc8051_ram_top1_oc8051_idata_n1960), .B(
        oc8051_ram_top1_oc8051_idata_n1961), .C(
        oc8051_ram_top1_oc8051_idata_n1962), .D(
        oc8051_ram_top1_oc8051_idata_n1963), .Y(
        oc8051_ram_top1_oc8051_idata_n1945) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3386 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1956) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3385 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1957) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3384 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1958) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3383 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1959) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3382 ( .A(
        oc8051_ram_top1_oc8051_idata_n1956), .B(
        oc8051_ram_top1_oc8051_idata_n1957), .C(
        oc8051_ram_top1_oc8051_idata_n1958), .D(
        oc8051_ram_top1_oc8051_idata_n1959), .Y(
        oc8051_ram_top1_oc8051_idata_n1946) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3381 ( .A0(
        oc8051_ram_top1_oc8051_idata_n320), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n312), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1955) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3380 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1955), .Y(
        oc8051_ram_top1_oc8051_idata_n1948) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3379 ( .A0(
        oc8051_ram_top1_oc8051_idata_n304), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n296), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1954) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3378 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1954), .Y(
        oc8051_ram_top1_oc8051_idata_n1949) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3377 ( .A0(
        oc8051_ram_top1_oc8051_idata_n288), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n280), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1953) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3376 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1953), .Y(
        oc8051_ram_top1_oc8051_idata_n1950) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3375 ( .A0(
        oc8051_ram_top1_oc8051_idata_n272), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n264), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1952) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3374 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1952), .Y(
        oc8051_ram_top1_oc8051_idata_n1951) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3373 ( .A(
        oc8051_ram_top1_oc8051_idata_n1948), .B(
        oc8051_ram_top1_oc8051_idata_n1949), .C(
        oc8051_ram_top1_oc8051_idata_n1950), .D(
        oc8051_ram_top1_oc8051_idata_n1951), .Y(
        oc8051_ram_top1_oc8051_idata_n1947) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3372 ( .A(
        oc8051_ram_top1_oc8051_idata_n1942), .B(
        oc8051_ram_top1_oc8051_idata_n1943), .C(
        oc8051_ram_top1_oc8051_idata_n1944), .D(
        oc8051_ram_top1_oc8051_idata_n1945), .E(
        oc8051_ram_top1_oc8051_idata_n1946), .F(
        oc8051_ram_top1_oc8051_idata_n1947), .Y(
        oc8051_ram_top1_oc8051_idata_n1855) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3371 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1938) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3370 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1939) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3369 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1940) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3368 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1941) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3367 ( .A(
        oc8051_ram_top1_oc8051_idata_n1938), .B(
        oc8051_ram_top1_oc8051_idata_n1939), .C(
        oc8051_ram_top1_oc8051_idata_n1940), .D(
        oc8051_ram_top1_oc8051_idata_n1941), .Y(
        oc8051_ram_top1_oc8051_idata_n1900) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3366 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1934) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3365 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1935) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3364 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1936) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3363 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1937) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3362 ( .A(
        oc8051_ram_top1_oc8051_idata_n1934), .B(
        oc8051_ram_top1_oc8051_idata_n1935), .C(
        oc8051_ram_top1_oc8051_idata_n1936), .D(
        oc8051_ram_top1_oc8051_idata_n1937), .Y(
        oc8051_ram_top1_oc8051_idata_n1901) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3361 ( .A(
        oc8051_ram_top1_oc8051_idata_n248), .Y(
        oc8051_ram_top1_oc8051_idata_n1931) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3360 ( .A(
        oc8051_ram_top1_oc8051_idata_n256), .Y(
        oc8051_ram_top1_oc8051_idata_n1932) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3359 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n849) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3358 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n858) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3357 ( .A0(
        oc8051_ram_top1_oc8051_idata_n849), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n858), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1933) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3356 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1931), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1932), .C0(
        oc8051_ram_top1_oc8051_idata_n1933), .Y(
        oc8051_ram_top1_oc8051_idata_n1922) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3355 ( .A(
        oc8051_ram_top1_oc8051_idata_n232), .Y(
        oc8051_ram_top1_oc8051_idata_n1928) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3354 ( .A(
        oc8051_ram_top1_oc8051_idata_n240), .Y(
        oc8051_ram_top1_oc8051_idata_n1929) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3353 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n828) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3352 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n838) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3351 ( .A0(
        oc8051_ram_top1_oc8051_idata_n828), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n838), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1930) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3350 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1928), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1929), .C0(
        oc8051_ram_top1_oc8051_idata_n1930), .Y(
        oc8051_ram_top1_oc8051_idata_n1923) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3349 ( .A0(
        oc8051_ram_top1_oc8051_idata_n224), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n216), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1927) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3348 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1927), .Y(
        oc8051_ram_top1_oc8051_idata_n1924) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3347 ( .A0(
        oc8051_ram_top1_oc8051_idata_n208), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n200), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1926) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3346 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1926), .Y(
        oc8051_ram_top1_oc8051_idata_n1925) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3345 ( .A(
        oc8051_ram_top1_oc8051_idata_n1922), .B(
        oc8051_ram_top1_oc8051_idata_n1923), .C(
        oc8051_ram_top1_oc8051_idata_n1924), .D(
        oc8051_ram_top1_oc8051_idata_n1925), .Y(
        oc8051_ram_top1_oc8051_idata_n1902) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3344 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1918) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3343 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1919) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3342 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1920) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3341 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1921) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3340 ( .A(
        oc8051_ram_top1_oc8051_idata_n1918), .B(
        oc8051_ram_top1_oc8051_idata_n1919), .C(
        oc8051_ram_top1_oc8051_idata_n1920), .D(
        oc8051_ram_top1_oc8051_idata_n1921), .Y(
        oc8051_ram_top1_oc8051_idata_n1903) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3339 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1914) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3338 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1915) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3337 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1916) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3336 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1917) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3335 ( .A(
        oc8051_ram_top1_oc8051_idata_n1914), .B(
        oc8051_ram_top1_oc8051_idata_n1915), .C(
        oc8051_ram_top1_oc8051_idata_n1916), .D(
        oc8051_ram_top1_oc8051_idata_n1917), .Y(
        oc8051_ram_top1_oc8051_idata_n1904) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3334 ( .A0(
        oc8051_ram_top1_oc8051_idata_n192), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n184), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1913) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3333 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1913), .Y(
        oc8051_ram_top1_oc8051_idata_n1906) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3332 ( .A0(
        oc8051_ram_top1_oc8051_idata_n176), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n168), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1912) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3331 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1912), .Y(
        oc8051_ram_top1_oc8051_idata_n1907) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3330 ( .A0(
        oc8051_ram_top1_oc8051_idata_n160), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n152), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1911) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3329 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1911), .Y(
        oc8051_ram_top1_oc8051_idata_n1908) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3328 ( .A0(
        oc8051_ram_top1_oc8051_idata_n144), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n136), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1910) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3327 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1910), .Y(
        oc8051_ram_top1_oc8051_idata_n1909) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3326 ( .A(
        oc8051_ram_top1_oc8051_idata_n1906), .B(
        oc8051_ram_top1_oc8051_idata_n1907), .C(
        oc8051_ram_top1_oc8051_idata_n1908), .D(
        oc8051_ram_top1_oc8051_idata_n1909), .Y(
        oc8051_ram_top1_oc8051_idata_n1905) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3325 ( .A(
        oc8051_ram_top1_oc8051_idata_n1900), .B(
        oc8051_ram_top1_oc8051_idata_n1901), .C(
        oc8051_ram_top1_oc8051_idata_n1902), .D(
        oc8051_ram_top1_oc8051_idata_n1903), .E(
        oc8051_ram_top1_oc8051_idata_n1904), .F(
        oc8051_ram_top1_oc8051_idata_n1905), .Y(
        oc8051_ram_top1_oc8051_idata_n1856) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3324 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1896) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3323 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1897) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3322 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1898) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3321 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1899) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3320 ( .A(
        oc8051_ram_top1_oc8051_idata_n1896), .B(
        oc8051_ram_top1_oc8051_idata_n1897), .C(
        oc8051_ram_top1_oc8051_idata_n1898), .D(
        oc8051_ram_top1_oc8051_idata_n1899), .Y(
        oc8051_ram_top1_oc8051_idata_n1858) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3319 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1892) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3318 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1893) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3317 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1894) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3316 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1895) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3315 ( .A(
        oc8051_ram_top1_oc8051_idata_n1892), .B(
        oc8051_ram_top1_oc8051_idata_n1893), .C(
        oc8051_ram_top1_oc8051_idata_n1894), .D(
        oc8051_ram_top1_oc8051_idata_n1895), .Y(
        oc8051_ram_top1_oc8051_idata_n1859) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3314 ( .A(
        oc8051_ram_top1_oc8051_idata_n120), .Y(
        oc8051_ram_top1_oc8051_idata_n1889) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3313 ( .A(
        oc8051_ram_top1_oc8051_idata_n128), .Y(
        oc8051_ram_top1_oc8051_idata_n1890) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3312 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n746) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3311 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n755) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3310 ( .A0(
        oc8051_ram_top1_oc8051_idata_n746), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n755), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1891) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3309 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1889), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1890), .C0(
        oc8051_ram_top1_oc8051_idata_n1891), .Y(
        oc8051_ram_top1_oc8051_idata_n1880) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3308 ( .A(
        oc8051_ram_top1_oc8051_idata_n104), .Y(
        oc8051_ram_top1_oc8051_idata_n1886) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3307 ( .A(
        oc8051_ram_top1_oc8051_idata_n112), .Y(
        oc8051_ram_top1_oc8051_idata_n1887) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3306 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n725) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3305 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n735) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3304 ( .A0(
        oc8051_ram_top1_oc8051_idata_n725), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n735), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1888) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3303 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1886), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1887), .C0(
        oc8051_ram_top1_oc8051_idata_n1888), .Y(
        oc8051_ram_top1_oc8051_idata_n1881) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3302 ( .A0(
        oc8051_ram_top1_oc8051_idata_n96), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n88), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1885) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3301 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1885), .Y(
        oc8051_ram_top1_oc8051_idata_n1882) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3300 ( .A0(
        oc8051_ram_top1_oc8051_idata_n80), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n72), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1884) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3299 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1884), .Y(
        oc8051_ram_top1_oc8051_idata_n1883) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3298 ( .A(
        oc8051_ram_top1_oc8051_idata_n1880), .B(
        oc8051_ram_top1_oc8051_idata_n1881), .C(
        oc8051_ram_top1_oc8051_idata_n1882), .D(
        oc8051_ram_top1_oc8051_idata_n1883), .Y(
        oc8051_ram_top1_oc8051_idata_n1860) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3297 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1876) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3296 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1877) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3295 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1878) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3294 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1879) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3293 ( .A(
        oc8051_ram_top1_oc8051_idata_n1876), .B(
        oc8051_ram_top1_oc8051_idata_n1877), .C(
        oc8051_ram_top1_oc8051_idata_n1878), .D(
        oc8051_ram_top1_oc8051_idata_n1879), .Y(
        oc8051_ram_top1_oc8051_idata_n1861) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3292 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1872) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3291 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1873) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3290 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1874) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3289 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1875) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3288 ( .A(
        oc8051_ram_top1_oc8051_idata_n1872), .B(
        oc8051_ram_top1_oc8051_idata_n1873), .C(
        oc8051_ram_top1_oc8051_idata_n1874), .D(
        oc8051_ram_top1_oc8051_idata_n1875), .Y(
        oc8051_ram_top1_oc8051_idata_n1862) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3287 ( .A0(
        oc8051_ram_top1_oc8051_idata_n64), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n56), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1871) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3286 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1871), .Y(
        oc8051_ram_top1_oc8051_idata_n1864) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3285 ( .A0(
        oc8051_ram_top1_oc8051_idata_n48), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n40), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1870) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3284 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1870), .Y(
        oc8051_ram_top1_oc8051_idata_n1865) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3283 ( .A0(
        oc8051_ram_top1_oc8051_idata_n32), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n24), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1869) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3282 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1869), .Y(
        oc8051_ram_top1_oc8051_idata_n1866) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3281 ( .A0(
        oc8051_ram_top1_oc8051_idata_n16), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n8), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1868) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3280 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__3_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__3_), .C0(
        oc8051_ram_top1_oc8051_idata_n1868), .Y(
        oc8051_ram_top1_oc8051_idata_n1867) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3279 ( .A(
        oc8051_ram_top1_oc8051_idata_n1864), .B(
        oc8051_ram_top1_oc8051_idata_n1865), .C(
        oc8051_ram_top1_oc8051_idata_n1866), .D(
        oc8051_ram_top1_oc8051_idata_n1867), .Y(
        oc8051_ram_top1_oc8051_idata_n1863) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3278 ( .A(
        oc8051_ram_top1_oc8051_idata_n1858), .B(
        oc8051_ram_top1_oc8051_idata_n1859), .C(
        oc8051_ram_top1_oc8051_idata_n1860), .D(
        oc8051_ram_top1_oc8051_idata_n1861), .E(
        oc8051_ram_top1_oc8051_idata_n1862), .F(
        oc8051_ram_top1_oc8051_idata_n1863), .Y(
        oc8051_ram_top1_oc8051_idata_n1857) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3277 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n1855), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n1856), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n1857), .Y(
        oc8051_ram_top1_oc8051_idata_n1854) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3276 ( .A0(
        oc8051_ram_top1_oc8051_idata_n579), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n1853), .C0(
        oc8051_ram_top1_oc8051_idata_n1854), .Y(
        oc8051_ram_top1_oc8051_idata_n2478) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3275 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1849) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3274 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1850) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3273 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1851) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3272 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1852) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3271 ( .A(
        oc8051_ram_top1_oc8051_idata_n1849), .B(
        oc8051_ram_top1_oc8051_idata_n1850), .C(
        oc8051_ram_top1_oc8051_idata_n1851), .D(
        oc8051_ram_top1_oc8051_idata_n1852), .Y(
        oc8051_ram_top1_oc8051_idata_n1811) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3270 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1845) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3269 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1846) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3268 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1847) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3267 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1848) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3266 ( .A(
        oc8051_ram_top1_oc8051_idata_n1845), .B(
        oc8051_ram_top1_oc8051_idata_n1846), .C(
        oc8051_ram_top1_oc8051_idata_n1847), .D(
        oc8051_ram_top1_oc8051_idata_n1848), .Y(
        oc8051_ram_top1_oc8051_idata_n1812) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3265 ( .A(
        oc8051_ram_top1_oc8051_idata_n503), .Y(
        oc8051_ram_top1_oc8051_idata_n1842) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3264 ( .A(
        oc8051_ram_top1_oc8051_idata_n511), .Y(
        oc8051_ram_top1_oc8051_idata_n1843) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3263 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1058) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3262 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1068) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3261 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1058), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1068), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1844) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3260 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1842), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1843), .C0(
        oc8051_ram_top1_oc8051_idata_n1844), .Y(
        oc8051_ram_top1_oc8051_idata_n1833) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3259 ( .A(
        oc8051_ram_top1_oc8051_idata_n487), .Y(
        oc8051_ram_top1_oc8051_idata_n1839) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3258 ( .A(
        oc8051_ram_top1_oc8051_idata_n495), .Y(
        oc8051_ram_top1_oc8051_idata_n1840) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3257 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1032) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3256 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1044) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3255 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1032), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1044), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1841) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3254 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1839), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1840), .C0(
        oc8051_ram_top1_oc8051_idata_n1841), .Y(
        oc8051_ram_top1_oc8051_idata_n1834) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3253 ( .A0(
        oc8051_ram_top1_oc8051_idata_n479), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n471), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1838) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3252 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1838), .Y(
        oc8051_ram_top1_oc8051_idata_n1835) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3251 ( .A0(
        oc8051_ram_top1_oc8051_idata_n463), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n455), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1837) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3250 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1837), .Y(
        oc8051_ram_top1_oc8051_idata_n1836) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3249 ( .A(
        oc8051_ram_top1_oc8051_idata_n1833), .B(
        oc8051_ram_top1_oc8051_idata_n1834), .C(
        oc8051_ram_top1_oc8051_idata_n1835), .D(
        oc8051_ram_top1_oc8051_idata_n1836), .Y(
        oc8051_ram_top1_oc8051_idata_n1813) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3248 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1829) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3247 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1830) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3246 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1831) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3245 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1832) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3244 ( .A(
        oc8051_ram_top1_oc8051_idata_n1829), .B(
        oc8051_ram_top1_oc8051_idata_n1830), .C(
        oc8051_ram_top1_oc8051_idata_n1831), .D(
        oc8051_ram_top1_oc8051_idata_n1832), .Y(
        oc8051_ram_top1_oc8051_idata_n1814) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3243 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1825) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3242 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1826) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3241 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1827) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3240 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1828) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3239 ( .A(
        oc8051_ram_top1_oc8051_idata_n1825), .B(
        oc8051_ram_top1_oc8051_idata_n1826), .C(
        oc8051_ram_top1_oc8051_idata_n1827), .D(
        oc8051_ram_top1_oc8051_idata_n1828), .Y(
        oc8051_ram_top1_oc8051_idata_n1815) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3238 ( .A0(
        oc8051_ram_top1_oc8051_idata_n447), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n439), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1824) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3237 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1824), .Y(
        oc8051_ram_top1_oc8051_idata_n1817) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3236 ( .A0(
        oc8051_ram_top1_oc8051_idata_n431), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n423), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1823) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3235 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1823), .Y(
        oc8051_ram_top1_oc8051_idata_n1818) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3234 ( .A0(
        oc8051_ram_top1_oc8051_idata_n415), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n407), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1822) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3233 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1822), .Y(
        oc8051_ram_top1_oc8051_idata_n1819) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3232 ( .A0(
        oc8051_ram_top1_oc8051_idata_n399), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n391), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1821) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3231 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1821), .Y(
        oc8051_ram_top1_oc8051_idata_n1820) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3230 ( .A(
        oc8051_ram_top1_oc8051_idata_n1817), .B(
        oc8051_ram_top1_oc8051_idata_n1818), .C(
        oc8051_ram_top1_oc8051_idata_n1819), .D(
        oc8051_ram_top1_oc8051_idata_n1820), .Y(
        oc8051_ram_top1_oc8051_idata_n1816) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3229 ( .A(
        oc8051_ram_top1_oc8051_idata_n1811), .B(
        oc8051_ram_top1_oc8051_idata_n1812), .C(
        oc8051_ram_top1_oc8051_idata_n1813), .D(
        oc8051_ram_top1_oc8051_idata_n1814), .E(
        oc8051_ram_top1_oc8051_idata_n1815), .F(
        oc8051_ram_top1_oc8051_idata_n1816), .Y(
        oc8051_ram_top1_oc8051_idata_n1810) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3228 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n1810), .B0(oc8051_ram_top1_rd_data_m[4]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n1679) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3227 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1806) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3226 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1807) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3225 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1808) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3224 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1809) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3223 ( .A(
        oc8051_ram_top1_oc8051_idata_n1806), .B(
        oc8051_ram_top1_oc8051_idata_n1807), .C(
        oc8051_ram_top1_oc8051_idata_n1808), .D(
        oc8051_ram_top1_oc8051_idata_n1809), .Y(
        oc8051_ram_top1_oc8051_idata_n1768) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3222 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1802) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3221 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1803) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3220 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1804) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3219 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1805) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3218 ( .A(
        oc8051_ram_top1_oc8051_idata_n1802), .B(
        oc8051_ram_top1_oc8051_idata_n1803), .C(
        oc8051_ram_top1_oc8051_idata_n1804), .D(
        oc8051_ram_top1_oc8051_idata_n1805), .Y(
        oc8051_ram_top1_oc8051_idata_n1769) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3217 ( .A(
        oc8051_ram_top1_oc8051_idata_n375), .Y(
        oc8051_ram_top1_oc8051_idata_n1799) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3216 ( .A(
        oc8051_ram_top1_oc8051_idata_n383), .Y(
        oc8051_ram_top1_oc8051_idata_n1800) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3215 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n950) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3214 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n959) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3213 ( .A0(
        oc8051_ram_top1_oc8051_idata_n950), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n959), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1801) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3212 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1799), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1800), .C0(
        oc8051_ram_top1_oc8051_idata_n1801), .Y(
        oc8051_ram_top1_oc8051_idata_n1790) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3211 ( .A(
        oc8051_ram_top1_oc8051_idata_n359), .Y(
        oc8051_ram_top1_oc8051_idata_n1796) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3210 ( .A(
        oc8051_ram_top1_oc8051_idata_n367), .Y(
        oc8051_ram_top1_oc8051_idata_n1797) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3209 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n929) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3208 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n939) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3207 ( .A0(
        oc8051_ram_top1_oc8051_idata_n929), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n939), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1798) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3206 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1796), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1797), .C0(
        oc8051_ram_top1_oc8051_idata_n1798), .Y(
        oc8051_ram_top1_oc8051_idata_n1791) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3205 ( .A0(
        oc8051_ram_top1_oc8051_idata_n351), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n343), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1795) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3204 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1795), .Y(
        oc8051_ram_top1_oc8051_idata_n1792) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3203 ( .A0(
        oc8051_ram_top1_oc8051_idata_n335), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n327), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1794) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3202 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1794), .Y(
        oc8051_ram_top1_oc8051_idata_n1793) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3201 ( .A(
        oc8051_ram_top1_oc8051_idata_n1790), .B(
        oc8051_ram_top1_oc8051_idata_n1791), .C(
        oc8051_ram_top1_oc8051_idata_n1792), .D(
        oc8051_ram_top1_oc8051_idata_n1793), .Y(
        oc8051_ram_top1_oc8051_idata_n1770) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3200 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1786) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3199 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1787) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3198 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1788) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3197 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1789) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3196 ( .A(
        oc8051_ram_top1_oc8051_idata_n1786), .B(
        oc8051_ram_top1_oc8051_idata_n1787), .C(
        oc8051_ram_top1_oc8051_idata_n1788), .D(
        oc8051_ram_top1_oc8051_idata_n1789), .Y(
        oc8051_ram_top1_oc8051_idata_n1771) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3195 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1782) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3194 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1783) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3193 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1784) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3192 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1785) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3191 ( .A(
        oc8051_ram_top1_oc8051_idata_n1782), .B(
        oc8051_ram_top1_oc8051_idata_n1783), .C(
        oc8051_ram_top1_oc8051_idata_n1784), .D(
        oc8051_ram_top1_oc8051_idata_n1785), .Y(
        oc8051_ram_top1_oc8051_idata_n1772) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3190 ( .A0(
        oc8051_ram_top1_oc8051_idata_n319), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n311), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1781) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3189 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1781), .Y(
        oc8051_ram_top1_oc8051_idata_n1774) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3188 ( .A0(
        oc8051_ram_top1_oc8051_idata_n303), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n295), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1780) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3187 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1780), .Y(
        oc8051_ram_top1_oc8051_idata_n1775) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3186 ( .A0(
        oc8051_ram_top1_oc8051_idata_n287), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n279), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1779) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3185 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1779), .Y(
        oc8051_ram_top1_oc8051_idata_n1776) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3184 ( .A0(
        oc8051_ram_top1_oc8051_idata_n271), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n263), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1778) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3183 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1778), .Y(
        oc8051_ram_top1_oc8051_idata_n1777) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3182 ( .A(
        oc8051_ram_top1_oc8051_idata_n1774), .B(
        oc8051_ram_top1_oc8051_idata_n1775), .C(
        oc8051_ram_top1_oc8051_idata_n1776), .D(
        oc8051_ram_top1_oc8051_idata_n1777), .Y(
        oc8051_ram_top1_oc8051_idata_n1773) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3181 ( .A(
        oc8051_ram_top1_oc8051_idata_n1768), .B(
        oc8051_ram_top1_oc8051_idata_n1769), .C(
        oc8051_ram_top1_oc8051_idata_n1770), .D(
        oc8051_ram_top1_oc8051_idata_n1771), .E(
        oc8051_ram_top1_oc8051_idata_n1772), .F(
        oc8051_ram_top1_oc8051_idata_n1773), .Y(
        oc8051_ram_top1_oc8051_idata_n1681) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3180 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1764) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3179 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1765) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3178 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1766) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3177 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1767) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3176 ( .A(
        oc8051_ram_top1_oc8051_idata_n1764), .B(
        oc8051_ram_top1_oc8051_idata_n1765), .C(
        oc8051_ram_top1_oc8051_idata_n1766), .D(
        oc8051_ram_top1_oc8051_idata_n1767), .Y(
        oc8051_ram_top1_oc8051_idata_n1726) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3175 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1760) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3174 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1761) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3173 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1762) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3172 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1763) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3171 ( .A(
        oc8051_ram_top1_oc8051_idata_n1760), .B(
        oc8051_ram_top1_oc8051_idata_n1761), .C(
        oc8051_ram_top1_oc8051_idata_n1762), .D(
        oc8051_ram_top1_oc8051_idata_n1763), .Y(
        oc8051_ram_top1_oc8051_idata_n1727) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3170 ( .A(
        oc8051_ram_top1_oc8051_idata_n247), .Y(
        oc8051_ram_top1_oc8051_idata_n1757) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3169 ( .A(
        oc8051_ram_top1_oc8051_idata_n255), .Y(
        oc8051_ram_top1_oc8051_idata_n1758) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3168 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n848) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3167 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n857) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3166 ( .A0(
        oc8051_ram_top1_oc8051_idata_n848), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n857), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1759) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3165 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1757), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1758), .C0(
        oc8051_ram_top1_oc8051_idata_n1759), .Y(
        oc8051_ram_top1_oc8051_idata_n1748) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3164 ( .A(
        oc8051_ram_top1_oc8051_idata_n231), .Y(
        oc8051_ram_top1_oc8051_idata_n1754) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3163 ( .A(
        oc8051_ram_top1_oc8051_idata_n239), .Y(
        oc8051_ram_top1_oc8051_idata_n1755) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3162 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n827) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3161 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n837) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3160 ( .A0(
        oc8051_ram_top1_oc8051_idata_n827), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n837), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1756) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3159 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1754), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1755), .C0(
        oc8051_ram_top1_oc8051_idata_n1756), .Y(
        oc8051_ram_top1_oc8051_idata_n1749) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3158 ( .A0(
        oc8051_ram_top1_oc8051_idata_n223), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n215), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1753) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3157 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1753), .Y(
        oc8051_ram_top1_oc8051_idata_n1750) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3156 ( .A0(
        oc8051_ram_top1_oc8051_idata_n207), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n199), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1752) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3155 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1752), .Y(
        oc8051_ram_top1_oc8051_idata_n1751) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3154 ( .A(
        oc8051_ram_top1_oc8051_idata_n1748), .B(
        oc8051_ram_top1_oc8051_idata_n1749), .C(
        oc8051_ram_top1_oc8051_idata_n1750), .D(
        oc8051_ram_top1_oc8051_idata_n1751), .Y(
        oc8051_ram_top1_oc8051_idata_n1728) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3153 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1744) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3152 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1745) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3151 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1746) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3150 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1747) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3149 ( .A(
        oc8051_ram_top1_oc8051_idata_n1744), .B(
        oc8051_ram_top1_oc8051_idata_n1745), .C(
        oc8051_ram_top1_oc8051_idata_n1746), .D(
        oc8051_ram_top1_oc8051_idata_n1747), .Y(
        oc8051_ram_top1_oc8051_idata_n1729) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3148 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1740) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3147 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1741) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3146 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1742) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3145 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1743) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3144 ( .A(
        oc8051_ram_top1_oc8051_idata_n1740), .B(
        oc8051_ram_top1_oc8051_idata_n1741), .C(
        oc8051_ram_top1_oc8051_idata_n1742), .D(
        oc8051_ram_top1_oc8051_idata_n1743), .Y(
        oc8051_ram_top1_oc8051_idata_n1730) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3143 ( .A0(
        oc8051_ram_top1_oc8051_idata_n191), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n183), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1739) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3142 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1739), .Y(
        oc8051_ram_top1_oc8051_idata_n1732) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3141 ( .A0(
        oc8051_ram_top1_oc8051_idata_n175), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n167), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1738) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3140 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1738), .Y(
        oc8051_ram_top1_oc8051_idata_n1733) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3139 ( .A0(
        oc8051_ram_top1_oc8051_idata_n159), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n151), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1737) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3138 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1737), .Y(
        oc8051_ram_top1_oc8051_idata_n1734) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3137 ( .A0(
        oc8051_ram_top1_oc8051_idata_n143), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n135), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1736) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3136 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1736), .Y(
        oc8051_ram_top1_oc8051_idata_n1735) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3135 ( .A(
        oc8051_ram_top1_oc8051_idata_n1732), .B(
        oc8051_ram_top1_oc8051_idata_n1733), .C(
        oc8051_ram_top1_oc8051_idata_n1734), .D(
        oc8051_ram_top1_oc8051_idata_n1735), .Y(
        oc8051_ram_top1_oc8051_idata_n1731) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3134 ( .A(
        oc8051_ram_top1_oc8051_idata_n1726), .B(
        oc8051_ram_top1_oc8051_idata_n1727), .C(
        oc8051_ram_top1_oc8051_idata_n1728), .D(
        oc8051_ram_top1_oc8051_idata_n1729), .E(
        oc8051_ram_top1_oc8051_idata_n1730), .F(
        oc8051_ram_top1_oc8051_idata_n1731), .Y(
        oc8051_ram_top1_oc8051_idata_n1682) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3133 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1722) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3132 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1723) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3131 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1724) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3130 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1725) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3129 ( .A(
        oc8051_ram_top1_oc8051_idata_n1722), .B(
        oc8051_ram_top1_oc8051_idata_n1723), .C(
        oc8051_ram_top1_oc8051_idata_n1724), .D(
        oc8051_ram_top1_oc8051_idata_n1725), .Y(
        oc8051_ram_top1_oc8051_idata_n1684) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3128 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1718) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3127 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1719) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3126 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1720) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3125 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1721) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3124 ( .A(
        oc8051_ram_top1_oc8051_idata_n1718), .B(
        oc8051_ram_top1_oc8051_idata_n1719), .C(
        oc8051_ram_top1_oc8051_idata_n1720), .D(
        oc8051_ram_top1_oc8051_idata_n1721), .Y(
        oc8051_ram_top1_oc8051_idata_n1685) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3123 ( .A(
        oc8051_ram_top1_oc8051_idata_n119), .Y(
        oc8051_ram_top1_oc8051_idata_n1715) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3122 ( .A(
        oc8051_ram_top1_oc8051_idata_n127), .Y(
        oc8051_ram_top1_oc8051_idata_n1716) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3121 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n745) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3120 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n754) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3119 ( .A0(
        oc8051_ram_top1_oc8051_idata_n745), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n754), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1717) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3118 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1715), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1716), .C0(
        oc8051_ram_top1_oc8051_idata_n1717), .Y(
        oc8051_ram_top1_oc8051_idata_n1706) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3117 ( .A(
        oc8051_ram_top1_oc8051_idata_n103), .Y(
        oc8051_ram_top1_oc8051_idata_n1712) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3116 ( .A(
        oc8051_ram_top1_oc8051_idata_n111), .Y(
        oc8051_ram_top1_oc8051_idata_n1713) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3115 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n724) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3114 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n734) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3113 ( .A0(
        oc8051_ram_top1_oc8051_idata_n724), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n734), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1714) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3112 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1712), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1713), .C0(
        oc8051_ram_top1_oc8051_idata_n1714), .Y(
        oc8051_ram_top1_oc8051_idata_n1707) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3111 ( .A0(
        oc8051_ram_top1_oc8051_idata_n95), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n87), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1711) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3110 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1711), .Y(
        oc8051_ram_top1_oc8051_idata_n1708) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3109 ( .A0(
        oc8051_ram_top1_oc8051_idata_n79), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n71), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1710) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3108 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1710), .Y(
        oc8051_ram_top1_oc8051_idata_n1709) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3107 ( .A(
        oc8051_ram_top1_oc8051_idata_n1706), .B(
        oc8051_ram_top1_oc8051_idata_n1707), .C(
        oc8051_ram_top1_oc8051_idata_n1708), .D(
        oc8051_ram_top1_oc8051_idata_n1709), .Y(
        oc8051_ram_top1_oc8051_idata_n1686) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3106 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1702) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3105 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1703) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3104 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1704) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3103 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1705) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3102 ( .A(
        oc8051_ram_top1_oc8051_idata_n1702), .B(
        oc8051_ram_top1_oc8051_idata_n1703), .C(
        oc8051_ram_top1_oc8051_idata_n1704), .D(
        oc8051_ram_top1_oc8051_idata_n1705), .Y(
        oc8051_ram_top1_oc8051_idata_n1687) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3101 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1698) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3100 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1699) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3099 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1700) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3098 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__4_), .Y(
        oc8051_ram_top1_oc8051_idata_n1701) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3097 ( .A(
        oc8051_ram_top1_oc8051_idata_n1698), .B(
        oc8051_ram_top1_oc8051_idata_n1699), .C(
        oc8051_ram_top1_oc8051_idata_n1700), .D(
        oc8051_ram_top1_oc8051_idata_n1701), .Y(
        oc8051_ram_top1_oc8051_idata_n1688) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3096 ( .A0(
        oc8051_ram_top1_oc8051_idata_n63), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n55), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1697) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3095 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1697), .Y(
        oc8051_ram_top1_oc8051_idata_n1690) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3094 ( .A0(
        oc8051_ram_top1_oc8051_idata_n47), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n39), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1696) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3093 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1696), .Y(
        oc8051_ram_top1_oc8051_idata_n1691) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3092 ( .A0(
        oc8051_ram_top1_oc8051_idata_n31), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n23), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1695) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3091 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1695), .Y(
        oc8051_ram_top1_oc8051_idata_n1692) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3090 ( .A0(
        oc8051_ram_top1_oc8051_idata_n15), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n7), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1694) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3089 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__4_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__4_), .C0(
        oc8051_ram_top1_oc8051_idata_n1694), .Y(
        oc8051_ram_top1_oc8051_idata_n1693) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3088 ( .A(
        oc8051_ram_top1_oc8051_idata_n1690), .B(
        oc8051_ram_top1_oc8051_idata_n1691), .C(
        oc8051_ram_top1_oc8051_idata_n1692), .D(
        oc8051_ram_top1_oc8051_idata_n1693), .Y(
        oc8051_ram_top1_oc8051_idata_n1689) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3087 ( .A(
        oc8051_ram_top1_oc8051_idata_n1684), .B(
        oc8051_ram_top1_oc8051_idata_n1685), .C(
        oc8051_ram_top1_oc8051_idata_n1686), .D(
        oc8051_ram_top1_oc8051_idata_n1687), .E(
        oc8051_ram_top1_oc8051_idata_n1688), .F(
        oc8051_ram_top1_oc8051_idata_n1689), .Y(
        oc8051_ram_top1_oc8051_idata_n1683) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3086 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n1681), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n1682), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n1683), .Y(
        oc8051_ram_top1_oc8051_idata_n1680) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3085 ( .A0(
        oc8051_ram_top1_oc8051_idata_n596), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n1679), .C0(
        oc8051_ram_top1_oc8051_idata_n1680), .Y(
        oc8051_ram_top1_oc8051_idata_n2479) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3084 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1675) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3083 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1676) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3082 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1677) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3081 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1678) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3080 ( .A(
        oc8051_ram_top1_oc8051_idata_n1675), .B(
        oc8051_ram_top1_oc8051_idata_n1676), .C(
        oc8051_ram_top1_oc8051_idata_n1677), .D(
        oc8051_ram_top1_oc8051_idata_n1678), .Y(
        oc8051_ram_top1_oc8051_idata_n1637) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3079 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1671) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3078 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1672) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3077 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1673) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3076 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1674) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3075 ( .A(
        oc8051_ram_top1_oc8051_idata_n1671), .B(
        oc8051_ram_top1_oc8051_idata_n1672), .C(
        oc8051_ram_top1_oc8051_idata_n1673), .D(
        oc8051_ram_top1_oc8051_idata_n1674), .Y(
        oc8051_ram_top1_oc8051_idata_n1638) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3074 ( .A(
        oc8051_ram_top1_oc8051_idata_n502), .Y(
        oc8051_ram_top1_oc8051_idata_n1668) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3073 ( .A(
        oc8051_ram_top1_oc8051_idata_n510), .Y(
        oc8051_ram_top1_oc8051_idata_n1669) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3072 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1057) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3071 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1067) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3070 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1057), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1067), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1670) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3069 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1668), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1669), .C0(
        oc8051_ram_top1_oc8051_idata_n1670), .Y(
        oc8051_ram_top1_oc8051_idata_n1659) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3068 ( .A(
        oc8051_ram_top1_oc8051_idata_n486), .Y(
        oc8051_ram_top1_oc8051_idata_n1665) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3067 ( .A(
        oc8051_ram_top1_oc8051_idata_n494), .Y(
        oc8051_ram_top1_oc8051_idata_n1666) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3066 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1031) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3065 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1043) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3064 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1031), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1043), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1667) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3063 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1665), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1666), .C0(
        oc8051_ram_top1_oc8051_idata_n1667), .Y(
        oc8051_ram_top1_oc8051_idata_n1660) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3062 ( .A0(
        oc8051_ram_top1_oc8051_idata_n478), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n470), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1664) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3061 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1664), .Y(
        oc8051_ram_top1_oc8051_idata_n1661) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3060 ( .A0(
        oc8051_ram_top1_oc8051_idata_n462), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n454), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1663) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3059 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1663), .Y(
        oc8051_ram_top1_oc8051_idata_n1662) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3058 ( .A(
        oc8051_ram_top1_oc8051_idata_n1659), .B(
        oc8051_ram_top1_oc8051_idata_n1660), .C(
        oc8051_ram_top1_oc8051_idata_n1661), .D(
        oc8051_ram_top1_oc8051_idata_n1662), .Y(
        oc8051_ram_top1_oc8051_idata_n1639) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3057 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1655) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3056 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1656) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3055 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1657) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3054 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1658) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3053 ( .A(
        oc8051_ram_top1_oc8051_idata_n1655), .B(
        oc8051_ram_top1_oc8051_idata_n1656), .C(
        oc8051_ram_top1_oc8051_idata_n1657), .D(
        oc8051_ram_top1_oc8051_idata_n1658), .Y(
        oc8051_ram_top1_oc8051_idata_n1640) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3052 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1651) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3051 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1652) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3050 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1653) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3049 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1654) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3048 ( .A(
        oc8051_ram_top1_oc8051_idata_n1651), .B(
        oc8051_ram_top1_oc8051_idata_n1652), .C(
        oc8051_ram_top1_oc8051_idata_n1653), .D(
        oc8051_ram_top1_oc8051_idata_n1654), .Y(
        oc8051_ram_top1_oc8051_idata_n1641) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3047 ( .A0(
        oc8051_ram_top1_oc8051_idata_n446), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n438), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1650) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3046 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1650), .Y(
        oc8051_ram_top1_oc8051_idata_n1643) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3045 ( .A0(
        oc8051_ram_top1_oc8051_idata_n430), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n422), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1649) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3044 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1649), .Y(
        oc8051_ram_top1_oc8051_idata_n1644) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3043 ( .A0(
        oc8051_ram_top1_oc8051_idata_n414), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n406), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1648) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3042 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1648), .Y(
        oc8051_ram_top1_oc8051_idata_n1645) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3041 ( .A0(
        oc8051_ram_top1_oc8051_idata_n398), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n390), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1647) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3040 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1647), .Y(
        oc8051_ram_top1_oc8051_idata_n1646) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3039 ( .A(
        oc8051_ram_top1_oc8051_idata_n1643), .B(
        oc8051_ram_top1_oc8051_idata_n1644), .C(
        oc8051_ram_top1_oc8051_idata_n1645), .D(
        oc8051_ram_top1_oc8051_idata_n1646), .Y(
        oc8051_ram_top1_oc8051_idata_n1642) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3038 ( .A(
        oc8051_ram_top1_oc8051_idata_n1637), .B(
        oc8051_ram_top1_oc8051_idata_n1638), .C(
        oc8051_ram_top1_oc8051_idata_n1639), .D(
        oc8051_ram_top1_oc8051_idata_n1640), .E(
        oc8051_ram_top1_oc8051_idata_n1641), .F(
        oc8051_ram_top1_oc8051_idata_n1642), .Y(
        oc8051_ram_top1_oc8051_idata_n1636) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3037 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n1636), .B0(oc8051_ram_top1_rd_data_m[5]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n1505) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3036 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1632) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3035 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1633) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3034 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1634) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3033 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1635) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3032 ( .A(
        oc8051_ram_top1_oc8051_idata_n1632), .B(
        oc8051_ram_top1_oc8051_idata_n1633), .C(
        oc8051_ram_top1_oc8051_idata_n1634), .D(
        oc8051_ram_top1_oc8051_idata_n1635), .Y(
        oc8051_ram_top1_oc8051_idata_n1594) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3031 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1628) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3030 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1629) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3029 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1630) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3028 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1631) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3027 ( .A(
        oc8051_ram_top1_oc8051_idata_n1628), .B(
        oc8051_ram_top1_oc8051_idata_n1629), .C(
        oc8051_ram_top1_oc8051_idata_n1630), .D(
        oc8051_ram_top1_oc8051_idata_n1631), .Y(
        oc8051_ram_top1_oc8051_idata_n1595) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3026 ( .A(
        oc8051_ram_top1_oc8051_idata_n374), .Y(
        oc8051_ram_top1_oc8051_idata_n1625) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3025 ( .A(
        oc8051_ram_top1_oc8051_idata_n382), .Y(
        oc8051_ram_top1_oc8051_idata_n1626) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3024 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n949) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3023 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n958) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3022 ( .A0(
        oc8051_ram_top1_oc8051_idata_n949), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n958), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1627) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3021 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1625), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1626), .C0(
        oc8051_ram_top1_oc8051_idata_n1627), .Y(
        oc8051_ram_top1_oc8051_idata_n1616) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3020 ( .A(
        oc8051_ram_top1_oc8051_idata_n358), .Y(
        oc8051_ram_top1_oc8051_idata_n1622) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3019 ( .A(
        oc8051_ram_top1_oc8051_idata_n366), .Y(
        oc8051_ram_top1_oc8051_idata_n1623) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3018 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n928) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u3017 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n938) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3016 ( .A0(
        oc8051_ram_top1_oc8051_idata_n928), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n938), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1624) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3015 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1622), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1623), .C0(
        oc8051_ram_top1_oc8051_idata_n1624), .Y(
        oc8051_ram_top1_oc8051_idata_n1617) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3014 ( .A0(
        oc8051_ram_top1_oc8051_idata_n350), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n342), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1621) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3013 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1621), .Y(
        oc8051_ram_top1_oc8051_idata_n1618) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3012 ( .A0(
        oc8051_ram_top1_oc8051_idata_n334), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n326), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1620) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3011 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1620), .Y(
        oc8051_ram_top1_oc8051_idata_n1619) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3010 ( .A(
        oc8051_ram_top1_oc8051_idata_n1616), .B(
        oc8051_ram_top1_oc8051_idata_n1617), .C(
        oc8051_ram_top1_oc8051_idata_n1618), .D(
        oc8051_ram_top1_oc8051_idata_n1619), .Y(
        oc8051_ram_top1_oc8051_idata_n1596) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3009 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1612) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3008 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1613) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3007 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1614) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3006 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1615) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3005 ( .A(
        oc8051_ram_top1_oc8051_idata_n1612), .B(
        oc8051_ram_top1_oc8051_idata_n1613), .C(
        oc8051_ram_top1_oc8051_idata_n1614), .D(
        oc8051_ram_top1_oc8051_idata_n1615), .Y(
        oc8051_ram_top1_oc8051_idata_n1597) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3004 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1608) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3003 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1609) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3002 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1610) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u3001 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1611) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u3000 ( .A(
        oc8051_ram_top1_oc8051_idata_n1608), .B(
        oc8051_ram_top1_oc8051_idata_n1609), .C(
        oc8051_ram_top1_oc8051_idata_n1610), .D(
        oc8051_ram_top1_oc8051_idata_n1611), .Y(
        oc8051_ram_top1_oc8051_idata_n1598) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2999 ( .A0(
        oc8051_ram_top1_oc8051_idata_n318), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n310), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1607) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2998 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1607), .Y(
        oc8051_ram_top1_oc8051_idata_n1600) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2997 ( .A0(
        oc8051_ram_top1_oc8051_idata_n302), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n294), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1606) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2996 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1606), .Y(
        oc8051_ram_top1_oc8051_idata_n1601) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2995 ( .A0(
        oc8051_ram_top1_oc8051_idata_n286), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n278), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1605) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2994 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1605), .Y(
        oc8051_ram_top1_oc8051_idata_n1602) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2993 ( .A0(
        oc8051_ram_top1_oc8051_idata_n270), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n262), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1604) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2992 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1604), .Y(
        oc8051_ram_top1_oc8051_idata_n1603) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2991 ( .A(
        oc8051_ram_top1_oc8051_idata_n1600), .B(
        oc8051_ram_top1_oc8051_idata_n1601), .C(
        oc8051_ram_top1_oc8051_idata_n1602), .D(
        oc8051_ram_top1_oc8051_idata_n1603), .Y(
        oc8051_ram_top1_oc8051_idata_n1599) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2990 ( .A(
        oc8051_ram_top1_oc8051_idata_n1594), .B(
        oc8051_ram_top1_oc8051_idata_n1595), .C(
        oc8051_ram_top1_oc8051_idata_n1596), .D(
        oc8051_ram_top1_oc8051_idata_n1597), .E(
        oc8051_ram_top1_oc8051_idata_n1598), .F(
        oc8051_ram_top1_oc8051_idata_n1599), .Y(
        oc8051_ram_top1_oc8051_idata_n1507) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2989 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1590) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2988 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1591) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2987 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1592) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2986 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1593) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2985 ( .A(
        oc8051_ram_top1_oc8051_idata_n1590), .B(
        oc8051_ram_top1_oc8051_idata_n1591), .C(
        oc8051_ram_top1_oc8051_idata_n1592), .D(
        oc8051_ram_top1_oc8051_idata_n1593), .Y(
        oc8051_ram_top1_oc8051_idata_n1552) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2984 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1586) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2983 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1587) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2982 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1588) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2981 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1589) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2980 ( .A(
        oc8051_ram_top1_oc8051_idata_n1586), .B(
        oc8051_ram_top1_oc8051_idata_n1587), .C(
        oc8051_ram_top1_oc8051_idata_n1588), .D(
        oc8051_ram_top1_oc8051_idata_n1589), .Y(
        oc8051_ram_top1_oc8051_idata_n1553) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2979 ( .A(
        oc8051_ram_top1_oc8051_idata_n246), .Y(
        oc8051_ram_top1_oc8051_idata_n1583) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2978 ( .A(
        oc8051_ram_top1_oc8051_idata_n254), .Y(
        oc8051_ram_top1_oc8051_idata_n1584) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2977 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n847) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2976 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n856) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2975 ( .A0(
        oc8051_ram_top1_oc8051_idata_n847), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n856), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1585) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2974 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1583), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1584), .C0(
        oc8051_ram_top1_oc8051_idata_n1585), .Y(
        oc8051_ram_top1_oc8051_idata_n1574) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2973 ( .A(
        oc8051_ram_top1_oc8051_idata_n230), .Y(
        oc8051_ram_top1_oc8051_idata_n1580) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2972 ( .A(
        oc8051_ram_top1_oc8051_idata_n238), .Y(
        oc8051_ram_top1_oc8051_idata_n1581) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2971 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n826) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2970 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n836) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2969 ( .A0(
        oc8051_ram_top1_oc8051_idata_n826), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n836), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1582) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2968 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1580), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1581), .C0(
        oc8051_ram_top1_oc8051_idata_n1582), .Y(
        oc8051_ram_top1_oc8051_idata_n1575) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2967 ( .A0(
        oc8051_ram_top1_oc8051_idata_n222), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n214), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1579) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2966 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1579), .Y(
        oc8051_ram_top1_oc8051_idata_n1576) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2965 ( .A0(
        oc8051_ram_top1_oc8051_idata_n206), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n198), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1578) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2964 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1578), .Y(
        oc8051_ram_top1_oc8051_idata_n1577) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2963 ( .A(
        oc8051_ram_top1_oc8051_idata_n1574), .B(
        oc8051_ram_top1_oc8051_idata_n1575), .C(
        oc8051_ram_top1_oc8051_idata_n1576), .D(
        oc8051_ram_top1_oc8051_idata_n1577), .Y(
        oc8051_ram_top1_oc8051_idata_n1554) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2962 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1570) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2961 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1571) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2960 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1572) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2959 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1573) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2958 ( .A(
        oc8051_ram_top1_oc8051_idata_n1570), .B(
        oc8051_ram_top1_oc8051_idata_n1571), .C(
        oc8051_ram_top1_oc8051_idata_n1572), .D(
        oc8051_ram_top1_oc8051_idata_n1573), .Y(
        oc8051_ram_top1_oc8051_idata_n1555) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2957 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1566) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2956 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1567) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2955 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1568) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2954 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1569) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2953 ( .A(
        oc8051_ram_top1_oc8051_idata_n1566), .B(
        oc8051_ram_top1_oc8051_idata_n1567), .C(
        oc8051_ram_top1_oc8051_idata_n1568), .D(
        oc8051_ram_top1_oc8051_idata_n1569), .Y(
        oc8051_ram_top1_oc8051_idata_n1556) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2952 ( .A0(
        oc8051_ram_top1_oc8051_idata_n190), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n182), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1565) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2951 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1565), .Y(
        oc8051_ram_top1_oc8051_idata_n1558) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2950 ( .A0(
        oc8051_ram_top1_oc8051_idata_n174), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n166), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1564) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2949 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1564), .Y(
        oc8051_ram_top1_oc8051_idata_n1559) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2948 ( .A0(
        oc8051_ram_top1_oc8051_idata_n158), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n150), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1563) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2947 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1563), .Y(
        oc8051_ram_top1_oc8051_idata_n1560) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2946 ( .A0(
        oc8051_ram_top1_oc8051_idata_n142), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n134), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1562) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2945 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1562), .Y(
        oc8051_ram_top1_oc8051_idata_n1561) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2944 ( .A(
        oc8051_ram_top1_oc8051_idata_n1558), .B(
        oc8051_ram_top1_oc8051_idata_n1559), .C(
        oc8051_ram_top1_oc8051_idata_n1560), .D(
        oc8051_ram_top1_oc8051_idata_n1561), .Y(
        oc8051_ram_top1_oc8051_idata_n1557) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2943 ( .A(
        oc8051_ram_top1_oc8051_idata_n1552), .B(
        oc8051_ram_top1_oc8051_idata_n1553), .C(
        oc8051_ram_top1_oc8051_idata_n1554), .D(
        oc8051_ram_top1_oc8051_idata_n1555), .E(
        oc8051_ram_top1_oc8051_idata_n1556), .F(
        oc8051_ram_top1_oc8051_idata_n1557), .Y(
        oc8051_ram_top1_oc8051_idata_n1508) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2942 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1548) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2941 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1549) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2940 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1550) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2939 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1551) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2938 ( .A(
        oc8051_ram_top1_oc8051_idata_n1548), .B(
        oc8051_ram_top1_oc8051_idata_n1549), .C(
        oc8051_ram_top1_oc8051_idata_n1550), .D(
        oc8051_ram_top1_oc8051_idata_n1551), .Y(
        oc8051_ram_top1_oc8051_idata_n1510) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2937 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1544) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2936 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1545) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2935 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1546) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2934 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1547) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2933 ( .A(
        oc8051_ram_top1_oc8051_idata_n1544), .B(
        oc8051_ram_top1_oc8051_idata_n1545), .C(
        oc8051_ram_top1_oc8051_idata_n1546), .D(
        oc8051_ram_top1_oc8051_idata_n1547), .Y(
        oc8051_ram_top1_oc8051_idata_n1511) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2932 ( .A(
        oc8051_ram_top1_oc8051_idata_n118), .Y(
        oc8051_ram_top1_oc8051_idata_n1541) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2931 ( .A(
        oc8051_ram_top1_oc8051_idata_n126), .Y(
        oc8051_ram_top1_oc8051_idata_n1542) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2930 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n744) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2929 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n753) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2928 ( .A0(
        oc8051_ram_top1_oc8051_idata_n744), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n753), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1543) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2927 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1541), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1542), .C0(
        oc8051_ram_top1_oc8051_idata_n1543), .Y(
        oc8051_ram_top1_oc8051_idata_n1532) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2926 ( .A(
        oc8051_ram_top1_oc8051_idata_n102), .Y(
        oc8051_ram_top1_oc8051_idata_n1538) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2925 ( .A(
        oc8051_ram_top1_oc8051_idata_n110), .Y(
        oc8051_ram_top1_oc8051_idata_n1539) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2924 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n723) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2923 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n733) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2922 ( .A0(
        oc8051_ram_top1_oc8051_idata_n723), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n733), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1540) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2921 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1538), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1539), .C0(
        oc8051_ram_top1_oc8051_idata_n1540), .Y(
        oc8051_ram_top1_oc8051_idata_n1533) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2920 ( .A0(
        oc8051_ram_top1_oc8051_idata_n94), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n86), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1537) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2919 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1537), .Y(
        oc8051_ram_top1_oc8051_idata_n1534) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2918 ( .A0(
        oc8051_ram_top1_oc8051_idata_n78), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n70), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1536) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2917 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1536), .Y(
        oc8051_ram_top1_oc8051_idata_n1535) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2916 ( .A(
        oc8051_ram_top1_oc8051_idata_n1532), .B(
        oc8051_ram_top1_oc8051_idata_n1533), .C(
        oc8051_ram_top1_oc8051_idata_n1534), .D(
        oc8051_ram_top1_oc8051_idata_n1535), .Y(
        oc8051_ram_top1_oc8051_idata_n1512) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2915 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1528) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2914 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1529) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2913 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1530) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2912 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1531) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2911 ( .A(
        oc8051_ram_top1_oc8051_idata_n1528), .B(
        oc8051_ram_top1_oc8051_idata_n1529), .C(
        oc8051_ram_top1_oc8051_idata_n1530), .D(
        oc8051_ram_top1_oc8051_idata_n1531), .Y(
        oc8051_ram_top1_oc8051_idata_n1513) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2910 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1524) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2909 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1525) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2908 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1526) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2907 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__5_), .Y(
        oc8051_ram_top1_oc8051_idata_n1527) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2906 ( .A(
        oc8051_ram_top1_oc8051_idata_n1524), .B(
        oc8051_ram_top1_oc8051_idata_n1525), .C(
        oc8051_ram_top1_oc8051_idata_n1526), .D(
        oc8051_ram_top1_oc8051_idata_n1527), .Y(
        oc8051_ram_top1_oc8051_idata_n1514) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2905 ( .A0(
        oc8051_ram_top1_oc8051_idata_n62), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n54), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1523) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2904 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1523), .Y(
        oc8051_ram_top1_oc8051_idata_n1516) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2903 ( .A0(
        oc8051_ram_top1_oc8051_idata_n46), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n38), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1522) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2902 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1522), .Y(
        oc8051_ram_top1_oc8051_idata_n1517) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2901 ( .A0(
        oc8051_ram_top1_oc8051_idata_n30), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n22), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1521) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2900 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1521), .Y(
        oc8051_ram_top1_oc8051_idata_n1518) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2899 ( .A0(
        oc8051_ram_top1_oc8051_idata_n14), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n6), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1520) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2898 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__5_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__5_), .C0(
        oc8051_ram_top1_oc8051_idata_n1520), .Y(
        oc8051_ram_top1_oc8051_idata_n1519) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2897 ( .A(
        oc8051_ram_top1_oc8051_idata_n1516), .B(
        oc8051_ram_top1_oc8051_idata_n1517), .C(
        oc8051_ram_top1_oc8051_idata_n1518), .D(
        oc8051_ram_top1_oc8051_idata_n1519), .Y(
        oc8051_ram_top1_oc8051_idata_n1515) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2896 ( .A(
        oc8051_ram_top1_oc8051_idata_n1510), .B(
        oc8051_ram_top1_oc8051_idata_n1511), .C(
        oc8051_ram_top1_oc8051_idata_n1512), .D(
        oc8051_ram_top1_oc8051_idata_n1513), .E(
        oc8051_ram_top1_oc8051_idata_n1514), .F(
        oc8051_ram_top1_oc8051_idata_n1515), .Y(
        oc8051_ram_top1_oc8051_idata_n1509) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2895 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n1507), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n1508), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n1509), .Y(
        oc8051_ram_top1_oc8051_idata_n1506) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2894 ( .A0(
        oc8051_ram_top1_oc8051_idata_n613), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n1505), .C0(
        oc8051_ram_top1_oc8051_idata_n1506), .Y(
        oc8051_ram_top1_oc8051_idata_n2480) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2893 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1501) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2892 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1502) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2891 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1503) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2890 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1504) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2889 ( .A(
        oc8051_ram_top1_oc8051_idata_n1501), .B(
        oc8051_ram_top1_oc8051_idata_n1502), .C(
        oc8051_ram_top1_oc8051_idata_n1503), .D(
        oc8051_ram_top1_oc8051_idata_n1504), .Y(
        oc8051_ram_top1_oc8051_idata_n1463) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2888 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1497) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2887 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1498) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2886 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1499) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2885 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1500) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2884 ( .A(
        oc8051_ram_top1_oc8051_idata_n1497), .B(
        oc8051_ram_top1_oc8051_idata_n1498), .C(
        oc8051_ram_top1_oc8051_idata_n1499), .D(
        oc8051_ram_top1_oc8051_idata_n1500), .Y(
        oc8051_ram_top1_oc8051_idata_n1464) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2883 ( .A(
        oc8051_ram_top1_oc8051_idata_n501), .Y(
        oc8051_ram_top1_oc8051_idata_n1494) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2882 ( .A(
        oc8051_ram_top1_oc8051_idata_n509), .Y(
        oc8051_ram_top1_oc8051_idata_n1495) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2881 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1056) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2880 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1066) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2879 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1056), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1066), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1496) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2878 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1494), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1495), .C0(
        oc8051_ram_top1_oc8051_idata_n1496), .Y(
        oc8051_ram_top1_oc8051_idata_n1485) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2877 ( .A(
        oc8051_ram_top1_oc8051_idata_n485), .Y(
        oc8051_ram_top1_oc8051_idata_n1491) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2876 ( .A(
        oc8051_ram_top1_oc8051_idata_n493), .Y(
        oc8051_ram_top1_oc8051_idata_n1492) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2875 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1030) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2874 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1042) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2873 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1030), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1042), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1493) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2872 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1491), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1492), .C0(
        oc8051_ram_top1_oc8051_idata_n1493), .Y(
        oc8051_ram_top1_oc8051_idata_n1486) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2871 ( .A0(
        oc8051_ram_top1_oc8051_idata_n477), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n469), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1490) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2870 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1490), .Y(
        oc8051_ram_top1_oc8051_idata_n1487) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2869 ( .A0(
        oc8051_ram_top1_oc8051_idata_n461), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n453), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1489) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2868 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1489), .Y(
        oc8051_ram_top1_oc8051_idata_n1488) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2867 ( .A(
        oc8051_ram_top1_oc8051_idata_n1485), .B(
        oc8051_ram_top1_oc8051_idata_n1486), .C(
        oc8051_ram_top1_oc8051_idata_n1487), .D(
        oc8051_ram_top1_oc8051_idata_n1488), .Y(
        oc8051_ram_top1_oc8051_idata_n1465) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2866 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1481) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2865 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1482) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2864 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1483) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2863 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1484) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2862 ( .A(
        oc8051_ram_top1_oc8051_idata_n1481), .B(
        oc8051_ram_top1_oc8051_idata_n1482), .C(
        oc8051_ram_top1_oc8051_idata_n1483), .D(
        oc8051_ram_top1_oc8051_idata_n1484), .Y(
        oc8051_ram_top1_oc8051_idata_n1466) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2861 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1477) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2860 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1478) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2859 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1479) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2858 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1480) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2857 ( .A(
        oc8051_ram_top1_oc8051_idata_n1477), .B(
        oc8051_ram_top1_oc8051_idata_n1478), .C(
        oc8051_ram_top1_oc8051_idata_n1479), .D(
        oc8051_ram_top1_oc8051_idata_n1480), .Y(
        oc8051_ram_top1_oc8051_idata_n1467) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2856 ( .A0(
        oc8051_ram_top1_oc8051_idata_n445), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n437), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1476) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2855 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1476), .Y(
        oc8051_ram_top1_oc8051_idata_n1469) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2854 ( .A0(
        oc8051_ram_top1_oc8051_idata_n429), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n421), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1475) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2853 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1475), .Y(
        oc8051_ram_top1_oc8051_idata_n1470) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2852 ( .A0(
        oc8051_ram_top1_oc8051_idata_n413), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n405), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1474) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2851 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1474), .Y(
        oc8051_ram_top1_oc8051_idata_n1471) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2850 ( .A0(
        oc8051_ram_top1_oc8051_idata_n397), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n389), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1473) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2849 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1473), .Y(
        oc8051_ram_top1_oc8051_idata_n1472) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2848 ( .A(
        oc8051_ram_top1_oc8051_idata_n1469), .B(
        oc8051_ram_top1_oc8051_idata_n1470), .C(
        oc8051_ram_top1_oc8051_idata_n1471), .D(
        oc8051_ram_top1_oc8051_idata_n1472), .Y(
        oc8051_ram_top1_oc8051_idata_n1468) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2847 ( .A(
        oc8051_ram_top1_oc8051_idata_n1463), .B(
        oc8051_ram_top1_oc8051_idata_n1464), .C(
        oc8051_ram_top1_oc8051_idata_n1465), .D(
        oc8051_ram_top1_oc8051_idata_n1466), .E(
        oc8051_ram_top1_oc8051_idata_n1467), .F(
        oc8051_ram_top1_oc8051_idata_n1468), .Y(
        oc8051_ram_top1_oc8051_idata_n1462) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2846 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n1462), .B0(oc8051_ram_top1_rd_data_m[6]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n1331) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2845 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1458) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2844 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1459) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2843 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1460) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2842 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1461) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2841 ( .A(
        oc8051_ram_top1_oc8051_idata_n1458), .B(
        oc8051_ram_top1_oc8051_idata_n1459), .C(
        oc8051_ram_top1_oc8051_idata_n1460), .D(
        oc8051_ram_top1_oc8051_idata_n1461), .Y(
        oc8051_ram_top1_oc8051_idata_n1420) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2840 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1454) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2839 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1455) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2838 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1456) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2837 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1457) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2836 ( .A(
        oc8051_ram_top1_oc8051_idata_n1454), .B(
        oc8051_ram_top1_oc8051_idata_n1455), .C(
        oc8051_ram_top1_oc8051_idata_n1456), .D(
        oc8051_ram_top1_oc8051_idata_n1457), .Y(
        oc8051_ram_top1_oc8051_idata_n1421) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2835 ( .A(
        oc8051_ram_top1_oc8051_idata_n373), .Y(
        oc8051_ram_top1_oc8051_idata_n1451) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2834 ( .A(
        oc8051_ram_top1_oc8051_idata_n381), .Y(
        oc8051_ram_top1_oc8051_idata_n1452) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2833 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n948) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2832 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n957) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2831 ( .A0(
        oc8051_ram_top1_oc8051_idata_n948), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n957), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1453) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2830 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1451), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1452), .C0(
        oc8051_ram_top1_oc8051_idata_n1453), .Y(
        oc8051_ram_top1_oc8051_idata_n1442) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2829 ( .A(
        oc8051_ram_top1_oc8051_idata_n357), .Y(
        oc8051_ram_top1_oc8051_idata_n1448) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2828 ( .A(
        oc8051_ram_top1_oc8051_idata_n365), .Y(
        oc8051_ram_top1_oc8051_idata_n1449) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2827 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n927) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2826 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n937) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2825 ( .A0(
        oc8051_ram_top1_oc8051_idata_n927), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n937), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1450) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2824 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1448), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1449), .C0(
        oc8051_ram_top1_oc8051_idata_n1450), .Y(
        oc8051_ram_top1_oc8051_idata_n1443) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2823 ( .A0(
        oc8051_ram_top1_oc8051_idata_n349), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n341), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1447) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2822 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1447), .Y(
        oc8051_ram_top1_oc8051_idata_n1444) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2821 ( .A0(
        oc8051_ram_top1_oc8051_idata_n333), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n325), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1446) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2820 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1446), .Y(
        oc8051_ram_top1_oc8051_idata_n1445) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2819 ( .A(
        oc8051_ram_top1_oc8051_idata_n1442), .B(
        oc8051_ram_top1_oc8051_idata_n1443), .C(
        oc8051_ram_top1_oc8051_idata_n1444), .D(
        oc8051_ram_top1_oc8051_idata_n1445), .Y(
        oc8051_ram_top1_oc8051_idata_n1422) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2818 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1438) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2817 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1439) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2816 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1440) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2815 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1441) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2814 ( .A(
        oc8051_ram_top1_oc8051_idata_n1438), .B(
        oc8051_ram_top1_oc8051_idata_n1439), .C(
        oc8051_ram_top1_oc8051_idata_n1440), .D(
        oc8051_ram_top1_oc8051_idata_n1441), .Y(
        oc8051_ram_top1_oc8051_idata_n1423) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2813 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1434) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2812 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1435) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2811 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1436) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2810 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1437) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2809 ( .A(
        oc8051_ram_top1_oc8051_idata_n1434), .B(
        oc8051_ram_top1_oc8051_idata_n1435), .C(
        oc8051_ram_top1_oc8051_idata_n1436), .D(
        oc8051_ram_top1_oc8051_idata_n1437), .Y(
        oc8051_ram_top1_oc8051_idata_n1424) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2808 ( .A0(
        oc8051_ram_top1_oc8051_idata_n317), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n309), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1433) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2807 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1433), .Y(
        oc8051_ram_top1_oc8051_idata_n1426) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2806 ( .A0(
        oc8051_ram_top1_oc8051_idata_n301), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n293), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1432) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2805 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1432), .Y(
        oc8051_ram_top1_oc8051_idata_n1427) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2804 ( .A0(
        oc8051_ram_top1_oc8051_idata_n285), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n277), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1431) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2803 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1431), .Y(
        oc8051_ram_top1_oc8051_idata_n1428) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2802 ( .A0(
        oc8051_ram_top1_oc8051_idata_n269), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n261), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1430) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2801 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1430), .Y(
        oc8051_ram_top1_oc8051_idata_n1429) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2800 ( .A(
        oc8051_ram_top1_oc8051_idata_n1426), .B(
        oc8051_ram_top1_oc8051_idata_n1427), .C(
        oc8051_ram_top1_oc8051_idata_n1428), .D(
        oc8051_ram_top1_oc8051_idata_n1429), .Y(
        oc8051_ram_top1_oc8051_idata_n1425) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2799 ( .A(
        oc8051_ram_top1_oc8051_idata_n1420), .B(
        oc8051_ram_top1_oc8051_idata_n1421), .C(
        oc8051_ram_top1_oc8051_idata_n1422), .D(
        oc8051_ram_top1_oc8051_idata_n1423), .E(
        oc8051_ram_top1_oc8051_idata_n1424), .F(
        oc8051_ram_top1_oc8051_idata_n1425), .Y(
        oc8051_ram_top1_oc8051_idata_n1333) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2798 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1416) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2797 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1417) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2796 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1418) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2795 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1419) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2794 ( .A(
        oc8051_ram_top1_oc8051_idata_n1416), .B(
        oc8051_ram_top1_oc8051_idata_n1417), .C(
        oc8051_ram_top1_oc8051_idata_n1418), .D(
        oc8051_ram_top1_oc8051_idata_n1419), .Y(
        oc8051_ram_top1_oc8051_idata_n1378) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2793 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1412) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2792 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1413) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2791 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1414) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2790 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1415) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2789 ( .A(
        oc8051_ram_top1_oc8051_idata_n1412), .B(
        oc8051_ram_top1_oc8051_idata_n1413), .C(
        oc8051_ram_top1_oc8051_idata_n1414), .D(
        oc8051_ram_top1_oc8051_idata_n1415), .Y(
        oc8051_ram_top1_oc8051_idata_n1379) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2788 ( .A(
        oc8051_ram_top1_oc8051_idata_n245), .Y(
        oc8051_ram_top1_oc8051_idata_n1409) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2787 ( .A(
        oc8051_ram_top1_oc8051_idata_n253), .Y(
        oc8051_ram_top1_oc8051_idata_n1410) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2786 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n846) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2785 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n855) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2784 ( .A0(
        oc8051_ram_top1_oc8051_idata_n846), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n855), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1411) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2783 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1409), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1410), .C0(
        oc8051_ram_top1_oc8051_idata_n1411), .Y(
        oc8051_ram_top1_oc8051_idata_n1400) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2782 ( .A(
        oc8051_ram_top1_oc8051_idata_n229), .Y(
        oc8051_ram_top1_oc8051_idata_n1406) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2781 ( .A(
        oc8051_ram_top1_oc8051_idata_n237), .Y(
        oc8051_ram_top1_oc8051_idata_n1407) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2780 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n825) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2779 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n835) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2778 ( .A0(
        oc8051_ram_top1_oc8051_idata_n825), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n835), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1408) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2777 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1406), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1407), .C0(
        oc8051_ram_top1_oc8051_idata_n1408), .Y(
        oc8051_ram_top1_oc8051_idata_n1401) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2776 ( .A0(
        oc8051_ram_top1_oc8051_idata_n221), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n213), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1405) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2775 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1405), .Y(
        oc8051_ram_top1_oc8051_idata_n1402) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2774 ( .A0(
        oc8051_ram_top1_oc8051_idata_n205), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n197), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1404) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2773 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1404), .Y(
        oc8051_ram_top1_oc8051_idata_n1403) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2772 ( .A(
        oc8051_ram_top1_oc8051_idata_n1400), .B(
        oc8051_ram_top1_oc8051_idata_n1401), .C(
        oc8051_ram_top1_oc8051_idata_n1402), .D(
        oc8051_ram_top1_oc8051_idata_n1403), .Y(
        oc8051_ram_top1_oc8051_idata_n1380) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2771 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1396) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2770 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1397) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2769 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1398) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2768 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1399) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2767 ( .A(
        oc8051_ram_top1_oc8051_idata_n1396), .B(
        oc8051_ram_top1_oc8051_idata_n1397), .C(
        oc8051_ram_top1_oc8051_idata_n1398), .D(
        oc8051_ram_top1_oc8051_idata_n1399), .Y(
        oc8051_ram_top1_oc8051_idata_n1381) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2766 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1392) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2765 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1393) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2764 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1394) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2763 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1395) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2762 ( .A(
        oc8051_ram_top1_oc8051_idata_n1392), .B(
        oc8051_ram_top1_oc8051_idata_n1393), .C(
        oc8051_ram_top1_oc8051_idata_n1394), .D(
        oc8051_ram_top1_oc8051_idata_n1395), .Y(
        oc8051_ram_top1_oc8051_idata_n1382) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2761 ( .A0(
        oc8051_ram_top1_oc8051_idata_n189), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n181), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1391) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2760 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1391), .Y(
        oc8051_ram_top1_oc8051_idata_n1384) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2759 ( .A0(
        oc8051_ram_top1_oc8051_idata_n173), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n165), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1390) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2758 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1390), .Y(
        oc8051_ram_top1_oc8051_idata_n1385) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2757 ( .A0(
        oc8051_ram_top1_oc8051_idata_n157), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n149), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1389) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2756 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1389), .Y(
        oc8051_ram_top1_oc8051_idata_n1386) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2755 ( .A0(
        oc8051_ram_top1_oc8051_idata_n141), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n133), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1388) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2754 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1388), .Y(
        oc8051_ram_top1_oc8051_idata_n1387) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2753 ( .A(
        oc8051_ram_top1_oc8051_idata_n1384), .B(
        oc8051_ram_top1_oc8051_idata_n1385), .C(
        oc8051_ram_top1_oc8051_idata_n1386), .D(
        oc8051_ram_top1_oc8051_idata_n1387), .Y(
        oc8051_ram_top1_oc8051_idata_n1383) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2752 ( .A(
        oc8051_ram_top1_oc8051_idata_n1378), .B(
        oc8051_ram_top1_oc8051_idata_n1379), .C(
        oc8051_ram_top1_oc8051_idata_n1380), .D(
        oc8051_ram_top1_oc8051_idata_n1381), .E(
        oc8051_ram_top1_oc8051_idata_n1382), .F(
        oc8051_ram_top1_oc8051_idata_n1383), .Y(
        oc8051_ram_top1_oc8051_idata_n1334) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2751 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1374) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2750 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1375) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2749 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1376) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2748 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1377) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2747 ( .A(
        oc8051_ram_top1_oc8051_idata_n1374), .B(
        oc8051_ram_top1_oc8051_idata_n1375), .C(
        oc8051_ram_top1_oc8051_idata_n1376), .D(
        oc8051_ram_top1_oc8051_idata_n1377), .Y(
        oc8051_ram_top1_oc8051_idata_n1336) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2746 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1370) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2745 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1371) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2744 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1372) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2743 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1373) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2742 ( .A(
        oc8051_ram_top1_oc8051_idata_n1370), .B(
        oc8051_ram_top1_oc8051_idata_n1371), .C(
        oc8051_ram_top1_oc8051_idata_n1372), .D(
        oc8051_ram_top1_oc8051_idata_n1373), .Y(
        oc8051_ram_top1_oc8051_idata_n1337) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2741 ( .A(
        oc8051_ram_top1_oc8051_idata_n117), .Y(
        oc8051_ram_top1_oc8051_idata_n1367) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2740 ( .A(
        oc8051_ram_top1_oc8051_idata_n125), .Y(
        oc8051_ram_top1_oc8051_idata_n1368) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2739 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n743) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2738 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n752) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2737 ( .A0(
        oc8051_ram_top1_oc8051_idata_n743), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n752), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1369) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2736 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1367), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1368), .C0(
        oc8051_ram_top1_oc8051_idata_n1369), .Y(
        oc8051_ram_top1_oc8051_idata_n1358) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2735 ( .A(
        oc8051_ram_top1_oc8051_idata_n101), .Y(
        oc8051_ram_top1_oc8051_idata_n1364) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2734 ( .A(
        oc8051_ram_top1_oc8051_idata_n109), .Y(
        oc8051_ram_top1_oc8051_idata_n1365) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2733 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n722) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2732 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n732) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2731 ( .A0(
        oc8051_ram_top1_oc8051_idata_n722), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n732), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1366) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2730 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1364), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1365), .C0(
        oc8051_ram_top1_oc8051_idata_n1366), .Y(
        oc8051_ram_top1_oc8051_idata_n1359) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2729 ( .A0(
        oc8051_ram_top1_oc8051_idata_n93), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n85), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1363) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2728 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1363), .Y(
        oc8051_ram_top1_oc8051_idata_n1360) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2727 ( .A0(
        oc8051_ram_top1_oc8051_idata_n77), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n69), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1362) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2726 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1362), .Y(
        oc8051_ram_top1_oc8051_idata_n1361) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2725 ( .A(
        oc8051_ram_top1_oc8051_idata_n1358), .B(
        oc8051_ram_top1_oc8051_idata_n1359), .C(
        oc8051_ram_top1_oc8051_idata_n1360), .D(
        oc8051_ram_top1_oc8051_idata_n1361), .Y(
        oc8051_ram_top1_oc8051_idata_n1338) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2724 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1354) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2723 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1355) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2722 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1356) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2721 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1357) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2720 ( .A(
        oc8051_ram_top1_oc8051_idata_n1354), .B(
        oc8051_ram_top1_oc8051_idata_n1355), .C(
        oc8051_ram_top1_oc8051_idata_n1356), .D(
        oc8051_ram_top1_oc8051_idata_n1357), .Y(
        oc8051_ram_top1_oc8051_idata_n1339) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2719 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1350) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2718 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1351) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2717 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1352) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2716 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__6_), .Y(
        oc8051_ram_top1_oc8051_idata_n1353) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2715 ( .A(
        oc8051_ram_top1_oc8051_idata_n1350), .B(
        oc8051_ram_top1_oc8051_idata_n1351), .C(
        oc8051_ram_top1_oc8051_idata_n1352), .D(
        oc8051_ram_top1_oc8051_idata_n1353), .Y(
        oc8051_ram_top1_oc8051_idata_n1340) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2714 ( .A0(
        oc8051_ram_top1_oc8051_idata_n61), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n53), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1349) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2713 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1349), .Y(
        oc8051_ram_top1_oc8051_idata_n1342) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2712 ( .A0(
        oc8051_ram_top1_oc8051_idata_n45), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n37), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1348) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2711 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1348), .Y(
        oc8051_ram_top1_oc8051_idata_n1343) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2710 ( .A0(
        oc8051_ram_top1_oc8051_idata_n29), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n21), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1347) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2709 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1347), .Y(
        oc8051_ram_top1_oc8051_idata_n1344) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2708 ( .A0(
        oc8051_ram_top1_oc8051_idata_n13), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n5), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1346) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2707 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__6_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__6_), .C0(
        oc8051_ram_top1_oc8051_idata_n1346), .Y(
        oc8051_ram_top1_oc8051_idata_n1345) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2706 ( .A(
        oc8051_ram_top1_oc8051_idata_n1342), .B(
        oc8051_ram_top1_oc8051_idata_n1343), .C(
        oc8051_ram_top1_oc8051_idata_n1344), .D(
        oc8051_ram_top1_oc8051_idata_n1345), .Y(
        oc8051_ram_top1_oc8051_idata_n1341) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2705 ( .A(
        oc8051_ram_top1_oc8051_idata_n1336), .B(
        oc8051_ram_top1_oc8051_idata_n1337), .C(
        oc8051_ram_top1_oc8051_idata_n1338), .D(
        oc8051_ram_top1_oc8051_idata_n1339), .E(
        oc8051_ram_top1_oc8051_idata_n1340), .F(
        oc8051_ram_top1_oc8051_idata_n1341), .Y(
        oc8051_ram_top1_oc8051_idata_n1335) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2704 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n1333), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n1334), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n1335), .Y(
        oc8051_ram_top1_oc8051_idata_n1332) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2703 ( .A0(
        oc8051_ram_top1_oc8051_idata_n630), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n1331), .C0(
        oc8051_ram_top1_oc8051_idata_n1332), .Y(
        oc8051_ram_top1_oc8051_idata_n2481) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2702 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_232__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_233__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1327) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2701 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_234__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_235__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1328) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2700 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_239__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_251__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1329) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2699 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_238__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_250__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1330) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2698 ( .A(
        oc8051_ram_top1_oc8051_idata_n1327), .B(
        oc8051_ram_top1_oc8051_idata_n1328), .C(
        oc8051_ram_top1_oc8051_idata_n1329), .D(
        oc8051_ram_top1_oc8051_idata_n1330), .Y(
        oc8051_ram_top1_oc8051_idata_n1289) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2697 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_237__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_249__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1323) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2696 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_236__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_248__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1324) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2695 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_255__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_254__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1325) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2694 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_253__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_252__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1326) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2693 ( .A(
        oc8051_ram_top1_oc8051_idata_n1323), .B(
        oc8051_ram_top1_oc8051_idata_n1324), .C(
        oc8051_ram_top1_oc8051_idata_n1325), .D(
        oc8051_ram_top1_oc8051_idata_n1326), .Y(
        oc8051_ram_top1_oc8051_idata_n1290) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2692 ( .A(
        oc8051_ram_top1_oc8051_idata_n500), .Y(
        oc8051_ram_top1_oc8051_idata_n1320) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2691 ( .A(
        oc8051_ram_top1_oc8051_idata_n508), .Y(
        oc8051_ram_top1_oc8051_idata_n1321) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2690 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_244__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1054) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2689 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_245__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1064) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2688 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1054), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n1064), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1322) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2687 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1320), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1321), .C0(
        oc8051_ram_top1_oc8051_idata_n1322), .Y(
        oc8051_ram_top1_oc8051_idata_n1311) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2686 ( .A(
        oc8051_ram_top1_oc8051_idata_n484), .Y(
        oc8051_ram_top1_oc8051_idata_n1317) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2685 ( .A(
        oc8051_ram_top1_oc8051_idata_n492), .Y(
        oc8051_ram_top1_oc8051_idata_n1318) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2684 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_240__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1028) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2683 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_241__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1040) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2682 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1028), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n1040), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1319) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2681 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1317), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1318), .C0(
        oc8051_ram_top1_oc8051_idata_n1319), .Y(
        oc8051_ram_top1_oc8051_idata_n1312) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2680 ( .A0(
        oc8051_ram_top1_oc8051_idata_n476), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n468), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1316) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2679 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_231__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_230__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1316), .Y(
        oc8051_ram_top1_oc8051_idata_n1313) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2678 ( .A0(
        oc8051_ram_top1_oc8051_idata_n460), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n452), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1315) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2677 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_227__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_226__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1315), .Y(
        oc8051_ram_top1_oc8051_idata_n1314) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2676 ( .A(
        oc8051_ram_top1_oc8051_idata_n1311), .B(
        oc8051_ram_top1_oc8051_idata_n1312), .C(
        oc8051_ram_top1_oc8051_idata_n1313), .D(
        oc8051_ram_top1_oc8051_idata_n1314), .Y(
        oc8051_ram_top1_oc8051_idata_n1291) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2675 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_223__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_222__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1307) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2674 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_221__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_220__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1308) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2673 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_219__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_218__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1309) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2672 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_217__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_216__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1310) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2671 ( .A(
        oc8051_ram_top1_oc8051_idata_n1307), .B(
        oc8051_ram_top1_oc8051_idata_n1308), .C(
        oc8051_ram_top1_oc8051_idata_n1309), .D(
        oc8051_ram_top1_oc8051_idata_n1310), .Y(
        oc8051_ram_top1_oc8051_idata_n1292) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2670 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_215__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_214__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1303) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2669 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_213__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_212__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1304) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2668 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_211__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_210__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1305) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2667 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_209__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_208__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1306) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2666 ( .A(
        oc8051_ram_top1_oc8051_idata_n1303), .B(
        oc8051_ram_top1_oc8051_idata_n1304), .C(
        oc8051_ram_top1_oc8051_idata_n1305), .D(
        oc8051_ram_top1_oc8051_idata_n1306), .Y(
        oc8051_ram_top1_oc8051_idata_n1293) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2665 ( .A0(
        oc8051_ram_top1_oc8051_idata_n444), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n436), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1302) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2664 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_205__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_204__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1302), .Y(
        oc8051_ram_top1_oc8051_idata_n1295) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2663 ( .A0(
        oc8051_ram_top1_oc8051_idata_n428), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n420), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1301) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2662 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_203__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_202__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1301), .Y(
        oc8051_ram_top1_oc8051_idata_n1296) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2661 ( .A0(
        oc8051_ram_top1_oc8051_idata_n412), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n404), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1300) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2660 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_199__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_198__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1300), .Y(
        oc8051_ram_top1_oc8051_idata_n1297) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2659 ( .A0(
        oc8051_ram_top1_oc8051_idata_n396), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n388), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1299) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2658 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_195__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_194__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1299), .Y(
        oc8051_ram_top1_oc8051_idata_n1298) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2657 ( .A(
        oc8051_ram_top1_oc8051_idata_n1295), .B(
        oc8051_ram_top1_oc8051_idata_n1296), .C(
        oc8051_ram_top1_oc8051_idata_n1297), .D(
        oc8051_ram_top1_oc8051_idata_n1298), .Y(
        oc8051_ram_top1_oc8051_idata_n1294) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2656 ( .A(
        oc8051_ram_top1_oc8051_idata_n1289), .B(
        oc8051_ram_top1_oc8051_idata_n1290), .C(
        oc8051_ram_top1_oc8051_idata_n1291), .D(
        oc8051_ram_top1_oc8051_idata_n1292), .E(
        oc8051_ram_top1_oc8051_idata_n1293), .F(
        oc8051_ram_top1_oc8051_idata_n1294), .Y(
        oc8051_ram_top1_oc8051_idata_n1287) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2655 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1286), .A1(
        oc8051_ram_top1_oc8051_idata_n1287), .B0(oc8051_ram_top1_rd_data_m[7]), 
        .B1(oc8051_ram_top1_oc8051_idata_n1288), .Y(
        oc8051_ram_top1_oc8051_idata_n1088) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2654 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_168__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_169__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1282) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2653 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_170__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_171__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1283) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2652 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_175__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_187__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1284) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2651 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_174__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_186__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1285) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2650 ( .A(
        oc8051_ram_top1_oc8051_idata_n1282), .B(
        oc8051_ram_top1_oc8051_idata_n1283), .C(
        oc8051_ram_top1_oc8051_idata_n1284), .D(
        oc8051_ram_top1_oc8051_idata_n1285), .Y(
        oc8051_ram_top1_oc8051_idata_n1244) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2649 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_173__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_185__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1278) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2648 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_172__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_184__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1279) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2647 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_191__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_190__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1280) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2646 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_189__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_188__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1281) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2645 ( .A(
        oc8051_ram_top1_oc8051_idata_n1278), .B(
        oc8051_ram_top1_oc8051_idata_n1279), .C(
        oc8051_ram_top1_oc8051_idata_n1280), .D(
        oc8051_ram_top1_oc8051_idata_n1281), .Y(
        oc8051_ram_top1_oc8051_idata_n1245) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2644 ( .A(
        oc8051_ram_top1_oc8051_idata_n372), .Y(
        oc8051_ram_top1_oc8051_idata_n1275) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2643 ( .A(
        oc8051_ram_top1_oc8051_idata_n380), .Y(
        oc8051_ram_top1_oc8051_idata_n1276) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2642 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_180__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n946) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2641 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_181__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n955) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2640 ( .A0(
        oc8051_ram_top1_oc8051_idata_n946), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n955), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1277) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2639 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1275), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1276), .C0(
        oc8051_ram_top1_oc8051_idata_n1277), .Y(
        oc8051_ram_top1_oc8051_idata_n1266) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2638 ( .A(
        oc8051_ram_top1_oc8051_idata_n356), .Y(
        oc8051_ram_top1_oc8051_idata_n1272) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2637 ( .A(
        oc8051_ram_top1_oc8051_idata_n364), .Y(
        oc8051_ram_top1_oc8051_idata_n1273) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2636 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_176__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n925) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2635 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_177__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n935) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2634 ( .A0(
        oc8051_ram_top1_oc8051_idata_n925), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n935), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1274) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2633 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1272), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1273), .C0(
        oc8051_ram_top1_oc8051_idata_n1274), .Y(
        oc8051_ram_top1_oc8051_idata_n1267) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2632 ( .A0(
        oc8051_ram_top1_oc8051_idata_n348), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n340), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1271) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2631 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_167__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_166__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1271), .Y(
        oc8051_ram_top1_oc8051_idata_n1268) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2630 ( .A0(
        oc8051_ram_top1_oc8051_idata_n332), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n324), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1270) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2629 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_163__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_162__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1270), .Y(
        oc8051_ram_top1_oc8051_idata_n1269) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2628 ( .A(
        oc8051_ram_top1_oc8051_idata_n1266), .B(
        oc8051_ram_top1_oc8051_idata_n1267), .C(
        oc8051_ram_top1_oc8051_idata_n1268), .D(
        oc8051_ram_top1_oc8051_idata_n1269), .Y(
        oc8051_ram_top1_oc8051_idata_n1246) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2627 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_159__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_158__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1262) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2626 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_157__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_156__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1263) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2625 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_155__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_154__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1264) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2624 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_153__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_152__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1265) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2623 ( .A(
        oc8051_ram_top1_oc8051_idata_n1262), .B(
        oc8051_ram_top1_oc8051_idata_n1263), .C(
        oc8051_ram_top1_oc8051_idata_n1264), .D(
        oc8051_ram_top1_oc8051_idata_n1265), .Y(
        oc8051_ram_top1_oc8051_idata_n1247) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2622 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_151__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_150__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1258) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2621 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_149__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_148__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1259) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2620 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_147__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_146__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1260) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2619 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_145__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_144__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1261) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2618 ( .A(
        oc8051_ram_top1_oc8051_idata_n1258), .B(
        oc8051_ram_top1_oc8051_idata_n1259), .C(
        oc8051_ram_top1_oc8051_idata_n1260), .D(
        oc8051_ram_top1_oc8051_idata_n1261), .Y(
        oc8051_ram_top1_oc8051_idata_n1248) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2617 ( .A0(
        oc8051_ram_top1_oc8051_idata_n316), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n308), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1257) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2616 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_141__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_140__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1257), .Y(
        oc8051_ram_top1_oc8051_idata_n1250) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2615 ( .A0(
        oc8051_ram_top1_oc8051_idata_n300), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n292), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1256) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2614 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_139__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_138__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1256), .Y(
        oc8051_ram_top1_oc8051_idata_n1251) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2613 ( .A0(
        oc8051_ram_top1_oc8051_idata_n284), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n276), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1255) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2612 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_135__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_134__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1255), .Y(
        oc8051_ram_top1_oc8051_idata_n1252) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2611 ( .A0(
        oc8051_ram_top1_oc8051_idata_n268), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n260), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1254) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2610 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_131__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_130__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1254), .Y(
        oc8051_ram_top1_oc8051_idata_n1253) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2609 ( .A(
        oc8051_ram_top1_oc8051_idata_n1250), .B(
        oc8051_ram_top1_oc8051_idata_n1251), .C(
        oc8051_ram_top1_oc8051_idata_n1252), .D(
        oc8051_ram_top1_oc8051_idata_n1253), .Y(
        oc8051_ram_top1_oc8051_idata_n1249) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2608 ( .A(
        oc8051_ram_top1_oc8051_idata_n1244), .B(
        oc8051_ram_top1_oc8051_idata_n1245), .C(
        oc8051_ram_top1_oc8051_idata_n1246), .D(
        oc8051_ram_top1_oc8051_idata_n1247), .E(
        oc8051_ram_top1_oc8051_idata_n1248), .F(
        oc8051_ram_top1_oc8051_idata_n1249), .Y(
        oc8051_ram_top1_oc8051_idata_n1091) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2607 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_104__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_105__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1240) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2606 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_106__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_107__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1241) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2605 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_111__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_123__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1242) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2604 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_110__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_122__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1243) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2603 ( .A(
        oc8051_ram_top1_oc8051_idata_n1240), .B(
        oc8051_ram_top1_oc8051_idata_n1241), .C(
        oc8051_ram_top1_oc8051_idata_n1242), .D(
        oc8051_ram_top1_oc8051_idata_n1243), .Y(
        oc8051_ram_top1_oc8051_idata_n1202) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2602 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_109__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_121__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1236) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2601 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_108__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_120__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1237) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2600 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_127__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_126__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1238) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2599 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_125__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_124__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1239) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2598 ( .A(
        oc8051_ram_top1_oc8051_idata_n1236), .B(
        oc8051_ram_top1_oc8051_idata_n1237), .C(
        oc8051_ram_top1_oc8051_idata_n1238), .D(
        oc8051_ram_top1_oc8051_idata_n1239), .Y(
        oc8051_ram_top1_oc8051_idata_n1203) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2597 ( .A(
        oc8051_ram_top1_oc8051_idata_n244), .Y(
        oc8051_ram_top1_oc8051_idata_n1233) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2596 ( .A(
        oc8051_ram_top1_oc8051_idata_n252), .Y(
        oc8051_ram_top1_oc8051_idata_n1234) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2595 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_116__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n844) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2594 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_117__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n853) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2593 ( .A0(
        oc8051_ram_top1_oc8051_idata_n844), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n853), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1235) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2592 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1233), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1234), .C0(
        oc8051_ram_top1_oc8051_idata_n1235), .Y(
        oc8051_ram_top1_oc8051_idata_n1224) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2591 ( .A(
        oc8051_ram_top1_oc8051_idata_n228), .Y(
        oc8051_ram_top1_oc8051_idata_n1230) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2590 ( .A(
        oc8051_ram_top1_oc8051_idata_n236), .Y(
        oc8051_ram_top1_oc8051_idata_n1231) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2589 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_112__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n823) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2588 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_113__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n833) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2587 ( .A0(
        oc8051_ram_top1_oc8051_idata_n823), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n833), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1232) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2586 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1230), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1231), .C0(
        oc8051_ram_top1_oc8051_idata_n1232), .Y(
        oc8051_ram_top1_oc8051_idata_n1225) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2585 ( .A0(
        oc8051_ram_top1_oc8051_idata_n220), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n212), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1229) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2584 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_103__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_102__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1229), .Y(
        oc8051_ram_top1_oc8051_idata_n1226) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2583 ( .A0(
        oc8051_ram_top1_oc8051_idata_n204), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n196), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1228) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2582 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_99__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_98__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1228), .Y(
        oc8051_ram_top1_oc8051_idata_n1227) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2581 ( .A(
        oc8051_ram_top1_oc8051_idata_n1224), .B(
        oc8051_ram_top1_oc8051_idata_n1225), .C(
        oc8051_ram_top1_oc8051_idata_n1226), .D(
        oc8051_ram_top1_oc8051_idata_n1227), .Y(
        oc8051_ram_top1_oc8051_idata_n1204) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2580 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_95__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_94__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1220) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2579 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_93__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_92__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1221) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2578 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_91__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_90__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1222) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2577 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_89__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_88__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1223) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2576 ( .A(
        oc8051_ram_top1_oc8051_idata_n1220), .B(
        oc8051_ram_top1_oc8051_idata_n1221), .C(
        oc8051_ram_top1_oc8051_idata_n1222), .D(
        oc8051_ram_top1_oc8051_idata_n1223), .Y(
        oc8051_ram_top1_oc8051_idata_n1205) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2575 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_87__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_86__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1216) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2574 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_85__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_84__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1217) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2573 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_83__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_82__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1218) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2572 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_81__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_80__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1219) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2571 ( .A(
        oc8051_ram_top1_oc8051_idata_n1216), .B(
        oc8051_ram_top1_oc8051_idata_n1217), .C(
        oc8051_ram_top1_oc8051_idata_n1218), .D(
        oc8051_ram_top1_oc8051_idata_n1219), .Y(
        oc8051_ram_top1_oc8051_idata_n1206) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2570 ( .A0(
        oc8051_ram_top1_oc8051_idata_n188), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n180), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1215) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2569 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_77__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_76__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1215), .Y(
        oc8051_ram_top1_oc8051_idata_n1208) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2568 ( .A0(
        oc8051_ram_top1_oc8051_idata_n172), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n164), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1214) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2567 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_75__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_74__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1214), .Y(
        oc8051_ram_top1_oc8051_idata_n1209) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2566 ( .A0(
        oc8051_ram_top1_oc8051_idata_n156), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n148), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1213) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2565 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_71__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_70__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1213), .Y(
        oc8051_ram_top1_oc8051_idata_n1210) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2564 ( .A0(
        oc8051_ram_top1_oc8051_idata_n140), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n132), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1212) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2563 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_67__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_66__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1212), .Y(
        oc8051_ram_top1_oc8051_idata_n1211) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2562 ( .A(
        oc8051_ram_top1_oc8051_idata_n1208), .B(
        oc8051_ram_top1_oc8051_idata_n1209), .C(
        oc8051_ram_top1_oc8051_idata_n1210), .D(
        oc8051_ram_top1_oc8051_idata_n1211), .Y(
        oc8051_ram_top1_oc8051_idata_n1207) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2561 ( .A(
        oc8051_ram_top1_oc8051_idata_n1202), .B(
        oc8051_ram_top1_oc8051_idata_n1203), .C(
        oc8051_ram_top1_oc8051_idata_n1204), .D(
        oc8051_ram_top1_oc8051_idata_n1205), .E(
        oc8051_ram_top1_oc8051_idata_n1206), .F(
        oc8051_ram_top1_oc8051_idata_n1207), .Y(
        oc8051_ram_top1_oc8051_idata_n1093) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2560 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1200), .A1(
        oc8051_ram_top1_oc8051_idata_buff_40__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1201), .B1(
        oc8051_ram_top1_oc8051_idata_buff_41__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1190) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2559 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1198), .A1(
        oc8051_ram_top1_oc8051_idata_buff_42__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1199), .B1(
        oc8051_ram_top1_oc8051_idata_buff_43__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1191) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2558 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1196), .A1(
        oc8051_ram_top1_oc8051_idata_buff_47__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1197), .B1(
        oc8051_ram_top1_oc8051_idata_buff_59__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1192) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2557 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1194), .A1(
        oc8051_ram_top1_oc8051_idata_buff_46__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1195), .B1(
        oc8051_ram_top1_oc8051_idata_buff_58__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1193) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2556 ( .A(
        oc8051_ram_top1_oc8051_idata_n1190), .B(
        oc8051_ram_top1_oc8051_idata_n1191), .C(
        oc8051_ram_top1_oc8051_idata_n1192), .D(
        oc8051_ram_top1_oc8051_idata_n1193), .Y(
        oc8051_ram_top1_oc8051_idata_n1096) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2555 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1188), .A1(
        oc8051_ram_top1_oc8051_idata_buff_45__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1189), .B1(
        oc8051_ram_top1_oc8051_idata_buff_57__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1178) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2554 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1186), .A1(
        oc8051_ram_top1_oc8051_idata_buff_44__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1187), .B1(
        oc8051_ram_top1_oc8051_idata_buff_56__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1179) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2553 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1184), .A1(
        oc8051_ram_top1_oc8051_idata_buff_63__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1185), .B1(
        oc8051_ram_top1_oc8051_idata_buff_62__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1180) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2552 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1182), .A1(
        oc8051_ram_top1_oc8051_idata_buff_61__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1183), .B1(
        oc8051_ram_top1_oc8051_idata_buff_60__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1181) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2551 ( .A(
        oc8051_ram_top1_oc8051_idata_n1178), .B(
        oc8051_ram_top1_oc8051_idata_n1179), .C(
        oc8051_ram_top1_oc8051_idata_n1180), .D(
        oc8051_ram_top1_oc8051_idata_n1181), .Y(
        oc8051_ram_top1_oc8051_idata_n1097) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2550 ( .A(
        oc8051_ram_top1_oc8051_idata_n116), .Y(
        oc8051_ram_top1_oc8051_idata_n1172) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2549 ( .A(
        oc8051_ram_top1_oc8051_idata_n124), .Y(
        oc8051_ram_top1_oc8051_idata_n1174) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2548 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_52__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n741) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2547 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_53__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n750) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2546 ( .A0(
        oc8051_ram_top1_oc8051_idata_n741), .A1(
        oc8051_ram_top1_oc8051_idata_n1176), .B0(
        oc8051_ram_top1_oc8051_idata_n750), .B1(
        oc8051_ram_top1_oc8051_idata_n1177), .Y(
        oc8051_ram_top1_oc8051_idata_n1175) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2545 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1171), .A1(
        oc8051_ram_top1_oc8051_idata_n1172), .B0(
        oc8051_ram_top1_oc8051_idata_n1173), .B1(
        oc8051_ram_top1_oc8051_idata_n1174), .C0(
        oc8051_ram_top1_oc8051_idata_n1175), .Y(
        oc8051_ram_top1_oc8051_idata_n1150) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2544 ( .A(
        oc8051_ram_top1_oc8051_idata_n100), .Y(
        oc8051_ram_top1_oc8051_idata_n1165) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2543 ( .A(
        oc8051_ram_top1_oc8051_idata_n108), .Y(
        oc8051_ram_top1_oc8051_idata_n1167) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2542 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_48__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n720) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2541 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_49__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n730) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2540 ( .A0(
        oc8051_ram_top1_oc8051_idata_n720), .A1(
        oc8051_ram_top1_oc8051_idata_n1169), .B0(
        oc8051_ram_top1_oc8051_idata_n730), .B1(
        oc8051_ram_top1_oc8051_idata_n1170), .Y(
        oc8051_ram_top1_oc8051_idata_n1168) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2539 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1164), .A1(
        oc8051_ram_top1_oc8051_idata_n1165), .B0(
        oc8051_ram_top1_oc8051_idata_n1166), .B1(
        oc8051_ram_top1_oc8051_idata_n1167), .C0(
        oc8051_ram_top1_oc8051_idata_n1168), .Y(
        oc8051_ram_top1_oc8051_idata_n1151) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2538 ( .A0(
        oc8051_ram_top1_oc8051_idata_n92), .A1(
        oc8051_ram_top1_oc8051_idata_n1162), .B0(
        oc8051_ram_top1_oc8051_idata_n84), .B1(
        oc8051_ram_top1_oc8051_idata_n1163), .Y(
        oc8051_ram_top1_oc8051_idata_n1161) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2537 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1159), .A1(
        oc8051_ram_top1_oc8051_idata_buff_39__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1160), .B1(
        oc8051_ram_top1_oc8051_idata_buff_38__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1161), .Y(
        oc8051_ram_top1_oc8051_idata_n1152) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2536 ( .A0(
        oc8051_ram_top1_oc8051_idata_n76), .A1(
        oc8051_ram_top1_oc8051_idata_n1157), .B0(
        oc8051_ram_top1_oc8051_idata_n68), .B1(
        oc8051_ram_top1_oc8051_idata_n1158), .Y(
        oc8051_ram_top1_oc8051_idata_n1156) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2535 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1154), .A1(
        oc8051_ram_top1_oc8051_idata_buff_35__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1155), .B1(
        oc8051_ram_top1_oc8051_idata_buff_34__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1156), .Y(
        oc8051_ram_top1_oc8051_idata_n1153) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2534 ( .A(
        oc8051_ram_top1_oc8051_idata_n1150), .B(
        oc8051_ram_top1_oc8051_idata_n1151), .C(
        oc8051_ram_top1_oc8051_idata_n1152), .D(
        oc8051_ram_top1_oc8051_idata_n1153), .Y(
        oc8051_ram_top1_oc8051_idata_n1098) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2533 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1148), .A1(
        oc8051_ram_top1_oc8051_idata_buff_31__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1149), .B1(
        oc8051_ram_top1_oc8051_idata_buff_30__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1138) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2532 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1146), .A1(
        oc8051_ram_top1_oc8051_idata_buff_29__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1147), .B1(
        oc8051_ram_top1_oc8051_idata_buff_28__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1139) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2531 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1144), .A1(
        oc8051_ram_top1_oc8051_idata_buff_27__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1145), .B1(
        oc8051_ram_top1_oc8051_idata_buff_26__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1140) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2530 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1142), .A1(
        oc8051_ram_top1_oc8051_idata_buff_25__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1143), .B1(
        oc8051_ram_top1_oc8051_idata_buff_24__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1141) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2529 ( .A(
        oc8051_ram_top1_oc8051_idata_n1138), .B(
        oc8051_ram_top1_oc8051_idata_n1139), .C(
        oc8051_ram_top1_oc8051_idata_n1140), .D(
        oc8051_ram_top1_oc8051_idata_n1141), .Y(
        oc8051_ram_top1_oc8051_idata_n1099) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2528 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1136), .A1(
        oc8051_ram_top1_oc8051_idata_buff_23__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1137), .B1(
        oc8051_ram_top1_oc8051_idata_buff_22__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1126) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2527 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1134), .A1(
        oc8051_ram_top1_oc8051_idata_buff_21__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1135), .B1(
        oc8051_ram_top1_oc8051_idata_buff_20__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1127) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2526 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1132), .A1(
        oc8051_ram_top1_oc8051_idata_buff_19__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1133), .B1(
        oc8051_ram_top1_oc8051_idata_buff_18__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1128) );
  AOI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2525 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1130), .A1(
        oc8051_ram_top1_oc8051_idata_buff_17__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1131), .B1(
        oc8051_ram_top1_oc8051_idata_buff_16__7_), .Y(
        oc8051_ram_top1_oc8051_idata_n1129) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2524 ( .A(
        oc8051_ram_top1_oc8051_idata_n1126), .B(
        oc8051_ram_top1_oc8051_idata_n1127), .C(
        oc8051_ram_top1_oc8051_idata_n1128), .D(
        oc8051_ram_top1_oc8051_idata_n1129), .Y(
        oc8051_ram_top1_oc8051_idata_n1100) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2523 ( .A0(
        oc8051_ram_top1_oc8051_idata_n60), .A1(
        oc8051_ram_top1_oc8051_idata_n1124), .B0(
        oc8051_ram_top1_oc8051_idata_n52), .B1(
        oc8051_ram_top1_oc8051_idata_n1125), .Y(
        oc8051_ram_top1_oc8051_idata_n1123) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2522 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1121), .A1(
        oc8051_ram_top1_oc8051_idata_buff_13__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1122), .B1(
        oc8051_ram_top1_oc8051_idata_buff_12__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1123), .Y(
        oc8051_ram_top1_oc8051_idata_n1102) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2521 ( .A0(
        oc8051_ram_top1_oc8051_idata_n44), .A1(
        oc8051_ram_top1_oc8051_idata_n1119), .B0(
        oc8051_ram_top1_oc8051_idata_n36), .B1(
        oc8051_ram_top1_oc8051_idata_n1120), .Y(
        oc8051_ram_top1_oc8051_idata_n1118) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2520 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1116), .A1(
        oc8051_ram_top1_oc8051_idata_buff_11__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1117), .B1(
        oc8051_ram_top1_oc8051_idata_buff_10__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1118), .Y(
        oc8051_ram_top1_oc8051_idata_n1103) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2519 ( .A0(
        oc8051_ram_top1_oc8051_idata_n28), .A1(
        oc8051_ram_top1_oc8051_idata_n1114), .B0(
        oc8051_ram_top1_oc8051_idata_n20), .B1(
        oc8051_ram_top1_oc8051_idata_n1115), .Y(
        oc8051_ram_top1_oc8051_idata_n1113) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2518 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1111), .A1(
        oc8051_ram_top1_oc8051_idata_buff_7__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1112), .B1(
        oc8051_ram_top1_oc8051_idata_buff_6__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1113), .Y(
        oc8051_ram_top1_oc8051_idata_n1104) );
  OAI22_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2517 ( .A0(
        oc8051_ram_top1_oc8051_idata_n12), .A1(
        oc8051_ram_top1_oc8051_idata_n1109), .B0(
        oc8051_ram_top1_oc8051_idata_n4), .B1(
        oc8051_ram_top1_oc8051_idata_n1110), .Y(
        oc8051_ram_top1_oc8051_idata_n1108) );
  AOI221_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2516 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1106), .A1(
        oc8051_ram_top1_oc8051_idata_buff_3__7_), .B0(
        oc8051_ram_top1_oc8051_idata_n1107), .B1(
        oc8051_ram_top1_oc8051_idata_buff_2__7_), .C0(
        oc8051_ram_top1_oc8051_idata_n1108), .Y(
        oc8051_ram_top1_oc8051_idata_n1105) );
  NAND4_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2515 ( .A(
        oc8051_ram_top1_oc8051_idata_n1102), .B(
        oc8051_ram_top1_oc8051_idata_n1103), .C(
        oc8051_ram_top1_oc8051_idata_n1104), .D(
        oc8051_ram_top1_oc8051_idata_n1105), .Y(
        oc8051_ram_top1_oc8051_idata_n1101) );
  OR6_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2514 ( .A(
        oc8051_ram_top1_oc8051_idata_n1096), .B(
        oc8051_ram_top1_oc8051_idata_n1097), .C(
        oc8051_ram_top1_oc8051_idata_n1098), .D(
        oc8051_ram_top1_oc8051_idata_n1099), .E(
        oc8051_ram_top1_oc8051_idata_n1100), .F(
        oc8051_ram_top1_oc8051_idata_n1101), .Y(
        oc8051_ram_top1_oc8051_idata_n1095) );
  AOI222_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2513 ( .A0(
        oc8051_ram_top1_oc8051_idata_n1090), .A1(
        oc8051_ram_top1_oc8051_idata_n1091), .B0(
        oc8051_ram_top1_oc8051_idata_n1092), .B1(
        oc8051_ram_top1_oc8051_idata_n1093), .C0(
        oc8051_ram_top1_oc8051_idata_n1094), .C1(
        oc8051_ram_top1_oc8051_idata_n1095), .Y(
        oc8051_ram_top1_oc8051_idata_n1089) );
  OAI211_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2512 ( .A0(
        oc8051_ram_top1_oc8051_idata_n647), .A1(
        oc8051_ram_top1_oc8051_idata_n1087), .B0(
        oc8051_ram_top1_oc8051_idata_n1088), .C0(
        oc8051_ram_top1_oc8051_idata_n1089), .Y(
        oc8051_ram_top1_oc8051_idata_n2482) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2511 ( .A(wr_addr[7]), .B(
        n_0_net_), .Y(oc8051_ram_top1_oc8051_idata_n974) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2510 ( .A(
        oc8051_ram_top1_wr_addr_m_6_), .Y(oc8051_ram_top1_oc8051_idata_n872)
         );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2509 ( .AN(
        oc8051_ram_top1_oc8051_idata_n974), .B(
        oc8051_ram_top1_oc8051_idata_n872), .Y(
        oc8051_ram_top1_oc8051_idata_n992) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2508 ( .A(
        oc8051_ram_top1_wr_addr_m_4_), .Y(oc8051_ram_top1_oc8051_idata_n1010)
         );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2507 ( .AN(
        oc8051_ram_top1_wr_addr_m_5_), .B(oc8051_ram_top1_oc8051_idata_n1010), 
        .Y(oc8051_ram_top1_oc8051_idata_n769) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2506 ( .A(
        oc8051_ram_top1_oc8051_idata_n992), .B(
        oc8051_ram_top1_oc8051_idata_n769), .Y(
        oc8051_ram_top1_oc8051_idata_n1037) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2505 ( .A(
        oc8051_ram_top1_wr_addr_m_2_), .Y(oc8051_ram_top1_oc8051_idata_n1075)
         );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2504 ( .AN(
        oc8051_ram_top1_wr_addr_m_3_), .B(oc8051_ram_top1_oc8051_idata_n1075), 
        .Y(oc8051_ram_top1_oc8051_idata_n1082) );
  INV_X0P5B_A12TS oc8051_ram_top1_oc8051_idata_u2503 ( .A(
        oc8051_ram_top1_wr_addr_m_0_), .Y(oc8051_ram_top1_oc8051_idata_n1084)
         );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2502 ( .AN(
        oc8051_ram_top1_wr_addr_m_1_), .B(oc8051_ram_top1_oc8051_idata_n1084), 
        .Y(oc8051_ram_top1_oc8051_idata_n1053) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2501 ( .A(
        oc8051_ram_top1_oc8051_idata_n1082), .B(
        oc8051_ram_top1_oc8051_idata_n1053), .Y(
        oc8051_ram_top1_oc8051_idata_n681) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2500 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n1086) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2499 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2483) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2498 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2484) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2497 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2485) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2496 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2486) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2495 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2487) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2494 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2488) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2493 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2489) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2492 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_255__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1086), .Y(
        oc8051_ram_top1_oc8051_idata_n2490) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2491 ( .AN(
        oc8051_ram_top1_wr_addr_m_1_), .B(oc8051_ram_top1_wr_addr_m_0_), .Y(
        oc8051_ram_top1_oc8051_idata_n1051) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2490 ( .A(
        oc8051_ram_top1_oc8051_idata_n1082), .B(
        oc8051_ram_top1_oc8051_idata_n1051), .Y(
        oc8051_ram_top1_oc8051_idata_n679) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2489 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n1085) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2488 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2491) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2487 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2492) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2486 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2493) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2485 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2494) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2484 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2495) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2483 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2496) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2482 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2497) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2481 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_254__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1085), .Y(
        oc8051_ram_top1_oc8051_idata_n2498) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2480 ( .A(
        oc8051_ram_top1_oc8051_idata_n1084), .B(oc8051_ram_top1_wr_addr_m_1_), 
        .Y(oc8051_ram_top1_oc8051_idata_n1049) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2479 ( .A(
        oc8051_ram_top1_oc8051_idata_n1082), .B(
        oc8051_ram_top1_oc8051_idata_n1049), .Y(
        oc8051_ram_top1_oc8051_idata_n677) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2478 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n1083) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2477 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2499) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2476 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2500) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2475 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2501) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2474 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2502) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2473 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2503) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2472 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2504) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2471 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2505) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2470 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_253__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1083), .Y(
        oc8051_ram_top1_oc8051_idata_n2506) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2469 ( .A(
        oc8051_ram_top1_wr_addr_m_0_), .B(oc8051_ram_top1_wr_addr_m_1_), .Y(
        oc8051_ram_top1_oc8051_idata_n1039) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2468 ( .A(
        oc8051_ram_top1_oc8051_idata_n1082), .B(
        oc8051_ram_top1_oc8051_idata_n1039), .Y(
        oc8051_ram_top1_oc8051_idata_n675) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2467 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n1081) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2466 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2507) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2465 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2508) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2464 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2509) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2463 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2510) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2462 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2511) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2461 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2512) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2460 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2513) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2459 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_252__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1081), .Y(
        oc8051_ram_top1_oc8051_idata_n2514) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2458 ( .AN(
        oc8051_ram_top1_wr_addr_m_3_), .B(oc8051_ram_top1_wr_addr_m_2_), .Y(
        oc8051_ram_top1_oc8051_idata_n1077) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2457 ( .A(
        oc8051_ram_top1_oc8051_idata_n1077), .B(
        oc8051_ram_top1_oc8051_idata_n1053), .Y(
        oc8051_ram_top1_oc8051_idata_n673) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2456 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n1080) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2455 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2515) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2454 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2516) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2453 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2517) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2452 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2518) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2451 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2519) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2450 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2520) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2449 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2521) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2448 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_251__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1080), .Y(
        oc8051_ram_top1_oc8051_idata_n2522) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2447 ( .A(
        oc8051_ram_top1_oc8051_idata_n1077), .B(
        oc8051_ram_top1_oc8051_idata_n1051), .Y(
        oc8051_ram_top1_oc8051_idata_n671) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2446 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n1079) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2445 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2523) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2444 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2524) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2443 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2525) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2442 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2526) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2441 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2527) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2440 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2528) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2439 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2529) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2438 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_250__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1079), .Y(
        oc8051_ram_top1_oc8051_idata_n2530) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2437 ( .A(
        oc8051_ram_top1_oc8051_idata_n1077), .B(
        oc8051_ram_top1_oc8051_idata_n1049), .Y(
        oc8051_ram_top1_oc8051_idata_n669) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2436 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n1078) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2435 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2531) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2434 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2532) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2433 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2533) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2432 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2534) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2431 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2535) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2430 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2536) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2429 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2537) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2428 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_249__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1078), .Y(
        oc8051_ram_top1_oc8051_idata_n2538) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2427 ( .A(
        oc8051_ram_top1_oc8051_idata_n1077), .B(
        oc8051_ram_top1_oc8051_idata_n1039), .Y(
        oc8051_ram_top1_oc8051_idata_n667) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2426 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n1076) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2425 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2539) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2424 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2540) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2423 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2541) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2422 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2542) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2421 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2543) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2420 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2544) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2419 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2545) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2418 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_248__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1076), .Y(
        oc8051_ram_top1_oc8051_idata_n2546) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2417 ( .A(
        oc8051_ram_top1_oc8051_idata_n1075), .B(oc8051_ram_top1_wr_addr_m_3_), 
        .Y(oc8051_ram_top1_oc8051_idata_n1063) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2416 ( .A(
        oc8051_ram_top1_oc8051_idata_n1063), .B(
        oc8051_ram_top1_oc8051_idata_n1053), .Y(
        oc8051_ram_top1_oc8051_idata_n665) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2415 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n1074) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2414 ( .A(
        oc8051_ram_top1_oc8051_idata_n515), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2547) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2413 ( .A(
        oc8051_ram_top1_oc8051_idata_n514), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2548) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2412 ( .A(
        oc8051_ram_top1_oc8051_idata_n513), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2549) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2411 ( .A(
        oc8051_ram_top1_oc8051_idata_n512), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2550) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2410 ( .A(
        oc8051_ram_top1_oc8051_idata_n511), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2551) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2409 ( .A(
        oc8051_ram_top1_oc8051_idata_n510), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2552) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2408 ( .A(
        oc8051_ram_top1_oc8051_idata_n509), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2553) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2407 ( .A(
        oc8051_ram_top1_oc8051_idata_n508), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1074), .Y(
        oc8051_ram_top1_oc8051_idata_n2554) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2406 ( .A(
        oc8051_ram_top1_oc8051_idata_n1063), .B(
        oc8051_ram_top1_oc8051_idata_n1051), .Y(
        oc8051_ram_top1_oc8051_idata_n663) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2405 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n1073) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2404 ( .A(
        oc8051_ram_top1_oc8051_idata_n507), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2555) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2403 ( .A(
        oc8051_ram_top1_oc8051_idata_n506), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2556) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2402 ( .A(
        oc8051_ram_top1_oc8051_idata_n505), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2557) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2401 ( .A(
        oc8051_ram_top1_oc8051_idata_n504), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2558) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2400 ( .A(
        oc8051_ram_top1_oc8051_idata_n503), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2559) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2399 ( .A(
        oc8051_ram_top1_oc8051_idata_n502), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2560) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2398 ( .A(
        oc8051_ram_top1_oc8051_idata_n501), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2561) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2397 ( .A(
        oc8051_ram_top1_oc8051_idata_n500), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1073), .Y(
        oc8051_ram_top1_oc8051_idata_n2562) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2396 ( .A(
        oc8051_ram_top1_oc8051_idata_n1063), .B(
        oc8051_ram_top1_oc8051_idata_n1049), .Y(
        oc8051_ram_top1_oc8051_idata_n661) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2395 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n1065) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2394 ( .A(
        oc8051_ram_top1_oc8051_idata_n1072), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2563) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2393 ( .A(
        oc8051_ram_top1_oc8051_idata_n1071), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2564) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2392 ( .A(
        oc8051_ram_top1_oc8051_idata_n1070), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2565) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2391 ( .A(
        oc8051_ram_top1_oc8051_idata_n1069), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2566) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2390 ( .A(
        oc8051_ram_top1_oc8051_idata_n1068), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2567) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2389 ( .A(
        oc8051_ram_top1_oc8051_idata_n1067), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2568) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2388 ( .A(
        oc8051_ram_top1_oc8051_idata_n1066), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2569) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2387 ( .A(
        oc8051_ram_top1_oc8051_idata_n1064), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1065), .Y(
        oc8051_ram_top1_oc8051_idata_n2570) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2386 ( .A(
        oc8051_ram_top1_oc8051_idata_n1063), .B(
        oc8051_ram_top1_oc8051_idata_n1039), .Y(
        oc8051_ram_top1_oc8051_idata_n659) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2385 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n1055) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2384 ( .A(
        oc8051_ram_top1_oc8051_idata_n1062), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2571) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2383 ( .A(
        oc8051_ram_top1_oc8051_idata_n1061), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2572) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2382 ( .A(
        oc8051_ram_top1_oc8051_idata_n1060), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2573) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2381 ( .A(
        oc8051_ram_top1_oc8051_idata_n1059), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2574) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2380 ( .A(
        oc8051_ram_top1_oc8051_idata_n1058), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2575) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2379 ( .A(
        oc8051_ram_top1_oc8051_idata_n1057), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2576) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2378 ( .A(
        oc8051_ram_top1_oc8051_idata_n1056), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2577) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2377 ( .A(
        oc8051_ram_top1_oc8051_idata_n1054), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1055), .Y(
        oc8051_ram_top1_oc8051_idata_n2578) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2376 ( .A(
        oc8051_ram_top1_wr_addr_m_2_), .B(oc8051_ram_top1_wr_addr_m_3_), .Y(
        oc8051_ram_top1_oc8051_idata_n1038) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2375 ( .A(
        oc8051_ram_top1_oc8051_idata_n1053), .B(
        oc8051_ram_top1_oc8051_idata_n1038), .Y(
        oc8051_ram_top1_oc8051_idata_n657) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2374 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n1052) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2373 ( .A(
        oc8051_ram_top1_oc8051_idata_n499), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2579) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2372 ( .A(
        oc8051_ram_top1_oc8051_idata_n498), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2580) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2371 ( .A(
        oc8051_ram_top1_oc8051_idata_n497), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2581) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2370 ( .A(
        oc8051_ram_top1_oc8051_idata_n496), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2582) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2369 ( .A(
        oc8051_ram_top1_oc8051_idata_n495), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2583) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2368 ( .A(
        oc8051_ram_top1_oc8051_idata_n494), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2584) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2367 ( .A(
        oc8051_ram_top1_oc8051_idata_n493), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2585) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2366 ( .A(
        oc8051_ram_top1_oc8051_idata_n492), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1052), .Y(
        oc8051_ram_top1_oc8051_idata_n2586) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2365 ( .A(
        oc8051_ram_top1_oc8051_idata_n1051), .B(
        oc8051_ram_top1_oc8051_idata_n1038), .Y(
        oc8051_ram_top1_oc8051_idata_n655) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2364 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n1050) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2363 ( .A(
        oc8051_ram_top1_oc8051_idata_n491), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2587) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2362 ( .A(
        oc8051_ram_top1_oc8051_idata_n490), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2588) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2361 ( .A(
        oc8051_ram_top1_oc8051_idata_n489), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2589) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2360 ( .A(
        oc8051_ram_top1_oc8051_idata_n488), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2590) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2359 ( .A(
        oc8051_ram_top1_oc8051_idata_n487), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2591) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2358 ( .A(
        oc8051_ram_top1_oc8051_idata_n486), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2592) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2357 ( .A(
        oc8051_ram_top1_oc8051_idata_n485), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2593) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2356 ( .A(
        oc8051_ram_top1_oc8051_idata_n484), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1050), .Y(
        oc8051_ram_top1_oc8051_idata_n2594) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2355 ( .A(
        oc8051_ram_top1_oc8051_idata_n1049), .B(
        oc8051_ram_top1_oc8051_idata_n1038), .Y(
        oc8051_ram_top1_oc8051_idata_n653) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2354 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n1041) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2353 ( .A(
        oc8051_ram_top1_oc8051_idata_n1048), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2595) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2352 ( .A(
        oc8051_ram_top1_oc8051_idata_n1047), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2596) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2351 ( .A(
        oc8051_ram_top1_oc8051_idata_n1046), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2597) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2350 ( .A(
        oc8051_ram_top1_oc8051_idata_n1045), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2598) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2349 ( .A(
        oc8051_ram_top1_oc8051_idata_n1044), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2599) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2348 ( .A(
        oc8051_ram_top1_oc8051_idata_n1043), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2600) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2347 ( .A(
        oc8051_ram_top1_oc8051_idata_n1042), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2601) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2346 ( .A(
        oc8051_ram_top1_oc8051_idata_n1040), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1041), .Y(
        oc8051_ram_top1_oc8051_idata_n2602) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2345 ( .A(
        oc8051_ram_top1_oc8051_idata_n1038), .B(
        oc8051_ram_top1_oc8051_idata_n1039), .Y(
        oc8051_ram_top1_oc8051_idata_n650) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2344 ( .A(
        oc8051_ram_top1_oc8051_idata_n1037), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n1029) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2343 ( .A(
        oc8051_ram_top1_oc8051_idata_n1036), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2603) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2342 ( .A(
        oc8051_ram_top1_oc8051_idata_n1035), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2604) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2341 ( .A(
        oc8051_ram_top1_oc8051_idata_n1034), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2605) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2340 ( .A(
        oc8051_ram_top1_oc8051_idata_n1033), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2606) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2339 ( .A(
        oc8051_ram_top1_oc8051_idata_n1032), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2607) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2338 ( .A(
        oc8051_ram_top1_oc8051_idata_n1031), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2608) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2337 ( .A(
        oc8051_ram_top1_oc8051_idata_n1030), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2609) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2336 ( .A(
        oc8051_ram_top1_oc8051_idata_n1028), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1029), .Y(
        oc8051_ram_top1_oc8051_idata_n2610) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2335 ( .AN(
        oc8051_ram_top1_wr_addr_m_5_), .B(oc8051_ram_top1_wr_addr_m_4_), .Y(
        oc8051_ram_top1_oc8051_idata_n719) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2334 ( .A(
        oc8051_ram_top1_oc8051_idata_n992), .B(
        oc8051_ram_top1_oc8051_idata_n719), .Y(
        oc8051_ram_top1_oc8051_idata_n1012) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2333 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n1027) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2332 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2611) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2331 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2612) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2330 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2613) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2329 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2614) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2328 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2615) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2327 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2616) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2326 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2617) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2325 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_239__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1027), .Y(
        oc8051_ram_top1_oc8051_idata_n2618) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2324 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n1026) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2323 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2619) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2322 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2620) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2321 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2621) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2320 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2622) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2319 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2623) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2318 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2624) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2317 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2625) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2316 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_238__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1026), .Y(
        oc8051_ram_top1_oc8051_idata_n2626) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2315 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n1025) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2314 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2627) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2313 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2628) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2312 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2629) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2311 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2630) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2310 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2631) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2309 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2632) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2308 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2633) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2307 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_237__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1025), .Y(
        oc8051_ram_top1_oc8051_idata_n2634) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2306 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n1024) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2305 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2635) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2304 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2636) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2303 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2637) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2302 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2638) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2301 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2639) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2300 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2640) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2299 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2641) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2298 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_236__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n1024), .Y(
        oc8051_ram_top1_oc8051_idata_n2642) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2297 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n1023) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2296 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2643) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2295 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2644) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2294 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2645) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2293 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2646) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2292 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2647) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2291 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2648) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2290 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2649) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2289 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_235__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n1023), .Y(
        oc8051_ram_top1_oc8051_idata_n2650) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2288 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n1022) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2287 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2651) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2286 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2652) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2285 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2653) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2284 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2654) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2283 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2655) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2282 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2656) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2281 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2657) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2280 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_234__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n1022), .Y(
        oc8051_ram_top1_oc8051_idata_n2658) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2279 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n1021) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2278 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2659) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2277 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2660) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2276 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2661) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2275 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2662) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2274 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2663) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2273 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2664) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2272 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2665) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2271 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_233__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n1021), .Y(
        oc8051_ram_top1_oc8051_idata_n2666) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2270 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n1020) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2269 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2667) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2268 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2668) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2267 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2669) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2266 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2670) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2265 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2671) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2264 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2672) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2263 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2673) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2262 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_232__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n1020), .Y(
        oc8051_ram_top1_oc8051_idata_n2674) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2261 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n1019) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2260 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2675) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2259 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2676) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2258 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2677) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2257 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2678) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2256 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2679) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2255 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2680) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2254 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2681) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2253 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_231__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n1019), .Y(
        oc8051_ram_top1_oc8051_idata_n2682) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2252 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n1018) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2251 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2683) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2250 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2684) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2249 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2685) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2248 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2686) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2247 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2687) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2246 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2688) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2245 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2689) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2244 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_230__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n1018), .Y(
        oc8051_ram_top1_oc8051_idata_n2690) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2243 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n1017) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2242 ( .A(
        oc8051_ram_top1_oc8051_idata_n483), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2691) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2241 ( .A(
        oc8051_ram_top1_oc8051_idata_n482), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2692) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2240 ( .A(
        oc8051_ram_top1_oc8051_idata_n481), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2693) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2239 ( .A(
        oc8051_ram_top1_oc8051_idata_n480), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2694) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2238 ( .A(
        oc8051_ram_top1_oc8051_idata_n479), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2695) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2237 ( .A(
        oc8051_ram_top1_oc8051_idata_n478), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2696) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2236 ( .A(
        oc8051_ram_top1_oc8051_idata_n477), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2697) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2235 ( .A(
        oc8051_ram_top1_oc8051_idata_n476), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1017), .Y(
        oc8051_ram_top1_oc8051_idata_n2698) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2234 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n1016) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2233 ( .A(
        oc8051_ram_top1_oc8051_idata_n475), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2699) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2232 ( .A(
        oc8051_ram_top1_oc8051_idata_n474), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2700) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2231 ( .A(
        oc8051_ram_top1_oc8051_idata_n473), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2701) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2230 ( .A(
        oc8051_ram_top1_oc8051_idata_n472), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2702) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2229 ( .A(
        oc8051_ram_top1_oc8051_idata_n471), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2703) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2228 ( .A(
        oc8051_ram_top1_oc8051_idata_n470), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2704) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2227 ( .A(
        oc8051_ram_top1_oc8051_idata_n469), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2705) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2226 ( .A(
        oc8051_ram_top1_oc8051_idata_n468), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1016), .Y(
        oc8051_ram_top1_oc8051_idata_n2706) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2225 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n1015) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2224 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2707) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2223 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2708) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2222 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2709) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2221 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2710) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2220 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2711) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2219 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2712) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2218 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2713) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2217 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_227__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n1015), .Y(
        oc8051_ram_top1_oc8051_idata_n2714) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2216 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n1014) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2215 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2715) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2214 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2716) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2213 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2717) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2212 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2718) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2211 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2719) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2210 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2720) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2209 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2721) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2208 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_226__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n1014), .Y(
        oc8051_ram_top1_oc8051_idata_n2722) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2207 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n1013) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2206 ( .A(
        oc8051_ram_top1_oc8051_idata_n467), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2723) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2205 ( .A(
        oc8051_ram_top1_oc8051_idata_n466), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2724) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2204 ( .A(
        oc8051_ram_top1_oc8051_idata_n465), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2725) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2203 ( .A(
        oc8051_ram_top1_oc8051_idata_n464), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2726) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2202 ( .A(
        oc8051_ram_top1_oc8051_idata_n463), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2727) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2201 ( .A(
        oc8051_ram_top1_oc8051_idata_n462), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2728) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2200 ( .A(
        oc8051_ram_top1_oc8051_idata_n461), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2729) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2199 ( .A(
        oc8051_ram_top1_oc8051_idata_n460), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1013), .Y(
        oc8051_ram_top1_oc8051_idata_n2730) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2198 ( .A(
        oc8051_ram_top1_oc8051_idata_n1012), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n1011) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2197 ( .A(
        oc8051_ram_top1_oc8051_idata_n459), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2731) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2196 ( .A(
        oc8051_ram_top1_oc8051_idata_n458), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2732) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2195 ( .A(
        oc8051_ram_top1_oc8051_idata_n457), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2733) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2194 ( .A(
        oc8051_ram_top1_oc8051_idata_n456), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2734) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2193 ( .A(
        oc8051_ram_top1_oc8051_idata_n455), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2735) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2192 ( .A(
        oc8051_ram_top1_oc8051_idata_n454), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2736) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2191 ( .A(
        oc8051_ram_top1_oc8051_idata_n453), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2737) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2190 ( .A(
        oc8051_ram_top1_oc8051_idata_n452), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n1011), .Y(
        oc8051_ram_top1_oc8051_idata_n2738) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2189 ( .A(
        oc8051_ram_top1_oc8051_idata_n1010), .B(oc8051_ram_top1_wr_addr_m_5_), 
        .Y(oc8051_ram_top1_oc8051_idata_n701) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2188 ( .A(
        oc8051_ram_top1_oc8051_idata_n992), .B(
        oc8051_ram_top1_oc8051_idata_n701), .Y(
        oc8051_ram_top1_oc8051_idata_n994) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2187 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n1009) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2186 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2739) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2185 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2740) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2184 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2741) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2183 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2742) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2182 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2743) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2181 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2744) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2180 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2745) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2179 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_223__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n1009), .Y(
        oc8051_ram_top1_oc8051_idata_n2746) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2178 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n1008) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2177 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2747) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2176 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2748) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2175 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2749) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2174 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2750) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2173 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2751) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2172 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2752) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2171 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2753) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2170 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_222__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1008), .Y(
        oc8051_ram_top1_oc8051_idata_n2754) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2169 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n1007) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2168 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2755) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2167 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2756) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2166 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2757) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2165 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2758) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2164 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2759) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2163 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2760) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2162 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2761) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2161 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_221__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n1007), .Y(
        oc8051_ram_top1_oc8051_idata_n2762) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2160 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n1006) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2159 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2763) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2158 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2764) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2157 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2765) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2156 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2766) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2155 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2767) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2154 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2768) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2153 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2769) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2152 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_220__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n1006), .Y(
        oc8051_ram_top1_oc8051_idata_n2770) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2151 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n1005) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2150 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2771) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2149 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2772) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2148 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2773) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2147 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2774) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2146 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2775) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2145 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2776) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2144 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2777) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2143 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_219__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n1005), .Y(
        oc8051_ram_top1_oc8051_idata_n2778) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2142 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n1004) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2141 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2779) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2140 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2780) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2139 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2781) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2138 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2782) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2137 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2783) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2136 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2784) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2135 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2785) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2134 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_218__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n1004), .Y(
        oc8051_ram_top1_oc8051_idata_n2786) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2133 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n1003) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2132 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2787) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2131 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2788) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2130 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2789) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2129 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2790) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2128 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2791) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2127 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2792) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2126 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2793) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2125 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_217__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n1003), .Y(
        oc8051_ram_top1_oc8051_idata_n2794) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2124 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n1002) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2123 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2795) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2122 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2796) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2121 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2797) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2120 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2798) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2119 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2799) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2118 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2800) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2117 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2801) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2116 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_216__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n1002), .Y(
        oc8051_ram_top1_oc8051_idata_n2802) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2115 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n1001) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2114 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2803) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2113 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2804) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2112 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2805) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2111 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2806) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2110 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2807) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2109 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2808) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2108 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2809) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2107 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_215__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n1001), .Y(
        oc8051_ram_top1_oc8051_idata_n2810) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2106 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n1000) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2105 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2811) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2104 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2812) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2103 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2813) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2102 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2814) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2101 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2815) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2100 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2816) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2099 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2817) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2098 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_214__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n1000), .Y(
        oc8051_ram_top1_oc8051_idata_n2818) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2097 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n999) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2096 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2819) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2095 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2820) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2094 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2821) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2093 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2822) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2092 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2823) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2091 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2824) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2090 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2825) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2089 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_213__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n999), .Y(
        oc8051_ram_top1_oc8051_idata_n2826) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2088 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n998) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2087 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2827) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2086 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2828) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2085 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2829) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2084 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2830) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2083 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2831) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2082 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2832) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2081 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2833) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2080 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_212__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n998), .Y(
        oc8051_ram_top1_oc8051_idata_n2834) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2079 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n997) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2078 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2835) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2077 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2836) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2076 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2837) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2075 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2838) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2074 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2839) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2073 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2840) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2072 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2841) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2071 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_211__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n997), .Y(
        oc8051_ram_top1_oc8051_idata_n2842) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2070 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n996) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2069 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2843) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2068 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2844) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2067 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2845) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2066 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2846) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2065 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2847) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2064 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2848) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2063 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2849) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2062 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_210__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n996), .Y(
        oc8051_ram_top1_oc8051_idata_n2850) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2061 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n995) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2060 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2851) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2059 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2852) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2058 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2853) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2057 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2854) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2056 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2855) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2055 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2856) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2054 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2857) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2053 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_209__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n995), .Y(
        oc8051_ram_top1_oc8051_idata_n2858) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2052 ( .A(
        oc8051_ram_top1_oc8051_idata_n994), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n993) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2051 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2859) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2050 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2860) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2049 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2861) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2048 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2862) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2047 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2863) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2046 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2864) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2045 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2865) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2044 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_208__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n993), .Y(
        oc8051_ram_top1_oc8051_idata_n2866) );
  NOR2_X0P5A_A12TS oc8051_ram_top1_oc8051_idata_u2043 ( .A(
        oc8051_ram_top1_wr_addr_m_4_), .B(oc8051_ram_top1_wr_addr_m_5_), .Y(
        oc8051_ram_top1_oc8051_idata_n683) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2042 ( .A(
        oc8051_ram_top1_oc8051_idata_n992), .B(
        oc8051_ram_top1_oc8051_idata_n683), .Y(
        oc8051_ram_top1_oc8051_idata_n976) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2041 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n991) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2040 ( .A(
        oc8051_ram_top1_oc8051_idata_n451), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2867) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2039 ( .A(
        oc8051_ram_top1_oc8051_idata_n450), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2868) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2038 ( .A(
        oc8051_ram_top1_oc8051_idata_n449), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2869) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2037 ( .A(
        oc8051_ram_top1_oc8051_idata_n448), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2870) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2036 ( .A(
        oc8051_ram_top1_oc8051_idata_n447), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2871) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2035 ( .A(
        oc8051_ram_top1_oc8051_idata_n446), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2872) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2034 ( .A(
        oc8051_ram_top1_oc8051_idata_n445), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2873) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2033 ( .A(
        oc8051_ram_top1_oc8051_idata_n444), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n991), .Y(
        oc8051_ram_top1_oc8051_idata_n2874) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2032 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n990) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2031 ( .A(
        oc8051_ram_top1_oc8051_idata_n443), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2875) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2030 ( .A(
        oc8051_ram_top1_oc8051_idata_n442), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2876) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2029 ( .A(
        oc8051_ram_top1_oc8051_idata_n441), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2877) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2028 ( .A(
        oc8051_ram_top1_oc8051_idata_n440), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2878) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2027 ( .A(
        oc8051_ram_top1_oc8051_idata_n439), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2879) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2026 ( .A(
        oc8051_ram_top1_oc8051_idata_n438), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2880) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2025 ( .A(
        oc8051_ram_top1_oc8051_idata_n437), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2881) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2024 ( .A(
        oc8051_ram_top1_oc8051_idata_n436), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n990), .Y(
        oc8051_ram_top1_oc8051_idata_n2882) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2023 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n989) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2022 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2883) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2021 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2884) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2020 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2885) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2019 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2886) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2018 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2887) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2017 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2888) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2016 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2889) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2015 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_205__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n989), .Y(
        oc8051_ram_top1_oc8051_idata_n2890) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2014 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n988) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2013 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2891) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2012 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2892) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2011 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2893) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2010 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2894) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2009 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2895) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2008 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2896) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2007 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2897) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2006 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_204__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n988), .Y(
        oc8051_ram_top1_oc8051_idata_n2898) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2005 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n987) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2004 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2899) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2003 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2900) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2002 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2901) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2001 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2902) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u2000 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2903) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1999 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2904) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1998 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2905) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1997 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_203__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n987), .Y(
        oc8051_ram_top1_oc8051_idata_n2906) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1996 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n986) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1995 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2907) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1994 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2908) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1993 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2909) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1992 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2910) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1991 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2911) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1990 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2912) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1989 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2913) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1988 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_202__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n986), .Y(
        oc8051_ram_top1_oc8051_idata_n2914) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1987 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n985) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1986 ( .A(
        oc8051_ram_top1_oc8051_idata_n435), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2915) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1985 ( .A(
        oc8051_ram_top1_oc8051_idata_n434), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2916) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1984 ( .A(
        oc8051_ram_top1_oc8051_idata_n433), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2917) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1983 ( .A(
        oc8051_ram_top1_oc8051_idata_n432), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2918) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1982 ( .A(
        oc8051_ram_top1_oc8051_idata_n431), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2919) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1981 ( .A(
        oc8051_ram_top1_oc8051_idata_n430), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2920) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1980 ( .A(
        oc8051_ram_top1_oc8051_idata_n429), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2921) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1979 ( .A(
        oc8051_ram_top1_oc8051_idata_n428), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n985), .Y(
        oc8051_ram_top1_oc8051_idata_n2922) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1978 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n984) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1977 ( .A(
        oc8051_ram_top1_oc8051_idata_n427), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2923) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1976 ( .A(
        oc8051_ram_top1_oc8051_idata_n426), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2924) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1975 ( .A(
        oc8051_ram_top1_oc8051_idata_n425), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2925) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1974 ( .A(
        oc8051_ram_top1_oc8051_idata_n424), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2926) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1973 ( .A(
        oc8051_ram_top1_oc8051_idata_n423), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2927) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1972 ( .A(
        oc8051_ram_top1_oc8051_idata_n422), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2928) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1971 ( .A(
        oc8051_ram_top1_oc8051_idata_n421), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2929) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1970 ( .A(
        oc8051_ram_top1_oc8051_idata_n420), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n984), .Y(
        oc8051_ram_top1_oc8051_idata_n2930) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1969 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n983) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1968 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2931) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1967 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2932) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1966 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2933) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1965 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2934) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1964 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2935) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1963 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2936) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1962 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2937) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1961 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_199__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n983), .Y(
        oc8051_ram_top1_oc8051_idata_n2938) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1960 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n982) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1959 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2939) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1958 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2940) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1957 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2941) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1956 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2942) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1955 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2943) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1954 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2944) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1953 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2945) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1952 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_198__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n982), .Y(
        oc8051_ram_top1_oc8051_idata_n2946) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1951 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n981) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1950 ( .A(
        oc8051_ram_top1_oc8051_idata_n419), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2947) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1949 ( .A(
        oc8051_ram_top1_oc8051_idata_n418), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2948) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1948 ( .A(
        oc8051_ram_top1_oc8051_idata_n417), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2949) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1947 ( .A(
        oc8051_ram_top1_oc8051_idata_n416), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2950) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1946 ( .A(
        oc8051_ram_top1_oc8051_idata_n415), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2951) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1945 ( .A(
        oc8051_ram_top1_oc8051_idata_n414), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2952) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1944 ( .A(
        oc8051_ram_top1_oc8051_idata_n413), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2953) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1943 ( .A(
        oc8051_ram_top1_oc8051_idata_n412), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n981), .Y(
        oc8051_ram_top1_oc8051_idata_n2954) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1942 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n980) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1941 ( .A(
        oc8051_ram_top1_oc8051_idata_n411), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2955) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1940 ( .A(
        oc8051_ram_top1_oc8051_idata_n410), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2956) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1939 ( .A(
        oc8051_ram_top1_oc8051_idata_n409), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2957) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1938 ( .A(
        oc8051_ram_top1_oc8051_idata_n408), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2958) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1937 ( .A(
        oc8051_ram_top1_oc8051_idata_n407), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2959) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1936 ( .A(
        oc8051_ram_top1_oc8051_idata_n406), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2960) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1935 ( .A(
        oc8051_ram_top1_oc8051_idata_n405), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2961) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1934 ( .A(
        oc8051_ram_top1_oc8051_idata_n404), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n980), .Y(
        oc8051_ram_top1_oc8051_idata_n2962) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1933 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n979) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1932 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2963) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1931 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2964) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1930 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2965) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1929 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2966) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1928 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2967) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1927 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2968) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1926 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2969) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1925 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_195__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n979), .Y(
        oc8051_ram_top1_oc8051_idata_n2970) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1924 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n978) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1923 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2971) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1922 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2972) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1921 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2973) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1920 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2974) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1919 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2975) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1918 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2976) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1917 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2977) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1916 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_194__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n978), .Y(
        oc8051_ram_top1_oc8051_idata_n2978) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1915 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n977) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1914 ( .A(
        oc8051_ram_top1_oc8051_idata_n403), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2979) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1913 ( .A(
        oc8051_ram_top1_oc8051_idata_n402), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2980) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1912 ( .A(
        oc8051_ram_top1_oc8051_idata_n401), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2981) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1911 ( .A(
        oc8051_ram_top1_oc8051_idata_n400), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2982) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1910 ( .A(
        oc8051_ram_top1_oc8051_idata_n399), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2983) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1909 ( .A(
        oc8051_ram_top1_oc8051_idata_n398), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2984) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1908 ( .A(
        oc8051_ram_top1_oc8051_idata_n397), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2985) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1907 ( .A(
        oc8051_ram_top1_oc8051_idata_n396), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n977), .Y(
        oc8051_ram_top1_oc8051_idata_n2986) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1906 ( .A(
        oc8051_ram_top1_oc8051_idata_n976), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n975) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1905 ( .A(
        oc8051_ram_top1_oc8051_idata_n395), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2987) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1904 ( .A(
        oc8051_ram_top1_oc8051_idata_n394), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2988) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1903 ( .A(
        oc8051_ram_top1_oc8051_idata_n393), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2989) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1902 ( .A(
        oc8051_ram_top1_oc8051_idata_n392), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2990) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1901 ( .A(
        oc8051_ram_top1_oc8051_idata_n391), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2991) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1900 ( .A(
        oc8051_ram_top1_oc8051_idata_n390), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2992) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1899 ( .A(
        oc8051_ram_top1_oc8051_idata_n389), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2993) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1898 ( .A(
        oc8051_ram_top1_oc8051_idata_n388), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n975), .Y(
        oc8051_ram_top1_oc8051_idata_n2994) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1897 ( .AN(
        oc8051_ram_top1_oc8051_idata_n974), .B(oc8051_ram_top1_wr_addr_m_6_), 
        .Y(oc8051_ram_top1_oc8051_idata_n890) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1896 ( .A(
        oc8051_ram_top1_oc8051_idata_n890), .B(
        oc8051_ram_top1_oc8051_idata_n769), .Y(
        oc8051_ram_top1_oc8051_idata_n934) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1895 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n973) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1894 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n2995) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1893 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n2996) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1892 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n2997) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1891 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n2998) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1890 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n2999) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1889 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n3000) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1888 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n3001) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1887 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_191__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n973), .Y(
        oc8051_ram_top1_oc8051_idata_n3002) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1886 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n972) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1885 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3003) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1884 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3004) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1883 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3005) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1882 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3006) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1881 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3007) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1880 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3008) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1879 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3009) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1878 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_190__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n972), .Y(
        oc8051_ram_top1_oc8051_idata_n3010) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1877 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n971) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1876 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3011) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1875 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3012) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1874 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3013) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1873 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3014) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1872 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3015) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1871 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3016) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1870 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3017) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1869 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_189__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n971), .Y(
        oc8051_ram_top1_oc8051_idata_n3018) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1868 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n970) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1867 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3019) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1866 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3020) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1865 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3021) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1864 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3022) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1863 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3023) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1862 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3024) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1861 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3025) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1860 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_188__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n970), .Y(
        oc8051_ram_top1_oc8051_idata_n3026) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1859 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n969) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1858 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3027) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1857 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3028) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1856 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3029) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1855 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3030) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1854 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3031) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1853 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3032) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1852 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3033) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1851 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_187__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n969), .Y(
        oc8051_ram_top1_oc8051_idata_n3034) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1850 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n968) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1849 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3035) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1848 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3036) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1847 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3037) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1846 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3038) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1845 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3039) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1844 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3040) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1843 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3041) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1842 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_186__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n968), .Y(
        oc8051_ram_top1_oc8051_idata_n3042) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1841 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n967) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1840 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3043) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1839 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3044) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1838 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3045) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1837 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3046) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1836 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3047) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1835 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3048) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1834 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3049) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1833 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_185__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n967), .Y(
        oc8051_ram_top1_oc8051_idata_n3050) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1832 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n966) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1831 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3051) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1830 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3052) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1829 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3053) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1828 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3054) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1827 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3055) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1826 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3056) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1825 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3057) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1824 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_184__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n966), .Y(
        oc8051_ram_top1_oc8051_idata_n3058) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1823 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n965) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1822 ( .A(
        oc8051_ram_top1_oc8051_idata_n387), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3059) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1821 ( .A(
        oc8051_ram_top1_oc8051_idata_n386), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3060) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1820 ( .A(
        oc8051_ram_top1_oc8051_idata_n385), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3061) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1819 ( .A(
        oc8051_ram_top1_oc8051_idata_n384), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3062) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1818 ( .A(
        oc8051_ram_top1_oc8051_idata_n383), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3063) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1817 ( .A(
        oc8051_ram_top1_oc8051_idata_n382), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3064) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1816 ( .A(
        oc8051_ram_top1_oc8051_idata_n381), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3065) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1815 ( .A(
        oc8051_ram_top1_oc8051_idata_n380), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n965), .Y(
        oc8051_ram_top1_oc8051_idata_n3066) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1814 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n964) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1813 ( .A(
        oc8051_ram_top1_oc8051_idata_n379), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3067) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1812 ( .A(
        oc8051_ram_top1_oc8051_idata_n378), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3068) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1811 ( .A(
        oc8051_ram_top1_oc8051_idata_n377), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3069) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1810 ( .A(
        oc8051_ram_top1_oc8051_idata_n376), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3070) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1809 ( .A(
        oc8051_ram_top1_oc8051_idata_n375), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3071) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1808 ( .A(
        oc8051_ram_top1_oc8051_idata_n374), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3072) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1807 ( .A(
        oc8051_ram_top1_oc8051_idata_n373), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3073) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1806 ( .A(
        oc8051_ram_top1_oc8051_idata_n372), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n964), .Y(
        oc8051_ram_top1_oc8051_idata_n3074) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1805 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n956) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1804 ( .A(
        oc8051_ram_top1_oc8051_idata_n963), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3075) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1803 ( .A(
        oc8051_ram_top1_oc8051_idata_n962), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3076) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1802 ( .A(
        oc8051_ram_top1_oc8051_idata_n961), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3077) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1801 ( .A(
        oc8051_ram_top1_oc8051_idata_n960), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3078) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1800 ( .A(
        oc8051_ram_top1_oc8051_idata_n959), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3079) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1799 ( .A(
        oc8051_ram_top1_oc8051_idata_n958), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3080) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1798 ( .A(
        oc8051_ram_top1_oc8051_idata_n957), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3081) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1797 ( .A(
        oc8051_ram_top1_oc8051_idata_n955), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n956), .Y(
        oc8051_ram_top1_oc8051_idata_n3082) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1796 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n947) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1795 ( .A(
        oc8051_ram_top1_oc8051_idata_n954), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3083) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1794 ( .A(
        oc8051_ram_top1_oc8051_idata_n953), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3084) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1793 ( .A(
        oc8051_ram_top1_oc8051_idata_n952), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3085) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1792 ( .A(
        oc8051_ram_top1_oc8051_idata_n951), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3086) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1791 ( .A(
        oc8051_ram_top1_oc8051_idata_n950), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3087) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1790 ( .A(
        oc8051_ram_top1_oc8051_idata_n949), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3088) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1789 ( .A(
        oc8051_ram_top1_oc8051_idata_n948), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3089) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1788 ( .A(
        oc8051_ram_top1_oc8051_idata_n946), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n947), .Y(
        oc8051_ram_top1_oc8051_idata_n3090) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1787 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n945) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1786 ( .A(
        oc8051_ram_top1_oc8051_idata_n371), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3091) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1785 ( .A(
        oc8051_ram_top1_oc8051_idata_n370), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3092) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1784 ( .A(
        oc8051_ram_top1_oc8051_idata_n369), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3093) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1783 ( .A(
        oc8051_ram_top1_oc8051_idata_n368), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3094) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1782 ( .A(
        oc8051_ram_top1_oc8051_idata_n367), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3095) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1781 ( .A(
        oc8051_ram_top1_oc8051_idata_n366), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3096) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1780 ( .A(
        oc8051_ram_top1_oc8051_idata_n365), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3097) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1779 ( .A(
        oc8051_ram_top1_oc8051_idata_n364), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n945), .Y(
        oc8051_ram_top1_oc8051_idata_n3098) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1778 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n944) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1777 ( .A(
        oc8051_ram_top1_oc8051_idata_n363), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3099) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1776 ( .A(
        oc8051_ram_top1_oc8051_idata_n362), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3100) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1775 ( .A(
        oc8051_ram_top1_oc8051_idata_n361), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3101) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1774 ( .A(
        oc8051_ram_top1_oc8051_idata_n360), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3102) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1773 ( .A(
        oc8051_ram_top1_oc8051_idata_n359), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3103) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1772 ( .A(
        oc8051_ram_top1_oc8051_idata_n358), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3104) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1771 ( .A(
        oc8051_ram_top1_oc8051_idata_n357), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3105) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1770 ( .A(
        oc8051_ram_top1_oc8051_idata_n356), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n944), .Y(
        oc8051_ram_top1_oc8051_idata_n3106) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1769 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n936) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1768 ( .A(
        oc8051_ram_top1_oc8051_idata_n943), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3107) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1767 ( .A(
        oc8051_ram_top1_oc8051_idata_n942), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3108) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1766 ( .A(
        oc8051_ram_top1_oc8051_idata_n941), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3109) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1765 ( .A(
        oc8051_ram_top1_oc8051_idata_n940), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3110) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1764 ( .A(
        oc8051_ram_top1_oc8051_idata_n939), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3111) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1763 ( .A(
        oc8051_ram_top1_oc8051_idata_n938), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3112) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1762 ( .A(
        oc8051_ram_top1_oc8051_idata_n937), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3113) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1761 ( .A(
        oc8051_ram_top1_oc8051_idata_n935), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n936), .Y(
        oc8051_ram_top1_oc8051_idata_n3114) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1760 ( .A(
        oc8051_ram_top1_oc8051_idata_n934), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n926) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1759 ( .A(
        oc8051_ram_top1_oc8051_idata_n933), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3115) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1758 ( .A(
        oc8051_ram_top1_oc8051_idata_n932), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3116) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1757 ( .A(
        oc8051_ram_top1_oc8051_idata_n931), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3117) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1756 ( .A(
        oc8051_ram_top1_oc8051_idata_n930), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3118) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1755 ( .A(
        oc8051_ram_top1_oc8051_idata_n929), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3119) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1754 ( .A(
        oc8051_ram_top1_oc8051_idata_n928), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3120) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1753 ( .A(
        oc8051_ram_top1_oc8051_idata_n927), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3121) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1752 ( .A(
        oc8051_ram_top1_oc8051_idata_n925), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n926), .Y(
        oc8051_ram_top1_oc8051_idata_n3122) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1751 ( .A(
        oc8051_ram_top1_oc8051_idata_n890), .B(
        oc8051_ram_top1_oc8051_idata_n719), .Y(
        oc8051_ram_top1_oc8051_idata_n909) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1750 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n924) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1749 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3123) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1748 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3124) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1747 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3125) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1746 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3126) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1745 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3127) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1744 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3128) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1743 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3129) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1742 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_175__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n924), .Y(
        oc8051_ram_top1_oc8051_idata_n3130) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1741 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n923) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1740 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3131) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1739 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3132) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1738 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3133) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1737 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3134) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1736 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3135) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1735 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3136) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1734 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3137) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1733 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_174__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n923), .Y(
        oc8051_ram_top1_oc8051_idata_n3138) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1732 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n922) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1731 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3139) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1730 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3140) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1729 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3141) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1728 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3142) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1727 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3143) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1726 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3144) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1725 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3145) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1724 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_173__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n922), .Y(
        oc8051_ram_top1_oc8051_idata_n3146) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1723 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n921) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1722 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3147) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1721 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3148) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1720 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3149) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1719 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3150) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1718 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3151) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1717 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3152) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1716 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3153) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1715 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_172__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n921), .Y(
        oc8051_ram_top1_oc8051_idata_n3154) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1714 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n920) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1713 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3155) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1712 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3156) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1711 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3157) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1710 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3158) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1709 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3159) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1708 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3160) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1707 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3161) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1706 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_171__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n920), .Y(
        oc8051_ram_top1_oc8051_idata_n3162) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1705 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n919) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1704 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3163) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1703 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3164) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1702 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3165) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1701 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3166) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1700 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3167) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1699 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3168) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1698 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3169) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1697 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_170__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n919), .Y(
        oc8051_ram_top1_oc8051_idata_n3170) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1696 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n918) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1695 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3171) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1694 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3172) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1693 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3173) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1692 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3174) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1691 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3175) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1690 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3176) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1689 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3177) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1688 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_169__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n918), .Y(
        oc8051_ram_top1_oc8051_idata_n3178) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1687 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n917) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1686 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3179) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1685 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3180) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1684 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3181) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1683 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3182) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1682 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3183) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1681 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3184) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1680 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3185) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1679 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_168__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n917), .Y(
        oc8051_ram_top1_oc8051_idata_n3186) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1678 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n916) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1677 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3187) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1676 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3188) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1675 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3189) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1674 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3190) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1673 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3191) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1672 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3192) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1671 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3193) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1670 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_167__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n916), .Y(
        oc8051_ram_top1_oc8051_idata_n3194) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1669 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n915) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1668 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3195) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1667 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3196) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1666 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3197) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1665 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3198) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1664 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3199) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1663 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3200) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1662 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3201) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1661 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_166__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n915), .Y(
        oc8051_ram_top1_oc8051_idata_n3202) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1660 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n914) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1659 ( .A(
        oc8051_ram_top1_oc8051_idata_n355), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3203) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1658 ( .A(
        oc8051_ram_top1_oc8051_idata_n354), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3204) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1657 ( .A(
        oc8051_ram_top1_oc8051_idata_n353), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3205) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1656 ( .A(
        oc8051_ram_top1_oc8051_idata_n352), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3206) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1655 ( .A(
        oc8051_ram_top1_oc8051_idata_n351), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3207) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1654 ( .A(
        oc8051_ram_top1_oc8051_idata_n350), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3208) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1653 ( .A(
        oc8051_ram_top1_oc8051_idata_n349), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3209) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1652 ( .A(
        oc8051_ram_top1_oc8051_idata_n348), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n914), .Y(
        oc8051_ram_top1_oc8051_idata_n3210) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1651 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n913) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1650 ( .A(
        oc8051_ram_top1_oc8051_idata_n347), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3211) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1649 ( .A(
        oc8051_ram_top1_oc8051_idata_n346), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3212) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1648 ( .A(
        oc8051_ram_top1_oc8051_idata_n345), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3213) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1647 ( .A(
        oc8051_ram_top1_oc8051_idata_n344), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3214) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1646 ( .A(
        oc8051_ram_top1_oc8051_idata_n343), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3215) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1645 ( .A(
        oc8051_ram_top1_oc8051_idata_n342), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3216) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1644 ( .A(
        oc8051_ram_top1_oc8051_idata_n341), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3217) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1643 ( .A(
        oc8051_ram_top1_oc8051_idata_n340), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n913), .Y(
        oc8051_ram_top1_oc8051_idata_n3218) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1642 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n912) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1641 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3219) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1640 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3220) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1639 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3221) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1638 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3222) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1637 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3223) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1636 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3224) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1635 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3225) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1634 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_163__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n912), .Y(
        oc8051_ram_top1_oc8051_idata_n3226) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1633 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n911) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1632 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3227) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1631 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3228) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1630 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3229) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1629 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3230) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1628 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3231) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1627 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3232) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1626 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3233) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1625 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_162__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n911), .Y(
        oc8051_ram_top1_oc8051_idata_n3234) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1624 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n910) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1623 ( .A(
        oc8051_ram_top1_oc8051_idata_n339), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3235) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1622 ( .A(
        oc8051_ram_top1_oc8051_idata_n338), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3236) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1621 ( .A(
        oc8051_ram_top1_oc8051_idata_n337), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3237) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1620 ( .A(
        oc8051_ram_top1_oc8051_idata_n336), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3238) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1619 ( .A(
        oc8051_ram_top1_oc8051_idata_n335), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3239) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1618 ( .A(
        oc8051_ram_top1_oc8051_idata_n334), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3240) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1617 ( .A(
        oc8051_ram_top1_oc8051_idata_n333), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3241) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1616 ( .A(
        oc8051_ram_top1_oc8051_idata_n332), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n910), .Y(
        oc8051_ram_top1_oc8051_idata_n3242) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1615 ( .A(
        oc8051_ram_top1_oc8051_idata_n909), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n908) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1614 ( .A(
        oc8051_ram_top1_oc8051_idata_n331), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3243) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1613 ( .A(
        oc8051_ram_top1_oc8051_idata_n330), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3244) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1612 ( .A(
        oc8051_ram_top1_oc8051_idata_n329), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3245) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1611 ( .A(
        oc8051_ram_top1_oc8051_idata_n328), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3246) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1610 ( .A(
        oc8051_ram_top1_oc8051_idata_n327), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3247) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1609 ( .A(
        oc8051_ram_top1_oc8051_idata_n326), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3248) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1608 ( .A(
        oc8051_ram_top1_oc8051_idata_n325), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3249) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1607 ( .A(
        oc8051_ram_top1_oc8051_idata_n324), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n908), .Y(
        oc8051_ram_top1_oc8051_idata_n3250) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1606 ( .A(
        oc8051_ram_top1_oc8051_idata_n890), .B(
        oc8051_ram_top1_oc8051_idata_n701), .Y(
        oc8051_ram_top1_oc8051_idata_n892) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1605 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n907) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1604 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3251) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1603 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3252) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1602 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3253) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1601 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3254) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1600 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3255) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1599 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3256) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1598 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3257) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1597 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_159__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n907), .Y(
        oc8051_ram_top1_oc8051_idata_n3258) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1596 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n906) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1595 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3259) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1594 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3260) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1593 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3261) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1592 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3262) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1591 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3263) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1590 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3264) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1589 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3265) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1588 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_158__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n906), .Y(
        oc8051_ram_top1_oc8051_idata_n3266) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1587 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n905) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1586 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3267) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1585 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3268) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1584 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3269) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1583 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3270) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1582 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3271) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1581 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3272) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1580 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3273) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1579 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_157__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n905), .Y(
        oc8051_ram_top1_oc8051_idata_n3274) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1578 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n904) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1577 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__0_), .B(
        oc8051_ram_top1_oc8051_idata_n522), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3275) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1576 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__1_), .B(
        oc8051_ram_top1_oc8051_idata_n539), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3276) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1575 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__2_), .B(
        oc8051_ram_top1_oc8051_idata_n556), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3277) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1574 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__3_), .B(
        oc8051_ram_top1_oc8051_idata_n573), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3278) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1573 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__4_), .B(
        oc8051_ram_top1_oc8051_idata_n590), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3279) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1572 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__5_), .B(
        oc8051_ram_top1_oc8051_idata_n607), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3280) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1571 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__6_), .B(
        oc8051_ram_top1_oc8051_idata_n624), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3281) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1570 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_156__7_), .B(
        oc8051_ram_top1_oc8051_idata_n641), .S0(
        oc8051_ram_top1_oc8051_idata_n904), .Y(
        oc8051_ram_top1_oc8051_idata_n3282) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1569 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n903) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1568 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__0_), .B(
        oc8051_ram_top1_oc8051_idata_n521), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3283) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1567 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__1_), .B(
        oc8051_ram_top1_oc8051_idata_n538), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3284) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1566 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__2_), .B(
        oc8051_ram_top1_oc8051_idata_n555), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3285) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1565 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__3_), .B(
        oc8051_ram_top1_oc8051_idata_n572), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3286) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1564 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__4_), .B(
        oc8051_ram_top1_oc8051_idata_n589), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3287) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1563 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__5_), .B(
        oc8051_ram_top1_oc8051_idata_n606), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3288) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1562 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__6_), .B(
        oc8051_ram_top1_oc8051_idata_n623), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3289) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1561 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_155__7_), .B(
        oc8051_ram_top1_oc8051_idata_n640), .S0(
        oc8051_ram_top1_oc8051_idata_n903), .Y(
        oc8051_ram_top1_oc8051_idata_n3290) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1560 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n902) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1559 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__0_), .B(oc8051_ram_top1_n1), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3291) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1558 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__1_), .B(oc8051_ram_top1_n2), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3292) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1557 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__2_), .B(oc8051_ram_top1_n3), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3293) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1556 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__3_), .B(oc8051_ram_top1_n4), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3294) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1555 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__4_), .B(oc8051_ram_top1_n5), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3295) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1554 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__5_), .B(oc8051_ram_top1_n6), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3296) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1553 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__6_), .B(oc8051_ram_top1_n7), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3297) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1552 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_154__7_), .B(oc8051_ram_top1_n8), 
        .S0(oc8051_ram_top1_oc8051_idata_n902), .Y(
        oc8051_ram_top1_oc8051_idata_n3298) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1551 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n901) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1550 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3299) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1549 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3300) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1548 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3301) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1547 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3302) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1546 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3303) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1545 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3304) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1544 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3305) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1543 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_153__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n901), .Y(
        oc8051_ram_top1_oc8051_idata_n3306) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1542 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n900) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1541 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3307) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1540 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3308) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1539 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3309) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1538 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3310) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1537 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3311) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1536 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3312) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1535 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3313) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1534 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_152__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n900), .Y(
        oc8051_ram_top1_oc8051_idata_n3314) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1533 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n899) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1532 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3315) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1531 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3316) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1530 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3317) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1529 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3318) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1528 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3319) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1527 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3320) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1526 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3321) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1525 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_151__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n899), .Y(
        oc8051_ram_top1_oc8051_idata_n3322) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1524 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n898) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1523 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3323) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1522 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3324) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1521 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3325) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1520 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3326) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1519 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3327) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1518 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3328) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1517 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3329) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1516 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_150__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n898), .Y(
        oc8051_ram_top1_oc8051_idata_n3330) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1515 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n897) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1514 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3331) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1513 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3332) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1512 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3333) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1511 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3334) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1510 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3335) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1509 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3336) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1508 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3337) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1507 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_149__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n897), .Y(
        oc8051_ram_top1_oc8051_idata_n3338) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1506 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n896) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1505 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3339) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1504 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3340) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1503 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3341) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1502 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3342) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1501 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3343) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1500 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3344) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1499 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3345) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1498 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_148__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n896), .Y(
        oc8051_ram_top1_oc8051_idata_n3346) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1497 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n895) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1496 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3347) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1495 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3348) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1494 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3349) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1493 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3350) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1492 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3351) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1491 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3352) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1490 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3353) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1489 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_147__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n895), .Y(
        oc8051_ram_top1_oc8051_idata_n3354) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1488 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n894) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1487 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3355) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1486 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3356) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1485 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3357) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1484 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3358) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1483 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3359) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1482 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3360) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1481 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3361) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1480 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_146__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n894), .Y(
        oc8051_ram_top1_oc8051_idata_n3362) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1479 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n893) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1478 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3363) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1477 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3364) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1476 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3365) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1475 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3366) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1474 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3367) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1473 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3368) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1472 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3369) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1471 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_145__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n893), .Y(
        oc8051_ram_top1_oc8051_idata_n3370) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1470 ( .A(
        oc8051_ram_top1_oc8051_idata_n892), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n891) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1469 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3371) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1468 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3372) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1467 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3373) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1466 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3374) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1465 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3375) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1464 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3376) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1463 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3377) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1462 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_144__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n891), .Y(
        oc8051_ram_top1_oc8051_idata_n3378) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1461 ( .A(
        oc8051_ram_top1_oc8051_idata_n890), .B(
        oc8051_ram_top1_oc8051_idata_n683), .Y(
        oc8051_ram_top1_oc8051_idata_n874) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1460 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n889) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1459 ( .A(
        oc8051_ram_top1_oc8051_idata_n323), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3379) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1458 ( .A(
        oc8051_ram_top1_oc8051_idata_n322), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3380) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1457 ( .A(
        oc8051_ram_top1_oc8051_idata_n321), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3381) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1456 ( .A(
        oc8051_ram_top1_oc8051_idata_n320), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3382) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1455 ( .A(
        oc8051_ram_top1_oc8051_idata_n319), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3383) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1454 ( .A(
        oc8051_ram_top1_oc8051_idata_n318), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3384) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1453 ( .A(
        oc8051_ram_top1_oc8051_idata_n317), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3385) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1452 ( .A(
        oc8051_ram_top1_oc8051_idata_n316), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n889), .Y(
        oc8051_ram_top1_oc8051_idata_n3386) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1451 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n888) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1450 ( .A(
        oc8051_ram_top1_oc8051_idata_n315), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3387) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1449 ( .A(
        oc8051_ram_top1_oc8051_idata_n314), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3388) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1448 ( .A(
        oc8051_ram_top1_oc8051_idata_n313), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3389) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1447 ( .A(
        oc8051_ram_top1_oc8051_idata_n312), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3390) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1446 ( .A(
        oc8051_ram_top1_oc8051_idata_n311), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3391) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1445 ( .A(
        oc8051_ram_top1_oc8051_idata_n310), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3392) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1444 ( .A(
        oc8051_ram_top1_oc8051_idata_n309), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3393) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1443 ( .A(
        oc8051_ram_top1_oc8051_idata_n308), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n888), .Y(
        oc8051_ram_top1_oc8051_idata_n3394) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1442 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n887) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1441 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3395) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1440 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3396) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1439 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3397) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1438 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3398) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1437 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3399) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1436 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3400) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1435 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3401) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1434 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_141__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n887), .Y(
        oc8051_ram_top1_oc8051_idata_n3402) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1433 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n886) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1432 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3403) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1431 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3404) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1430 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3405) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1429 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3406) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1428 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3407) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1427 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3408) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1426 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3409) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1425 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_140__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n886), .Y(
        oc8051_ram_top1_oc8051_idata_n3410) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1424 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n885) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1423 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3411) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1422 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3412) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1421 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3413) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1420 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3414) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1419 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3415) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1418 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3416) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1417 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3417) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1416 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_139__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n885), .Y(
        oc8051_ram_top1_oc8051_idata_n3418) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1415 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n884) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1414 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3419) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1413 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3420) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1412 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3421) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1411 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3422) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1410 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3423) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1409 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3424) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1408 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3425) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1407 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_138__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n884), .Y(
        oc8051_ram_top1_oc8051_idata_n3426) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1406 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n883) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1405 ( .A(
        oc8051_ram_top1_oc8051_idata_n307), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3427) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1404 ( .A(
        oc8051_ram_top1_oc8051_idata_n306), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3428) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1403 ( .A(
        oc8051_ram_top1_oc8051_idata_n305), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3429) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1402 ( .A(
        oc8051_ram_top1_oc8051_idata_n304), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3430) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1401 ( .A(
        oc8051_ram_top1_oc8051_idata_n303), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3431) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1400 ( .A(
        oc8051_ram_top1_oc8051_idata_n302), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3432) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1399 ( .A(
        oc8051_ram_top1_oc8051_idata_n301), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3433) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1398 ( .A(
        oc8051_ram_top1_oc8051_idata_n300), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n883), .Y(
        oc8051_ram_top1_oc8051_idata_n3434) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1397 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n882) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1396 ( .A(
        oc8051_ram_top1_oc8051_idata_n299), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3435) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1395 ( .A(
        oc8051_ram_top1_oc8051_idata_n298), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3436) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1394 ( .A(
        oc8051_ram_top1_oc8051_idata_n297), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3437) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1393 ( .A(
        oc8051_ram_top1_oc8051_idata_n296), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3438) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1392 ( .A(
        oc8051_ram_top1_oc8051_idata_n295), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3439) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1391 ( .A(
        oc8051_ram_top1_oc8051_idata_n294), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3440) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1390 ( .A(
        oc8051_ram_top1_oc8051_idata_n293), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3441) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1389 ( .A(
        oc8051_ram_top1_oc8051_idata_n292), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n882), .Y(
        oc8051_ram_top1_oc8051_idata_n3442) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1388 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n881) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1387 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__0_), .B(
        oc8051_ram_top1_oc8051_idata_n520), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3443) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1386 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__1_), .B(
        oc8051_ram_top1_oc8051_idata_n537), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3444) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1385 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__2_), .B(
        oc8051_ram_top1_oc8051_idata_n554), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3445) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1384 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__3_), .B(
        oc8051_ram_top1_oc8051_idata_n571), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3446) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1383 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__4_), .B(
        oc8051_ram_top1_oc8051_idata_n588), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3447) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1382 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__5_), .B(
        oc8051_ram_top1_oc8051_idata_n605), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3448) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1381 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__6_), .B(
        oc8051_ram_top1_oc8051_idata_n622), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3449) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1380 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_135__7_), .B(
        oc8051_ram_top1_oc8051_idata_n639), .S0(
        oc8051_ram_top1_oc8051_idata_n881), .Y(
        oc8051_ram_top1_oc8051_idata_n3450) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1379 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n880) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1378 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3451) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1377 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3452) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1376 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3453) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1375 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3454) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1374 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3455) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1373 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3456) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1372 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3457) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1371 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_134__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n880), .Y(
        oc8051_ram_top1_oc8051_idata_n3458) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1370 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n879) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1369 ( .A(
        oc8051_ram_top1_oc8051_idata_n291), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3459) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1368 ( .A(
        oc8051_ram_top1_oc8051_idata_n290), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3460) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1367 ( .A(
        oc8051_ram_top1_oc8051_idata_n289), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3461) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1366 ( .A(
        oc8051_ram_top1_oc8051_idata_n288), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3462) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1365 ( .A(
        oc8051_ram_top1_oc8051_idata_n287), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3463) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1364 ( .A(
        oc8051_ram_top1_oc8051_idata_n286), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3464) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1363 ( .A(
        oc8051_ram_top1_oc8051_idata_n285), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3465) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1362 ( .A(
        oc8051_ram_top1_oc8051_idata_n284), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n879), .Y(
        oc8051_ram_top1_oc8051_idata_n3466) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1361 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n878) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1360 ( .A(
        oc8051_ram_top1_oc8051_idata_n283), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3467) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1359 ( .A(
        oc8051_ram_top1_oc8051_idata_n282), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3468) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1358 ( .A(
        oc8051_ram_top1_oc8051_idata_n281), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3469) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1357 ( .A(
        oc8051_ram_top1_oc8051_idata_n280), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3470) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1356 ( .A(
        oc8051_ram_top1_oc8051_idata_n279), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3471) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1355 ( .A(
        oc8051_ram_top1_oc8051_idata_n278), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3472) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1354 ( .A(
        oc8051_ram_top1_oc8051_idata_n277), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3473) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1353 ( .A(
        oc8051_ram_top1_oc8051_idata_n276), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n878), .Y(
        oc8051_ram_top1_oc8051_idata_n3474) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1352 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n877) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1351 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3475) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1350 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3476) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1349 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3477) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1348 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3478) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1347 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3479) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1346 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3480) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1345 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3481) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1344 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_131__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n877), .Y(
        oc8051_ram_top1_oc8051_idata_n3482) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1343 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n876) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1342 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3483) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1341 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3484) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1340 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3485) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1339 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3486) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1338 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3487) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1337 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3488) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1336 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3489) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1335 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_130__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n876), .Y(
        oc8051_ram_top1_oc8051_idata_n3490) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1334 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n875) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1333 ( .A(
        oc8051_ram_top1_oc8051_idata_n275), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3491) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1332 ( .A(
        oc8051_ram_top1_oc8051_idata_n274), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3492) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1331 ( .A(
        oc8051_ram_top1_oc8051_idata_n273), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3493) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1330 ( .A(
        oc8051_ram_top1_oc8051_idata_n272), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3494) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1329 ( .A(
        oc8051_ram_top1_oc8051_idata_n271), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3495) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1328 ( .A(
        oc8051_ram_top1_oc8051_idata_n270), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3496) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1327 ( .A(
        oc8051_ram_top1_oc8051_idata_n269), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3497) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1326 ( .A(
        oc8051_ram_top1_oc8051_idata_n268), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n875), .Y(
        oc8051_ram_top1_oc8051_idata_n3498) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1325 ( .A(
        oc8051_ram_top1_oc8051_idata_n874), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n873) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1324 ( .A(
        oc8051_ram_top1_oc8051_idata_n267), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3499) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1323 ( .A(
        oc8051_ram_top1_oc8051_idata_n266), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3500) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1322 ( .A(
        oc8051_ram_top1_oc8051_idata_n265), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3501) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1321 ( .A(
        oc8051_ram_top1_oc8051_idata_n264), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3502) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1320 ( .A(
        oc8051_ram_top1_oc8051_idata_n263), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3503) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1319 ( .A(
        oc8051_ram_top1_oc8051_idata_n262), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3504) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1318 ( .A(
        oc8051_ram_top1_oc8051_idata_n261), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3505) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1317 ( .A(
        oc8051_ram_top1_oc8051_idata_n260), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n873), .Y(
        oc8051_ram_top1_oc8051_idata_n3506) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1316 ( .AN(n_0_net_), .B(
        wr_addr[7]), .Y(oc8051_ram_top1_oc8051_idata_n770) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1315 ( .AN(
        oc8051_ram_top1_oc8051_idata_n770), .B(
        oc8051_ram_top1_oc8051_idata_n872), .Y(
        oc8051_ram_top1_oc8051_idata_n788) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1314 ( .A(
        oc8051_ram_top1_oc8051_idata_n788), .B(
        oc8051_ram_top1_oc8051_idata_n769), .Y(
        oc8051_ram_top1_oc8051_idata_n832) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1313 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n871) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1312 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3507) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1311 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3508) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1310 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3509) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1309 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3510) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1308 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3511) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1307 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3512) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1306 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3513) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1305 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_127__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n871), .Y(
        oc8051_ram_top1_oc8051_idata_n3514) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1304 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n870) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1303 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3515) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1302 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3516) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1301 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3517) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1300 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3518) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1299 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3519) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1298 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3520) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1297 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3521) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1296 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_126__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n870), .Y(
        oc8051_ram_top1_oc8051_idata_n3522) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1295 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n869) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1294 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3523) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1293 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3524) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1292 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3525) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1291 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3526) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1290 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3527) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1289 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3528) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1288 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3529) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1287 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_125__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n869), .Y(
        oc8051_ram_top1_oc8051_idata_n3530) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1286 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n868) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1285 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3531) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1284 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3532) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1283 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3533) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1282 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3534) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1281 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3535) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1280 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3536) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1279 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3537) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1278 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_124__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n868), .Y(
        oc8051_ram_top1_oc8051_idata_n3538) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1277 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n867) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1276 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3539) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1275 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3540) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1274 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3541) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1273 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3542) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1272 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3543) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1271 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3544) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1270 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3545) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1269 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_123__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n867), .Y(
        oc8051_ram_top1_oc8051_idata_n3546) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1268 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n866) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1267 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3547) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1266 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3548) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1265 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3549) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1264 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3550) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1263 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3551) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1262 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3552) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1261 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3553) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1260 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_122__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n866), .Y(
        oc8051_ram_top1_oc8051_idata_n3554) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1259 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n865) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1258 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3555) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1257 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3556) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1256 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3557) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1255 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3558) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1254 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3559) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1253 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3560) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1252 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3561) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1251 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_121__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n865), .Y(
        oc8051_ram_top1_oc8051_idata_n3562) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1250 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n864) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1249 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3563) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1248 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3564) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1247 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3565) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1246 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3566) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1245 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3567) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1244 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3568) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1243 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3569) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1242 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_120__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n864), .Y(
        oc8051_ram_top1_oc8051_idata_n3570) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1241 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n863) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1240 ( .A(
        oc8051_ram_top1_oc8051_idata_n259), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3571) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1239 ( .A(
        oc8051_ram_top1_oc8051_idata_n258), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3572) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1238 ( .A(
        oc8051_ram_top1_oc8051_idata_n257), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3573) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1237 ( .A(
        oc8051_ram_top1_oc8051_idata_n256), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3574) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1236 ( .A(
        oc8051_ram_top1_oc8051_idata_n255), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3575) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1235 ( .A(
        oc8051_ram_top1_oc8051_idata_n254), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3576) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1234 ( .A(
        oc8051_ram_top1_oc8051_idata_n253), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3577) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1233 ( .A(
        oc8051_ram_top1_oc8051_idata_n252), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n863), .Y(
        oc8051_ram_top1_oc8051_idata_n3578) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1232 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n862) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1231 ( .A(
        oc8051_ram_top1_oc8051_idata_n251), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3579) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1230 ( .A(
        oc8051_ram_top1_oc8051_idata_n250), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3580) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1229 ( .A(
        oc8051_ram_top1_oc8051_idata_n249), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3581) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1228 ( .A(
        oc8051_ram_top1_oc8051_idata_n248), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3582) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1227 ( .A(
        oc8051_ram_top1_oc8051_idata_n247), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3583) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1226 ( .A(
        oc8051_ram_top1_oc8051_idata_n246), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3584) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1225 ( .A(
        oc8051_ram_top1_oc8051_idata_n245), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3585) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1224 ( .A(
        oc8051_ram_top1_oc8051_idata_n244), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n862), .Y(
        oc8051_ram_top1_oc8051_idata_n3586) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1223 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n854) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1222 ( .A(
        oc8051_ram_top1_oc8051_idata_n861), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3587) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1221 ( .A(
        oc8051_ram_top1_oc8051_idata_n860), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3588) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1220 ( .A(
        oc8051_ram_top1_oc8051_idata_n859), .B(
        oc8051_ram_top1_oc8051_idata_n562), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3589) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1219 ( .A(
        oc8051_ram_top1_oc8051_idata_n858), .B(
        oc8051_ram_top1_oc8051_idata_n579), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3590) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1218 ( .A(
        oc8051_ram_top1_oc8051_idata_n857), .B(
        oc8051_ram_top1_oc8051_idata_n596), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3591) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1217 ( .A(
        oc8051_ram_top1_oc8051_idata_n856), .B(
        oc8051_ram_top1_oc8051_idata_n613), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3592) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1216 ( .A(
        oc8051_ram_top1_oc8051_idata_n855), .B(
        oc8051_ram_top1_oc8051_idata_n630), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3593) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1215 ( .A(
        oc8051_ram_top1_oc8051_idata_n853), .B(
        oc8051_ram_top1_oc8051_idata_n647), .S0(
        oc8051_ram_top1_oc8051_idata_n854), .Y(
        oc8051_ram_top1_oc8051_idata_n3594) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1214 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n845) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1213 ( .A(
        oc8051_ram_top1_oc8051_idata_n852), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3595) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1212 ( .A(
        oc8051_ram_top1_oc8051_idata_n851), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3596) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1211 ( .A(
        oc8051_ram_top1_oc8051_idata_n850), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3597) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1210 ( .A(
        oc8051_ram_top1_oc8051_idata_n849), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3598) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1209 ( .A(
        oc8051_ram_top1_oc8051_idata_n848), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3599) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1208 ( .A(
        oc8051_ram_top1_oc8051_idata_n847), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3600) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1207 ( .A(
        oc8051_ram_top1_oc8051_idata_n846), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3601) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1206 ( .A(
        oc8051_ram_top1_oc8051_idata_n844), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n845), .Y(
        oc8051_ram_top1_oc8051_idata_n3602) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1205 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n843) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1204 ( .A(
        oc8051_ram_top1_oc8051_idata_n243), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3603) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1203 ( .A(
        oc8051_ram_top1_oc8051_idata_n242), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3604) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1202 ( .A(
        oc8051_ram_top1_oc8051_idata_n241), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3605) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1201 ( .A(
        oc8051_ram_top1_oc8051_idata_n240), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3606) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1200 ( .A(
        oc8051_ram_top1_oc8051_idata_n239), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3607) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1199 ( .A(
        oc8051_ram_top1_oc8051_idata_n238), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3608) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1198 ( .A(
        oc8051_ram_top1_oc8051_idata_n237), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3609) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1197 ( .A(
        oc8051_ram_top1_oc8051_idata_n236), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n843), .Y(
        oc8051_ram_top1_oc8051_idata_n3610) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1196 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n842) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1195 ( .A(
        oc8051_ram_top1_oc8051_idata_n235), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3611) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1194 ( .A(
        oc8051_ram_top1_oc8051_idata_n234), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3612) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1193 ( .A(
        oc8051_ram_top1_oc8051_idata_n233), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3613) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1192 ( .A(
        oc8051_ram_top1_oc8051_idata_n232), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3614) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1191 ( .A(
        oc8051_ram_top1_oc8051_idata_n231), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3615) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1190 ( .A(
        oc8051_ram_top1_oc8051_idata_n230), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3616) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1189 ( .A(
        oc8051_ram_top1_oc8051_idata_n229), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3617) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1188 ( .A(
        oc8051_ram_top1_oc8051_idata_n228), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n842), .Y(
        oc8051_ram_top1_oc8051_idata_n3618) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1187 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n834) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1186 ( .A(
        oc8051_ram_top1_oc8051_idata_n841), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3619) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1185 ( .A(
        oc8051_ram_top1_oc8051_idata_n840), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3620) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1184 ( .A(
        oc8051_ram_top1_oc8051_idata_n839), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3621) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1183 ( .A(
        oc8051_ram_top1_oc8051_idata_n838), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3622) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1182 ( .A(
        oc8051_ram_top1_oc8051_idata_n837), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3623) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1181 ( .A(
        oc8051_ram_top1_oc8051_idata_n836), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3624) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1180 ( .A(
        oc8051_ram_top1_oc8051_idata_n835), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3625) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1179 ( .A(
        oc8051_ram_top1_oc8051_idata_n833), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n834), .Y(
        oc8051_ram_top1_oc8051_idata_n3626) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1178 ( .A(
        oc8051_ram_top1_oc8051_idata_n832), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n824) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1177 ( .A(
        oc8051_ram_top1_oc8051_idata_n831), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3627) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1176 ( .A(
        oc8051_ram_top1_oc8051_idata_n830), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3628) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1175 ( .A(
        oc8051_ram_top1_oc8051_idata_n829), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3629) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1174 ( .A(
        oc8051_ram_top1_oc8051_idata_n828), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3630) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1173 ( .A(
        oc8051_ram_top1_oc8051_idata_n827), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3631) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1172 ( .A(
        oc8051_ram_top1_oc8051_idata_n826), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3632) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1171 ( .A(
        oc8051_ram_top1_oc8051_idata_n825), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3633) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1170 ( .A(
        oc8051_ram_top1_oc8051_idata_n823), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n824), .Y(
        oc8051_ram_top1_oc8051_idata_n3634) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1169 ( .A(
        oc8051_ram_top1_oc8051_idata_n788), .B(
        oc8051_ram_top1_oc8051_idata_n719), .Y(
        oc8051_ram_top1_oc8051_idata_n807) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1168 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n822) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1167 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3635) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1166 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3636) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1165 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3637) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1164 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3638) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1163 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3639) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1162 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3640) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1161 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3641) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1160 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_111__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n822), .Y(
        oc8051_ram_top1_oc8051_idata_n3642) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1159 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n821) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1158 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__0_), .B(
        oc8051_ram_top1_oc8051_idata_n519), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3643) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1157 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__1_), .B(
        oc8051_ram_top1_oc8051_idata_n536), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3644) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1156 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__2_), .B(
        oc8051_ram_top1_oc8051_idata_n553), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3645) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1155 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__3_), .B(
        oc8051_ram_top1_oc8051_idata_n570), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3646) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1154 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__4_), .B(
        oc8051_ram_top1_oc8051_idata_n587), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3647) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1153 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__5_), .B(
        oc8051_ram_top1_oc8051_idata_n604), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3648) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1152 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__6_), .B(
        oc8051_ram_top1_oc8051_idata_n621), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3649) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1151 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_110__7_), .B(
        oc8051_ram_top1_oc8051_idata_n638), .S0(
        oc8051_ram_top1_oc8051_idata_n821), .Y(
        oc8051_ram_top1_oc8051_idata_n3650) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1150 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n820) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1149 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3651) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1148 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3652) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1147 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3653) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1146 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3654) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1145 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3655) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1144 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3656) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1143 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3657) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1142 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_109__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n820), .Y(
        oc8051_ram_top1_oc8051_idata_n3658) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1141 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n819) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1140 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3659) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1139 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3660) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1138 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3661) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1137 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3662) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1136 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3663) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1135 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3664) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1134 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3665) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1133 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_108__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n819), .Y(
        oc8051_ram_top1_oc8051_idata_n3666) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1132 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n818) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1131 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3667) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1130 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3668) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1129 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3669) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1128 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3670) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1127 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3671) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1126 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3672) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1125 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3673) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1124 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_107__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n818), .Y(
        oc8051_ram_top1_oc8051_idata_n3674) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1123 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n817) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1122 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3675) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1121 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3676) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1120 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3677) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1119 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3678) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1118 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3679) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1117 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3680) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1116 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3681) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1115 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_106__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n817), .Y(
        oc8051_ram_top1_oc8051_idata_n3682) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1114 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n816) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1113 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3683) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1112 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3684) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1111 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3685) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1110 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3686) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1109 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3687) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1108 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3688) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1107 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3689) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1106 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_105__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n816), .Y(
        oc8051_ram_top1_oc8051_idata_n3690) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1105 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n815) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1104 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3691) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1103 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3692) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1102 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3693) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1101 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3694) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1100 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3695) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1099 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3696) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1098 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3697) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1097 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_104__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n815), .Y(
        oc8051_ram_top1_oc8051_idata_n3698) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1096 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n814) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1095 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3699) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1094 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3700) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1093 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3701) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1092 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3702) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1091 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3703) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1090 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3704) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1089 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3705) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1088 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_103__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n814), .Y(
        oc8051_ram_top1_oc8051_idata_n3706) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1087 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n813) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1086 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3707) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1085 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3708) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1084 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3709) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1083 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3710) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1082 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3711) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1081 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3712) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1080 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3713) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1079 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_102__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n813), .Y(
        oc8051_ram_top1_oc8051_idata_n3714) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1078 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n812) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1077 ( .A(
        oc8051_ram_top1_oc8051_idata_n227), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3715) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1076 ( .A(
        oc8051_ram_top1_oc8051_idata_n226), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3716) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1075 ( .A(
        oc8051_ram_top1_oc8051_idata_n225), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3717) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1074 ( .A(
        oc8051_ram_top1_oc8051_idata_n224), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3718) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1073 ( .A(
        oc8051_ram_top1_oc8051_idata_n223), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3719) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1072 ( .A(
        oc8051_ram_top1_oc8051_idata_n222), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3720) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1071 ( .A(
        oc8051_ram_top1_oc8051_idata_n221), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3721) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1070 ( .A(
        oc8051_ram_top1_oc8051_idata_n220), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n812), .Y(
        oc8051_ram_top1_oc8051_idata_n3722) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1069 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n811) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1068 ( .A(
        oc8051_ram_top1_oc8051_idata_n219), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3723) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1067 ( .A(
        oc8051_ram_top1_oc8051_idata_n218), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3724) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1066 ( .A(
        oc8051_ram_top1_oc8051_idata_n217), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3725) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1065 ( .A(
        oc8051_ram_top1_oc8051_idata_n216), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3726) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1064 ( .A(
        oc8051_ram_top1_oc8051_idata_n215), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3727) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1063 ( .A(
        oc8051_ram_top1_oc8051_idata_n214), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3728) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1062 ( .A(
        oc8051_ram_top1_oc8051_idata_n213), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3729) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1061 ( .A(
        oc8051_ram_top1_oc8051_idata_n212), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n811), .Y(
        oc8051_ram_top1_oc8051_idata_n3730) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1060 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n810) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1059 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3731) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1058 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3732) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1057 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3733) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1056 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3734) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1055 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3735) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1054 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3736) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1053 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3737) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1052 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_99__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n810), .Y(
        oc8051_ram_top1_oc8051_idata_n3738) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1051 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n809) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1050 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3739) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1049 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3740) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1048 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3741) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1047 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3742) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1046 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3743) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1045 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3744) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1044 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3745) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1043 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_98__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n809), .Y(
        oc8051_ram_top1_oc8051_idata_n3746) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1042 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n808) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1041 ( .A(
        oc8051_ram_top1_oc8051_idata_n211), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3747) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1040 ( .A(
        oc8051_ram_top1_oc8051_idata_n210), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3748) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1039 ( .A(
        oc8051_ram_top1_oc8051_idata_n209), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3749) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1038 ( .A(
        oc8051_ram_top1_oc8051_idata_n208), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3750) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1037 ( .A(
        oc8051_ram_top1_oc8051_idata_n207), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3751) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1036 ( .A(
        oc8051_ram_top1_oc8051_idata_n206), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3752) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1035 ( .A(
        oc8051_ram_top1_oc8051_idata_n205), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3753) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1034 ( .A(
        oc8051_ram_top1_oc8051_idata_n204), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n808), .Y(
        oc8051_ram_top1_oc8051_idata_n3754) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1033 ( .A(
        oc8051_ram_top1_oc8051_idata_n807), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n806) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1032 ( .A(
        oc8051_ram_top1_oc8051_idata_n203), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3755) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1031 ( .A(
        oc8051_ram_top1_oc8051_idata_n202), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3756) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1030 ( .A(
        oc8051_ram_top1_oc8051_idata_n201), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3757) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1029 ( .A(
        oc8051_ram_top1_oc8051_idata_n200), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3758) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1028 ( .A(
        oc8051_ram_top1_oc8051_idata_n199), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3759) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1027 ( .A(
        oc8051_ram_top1_oc8051_idata_n198), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3760) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1026 ( .A(
        oc8051_ram_top1_oc8051_idata_n197), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3761) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1025 ( .A(
        oc8051_ram_top1_oc8051_idata_n196), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n806), .Y(
        oc8051_ram_top1_oc8051_idata_n3762) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1024 ( .A(
        oc8051_ram_top1_oc8051_idata_n788), .B(
        oc8051_ram_top1_oc8051_idata_n701), .Y(
        oc8051_ram_top1_oc8051_idata_n790) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1023 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n805) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1022 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3763) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1021 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3764) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1020 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3765) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1019 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3766) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1018 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3767) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1017 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3768) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1016 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3769) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1015 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_95__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n805), .Y(
        oc8051_ram_top1_oc8051_idata_n3770) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1014 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n804) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1013 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3771) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1012 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3772) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1011 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3773) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1010 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3774) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1009 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3775) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1008 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3776) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1007 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3777) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1006 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_94__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n804), .Y(
        oc8051_ram_top1_oc8051_idata_n3778) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1005 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n803) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1004 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__0_), .B(
        oc8051_ram_top1_oc8051_idata_n518), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3779) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1003 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__1_), .B(
        oc8051_ram_top1_oc8051_idata_n535), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3780) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1002 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__2_), .B(
        oc8051_ram_top1_oc8051_idata_n552), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3781) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1001 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__3_), .B(
        oc8051_ram_top1_oc8051_idata_n569), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3782) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u1000 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__4_), .B(
        oc8051_ram_top1_oc8051_idata_n586), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3783) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u999 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__5_), .B(
        oc8051_ram_top1_oc8051_idata_n603), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3784) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u998 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__6_), .B(
        oc8051_ram_top1_oc8051_idata_n620), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3785) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u997 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_93__7_), .B(
        oc8051_ram_top1_oc8051_idata_n637), .S0(
        oc8051_ram_top1_oc8051_idata_n803), .Y(
        oc8051_ram_top1_oc8051_idata_n3786) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u996 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n802) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u995 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3787) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u994 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3788) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u993 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3789) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u992 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3790) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u991 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3791) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u990 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3792) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u989 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3793) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u988 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_92__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n802), .Y(
        oc8051_ram_top1_oc8051_idata_n3794) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u987 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n801) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u986 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3795) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u985 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3796) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u984 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3797) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u983 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3798) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u982 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3799) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u981 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3800) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u980 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3801) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u979 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_91__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n801), .Y(
        oc8051_ram_top1_oc8051_idata_n3802) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u978 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n800) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u977 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3803) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u976 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3804) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u975 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3805) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u974 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3806) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u973 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3807) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u972 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3808) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u971 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3809) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u970 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_90__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n800), .Y(
        oc8051_ram_top1_oc8051_idata_n3810) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u969 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n799) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u968 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3811) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u967 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3812) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u966 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3813) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u965 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3814) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u964 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3815) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u963 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3816) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u962 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3817) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u961 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_89__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n799), .Y(
        oc8051_ram_top1_oc8051_idata_n3818) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u960 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n798) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u959 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3819) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u958 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3820) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u957 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3821) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u956 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3822) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u955 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3823) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u954 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3824) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u953 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3825) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u952 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_88__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n798), .Y(
        oc8051_ram_top1_oc8051_idata_n3826) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u951 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n797) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u950 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3827) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u949 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3828) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u948 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3829) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u947 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3830) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u946 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3831) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u945 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3832) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u944 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3833) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u943 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_87__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n797), .Y(
        oc8051_ram_top1_oc8051_idata_n3834) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u942 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n796) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u941 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3835) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u940 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3836) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u939 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3837) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u938 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3838) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u937 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3839) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u936 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3840) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u935 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3841) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u934 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_86__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n796), .Y(
        oc8051_ram_top1_oc8051_idata_n3842) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u933 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n795) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u932 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3843) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u931 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3844) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u930 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3845) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u929 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3846) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u928 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3847) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u927 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3848) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u926 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3849) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u925 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_85__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n795), .Y(
        oc8051_ram_top1_oc8051_idata_n3850) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u924 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n794) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u923 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3851) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u922 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3852) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u921 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3853) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u920 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3854) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u919 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3855) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u918 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3856) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u917 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3857) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u916 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_84__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n794), .Y(
        oc8051_ram_top1_oc8051_idata_n3858) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u915 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n793) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u914 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3859) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u913 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3860) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u912 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3861) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u911 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3862) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u910 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3863) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u909 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3864) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u908 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3865) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u907 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_83__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n793), .Y(
        oc8051_ram_top1_oc8051_idata_n3866) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u906 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n792) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u905 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3867) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u904 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3868) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u903 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3869) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u902 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3870) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u901 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3871) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u900 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3872) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u899 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3873) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u898 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_82__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n792), .Y(
        oc8051_ram_top1_oc8051_idata_n3874) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u897 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n791) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u896 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3875) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u895 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3876) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u894 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3877) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u893 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3878) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u892 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3879) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u891 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3880) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u890 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3881) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u889 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_81__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n791), .Y(
        oc8051_ram_top1_oc8051_idata_n3882) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u888 ( .A(
        oc8051_ram_top1_oc8051_idata_n790), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n789) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u887 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__0_), .B(
        oc8051_ram_top1_oc8051_idata_n517), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3883) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u886 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__1_), .B(
        oc8051_ram_top1_oc8051_idata_n534), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3884) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u885 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__2_), .B(
        oc8051_ram_top1_oc8051_idata_n551), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3885) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u884 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__3_), .B(
        oc8051_ram_top1_oc8051_idata_n568), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3886) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u883 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__4_), .B(
        oc8051_ram_top1_oc8051_idata_n585), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3887) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u882 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__5_), .B(
        oc8051_ram_top1_oc8051_idata_n602), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3888) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u881 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__6_), .B(
        oc8051_ram_top1_oc8051_idata_n619), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3889) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u880 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_80__7_), .B(
        oc8051_ram_top1_oc8051_idata_n636), .S0(
        oc8051_ram_top1_oc8051_idata_n789), .Y(
        oc8051_ram_top1_oc8051_idata_n3890) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u879 ( .A(
        oc8051_ram_top1_oc8051_idata_n788), .B(
        oc8051_ram_top1_oc8051_idata_n683), .Y(
        oc8051_ram_top1_oc8051_idata_n772) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u878 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n787) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u877 ( .A(
        oc8051_ram_top1_oc8051_idata_n195), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3891) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u876 ( .A(
        oc8051_ram_top1_oc8051_idata_n194), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3892) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u875 ( .A(
        oc8051_ram_top1_oc8051_idata_n193), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3893) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u874 ( .A(
        oc8051_ram_top1_oc8051_idata_n192), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3894) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u873 ( .A(
        oc8051_ram_top1_oc8051_idata_n191), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3895) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u872 ( .A(
        oc8051_ram_top1_oc8051_idata_n190), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3896) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u871 ( .A(
        oc8051_ram_top1_oc8051_idata_n189), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3897) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u870 ( .A(
        oc8051_ram_top1_oc8051_idata_n188), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n787), .Y(
        oc8051_ram_top1_oc8051_idata_n3898) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u869 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n786) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u868 ( .A(
        oc8051_ram_top1_oc8051_idata_n187), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3899) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u867 ( .A(
        oc8051_ram_top1_oc8051_idata_n186), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3900) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u866 ( .A(
        oc8051_ram_top1_oc8051_idata_n185), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3901) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u865 ( .A(
        oc8051_ram_top1_oc8051_idata_n184), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3902) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u864 ( .A(
        oc8051_ram_top1_oc8051_idata_n183), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3903) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u863 ( .A(
        oc8051_ram_top1_oc8051_idata_n182), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3904) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u862 ( .A(
        oc8051_ram_top1_oc8051_idata_n181), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3905) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u861 ( .A(
        oc8051_ram_top1_oc8051_idata_n180), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n786), .Y(
        oc8051_ram_top1_oc8051_idata_n3906) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u860 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n785) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u859 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3907) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u858 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3908) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u857 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3909) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u856 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3910) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u855 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3911) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u854 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3912) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u853 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3913) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u852 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_77__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n785), .Y(
        oc8051_ram_top1_oc8051_idata_n3914) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u851 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n784) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u850 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3915) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u849 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3916) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u848 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3917) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u847 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3918) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u846 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3919) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u845 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3920) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u844 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3921) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u843 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_76__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n784), .Y(
        oc8051_ram_top1_oc8051_idata_n3922) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u842 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n783) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u841 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3923) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u840 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3924) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u839 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3925) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u838 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3926) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u837 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3927) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u836 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3928) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u835 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3929) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u834 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_75__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n783), .Y(
        oc8051_ram_top1_oc8051_idata_n3930) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u833 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n782) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u832 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3931) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u831 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3932) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u830 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3933) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u829 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3934) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u828 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3935) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u827 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3936) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u826 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3937) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u825 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_74__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n782), .Y(
        oc8051_ram_top1_oc8051_idata_n3938) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u824 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n781) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u823 ( .A(
        oc8051_ram_top1_oc8051_idata_n179), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3939) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u822 ( .A(
        oc8051_ram_top1_oc8051_idata_n178), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3940) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u821 ( .A(
        oc8051_ram_top1_oc8051_idata_n177), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3941) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u820 ( .A(
        oc8051_ram_top1_oc8051_idata_n176), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3942) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u819 ( .A(
        oc8051_ram_top1_oc8051_idata_n175), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3943) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u818 ( .A(
        oc8051_ram_top1_oc8051_idata_n174), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3944) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u817 ( .A(
        oc8051_ram_top1_oc8051_idata_n173), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3945) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u816 ( .A(
        oc8051_ram_top1_oc8051_idata_n172), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n781), .Y(
        oc8051_ram_top1_oc8051_idata_n3946) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u815 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n780) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u814 ( .A(
        oc8051_ram_top1_oc8051_idata_n171), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3947) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u813 ( .A(
        oc8051_ram_top1_oc8051_idata_n170), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3948) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u812 ( .A(
        oc8051_ram_top1_oc8051_idata_n169), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3949) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u811 ( .A(
        oc8051_ram_top1_oc8051_idata_n168), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3950) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u810 ( .A(
        oc8051_ram_top1_oc8051_idata_n167), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3951) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u809 ( .A(
        oc8051_ram_top1_oc8051_idata_n166), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3952) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u808 ( .A(
        oc8051_ram_top1_oc8051_idata_n165), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3953) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u807 ( .A(
        oc8051_ram_top1_oc8051_idata_n164), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n780), .Y(
        oc8051_ram_top1_oc8051_idata_n3954) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u806 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n779) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u805 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3955) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u804 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3956) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u803 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3957) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u802 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3958) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u801 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3959) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u800 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3960) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u799 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3961) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u798 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_71__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n779), .Y(
        oc8051_ram_top1_oc8051_idata_n3962) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u797 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n778) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u796 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3963) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u795 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3964) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u794 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3965) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u793 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3966) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u792 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3967) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u791 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3968) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u790 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3969) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u789 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_70__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n778), .Y(
        oc8051_ram_top1_oc8051_idata_n3970) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u788 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n777) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u787 ( .A(
        oc8051_ram_top1_oc8051_idata_n163), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3971) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u786 ( .A(
        oc8051_ram_top1_oc8051_idata_n162), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3972) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u785 ( .A(
        oc8051_ram_top1_oc8051_idata_n161), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3973) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u784 ( .A(
        oc8051_ram_top1_oc8051_idata_n160), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3974) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u783 ( .A(
        oc8051_ram_top1_oc8051_idata_n159), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3975) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u782 ( .A(
        oc8051_ram_top1_oc8051_idata_n158), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3976) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u781 ( .A(
        oc8051_ram_top1_oc8051_idata_n157), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3977) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u780 ( .A(
        oc8051_ram_top1_oc8051_idata_n156), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n777), .Y(
        oc8051_ram_top1_oc8051_idata_n3978) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u779 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n776) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u778 ( .A(
        oc8051_ram_top1_oc8051_idata_n155), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3979) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u777 ( .A(
        oc8051_ram_top1_oc8051_idata_n154), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3980) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u776 ( .A(
        oc8051_ram_top1_oc8051_idata_n153), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3981) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u775 ( .A(
        oc8051_ram_top1_oc8051_idata_n152), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3982) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u774 ( .A(
        oc8051_ram_top1_oc8051_idata_n151), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3983) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u773 ( .A(
        oc8051_ram_top1_oc8051_idata_n150), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3984) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u772 ( .A(
        oc8051_ram_top1_oc8051_idata_n149), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3985) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u771 ( .A(
        oc8051_ram_top1_oc8051_idata_n148), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n776), .Y(
        oc8051_ram_top1_oc8051_idata_n3986) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u770 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n775) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u769 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3987) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u768 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3988) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u767 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3989) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u766 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3990) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u765 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3991) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u764 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3992) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u763 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3993) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u762 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_67__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n775), .Y(
        oc8051_ram_top1_oc8051_idata_n3994) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u761 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n774) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u760 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n3995) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u759 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n3996) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u758 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n3997) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u757 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n3998) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u756 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n3999) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u755 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n4000) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u754 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n4001) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u753 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_66__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n774), .Y(
        oc8051_ram_top1_oc8051_idata_n4002) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u752 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n773) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u751 ( .A(
        oc8051_ram_top1_oc8051_idata_n147), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4003) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u750 ( .A(
        oc8051_ram_top1_oc8051_idata_n146), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4004) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u749 ( .A(
        oc8051_ram_top1_oc8051_idata_n145), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4005) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u748 ( .A(
        oc8051_ram_top1_oc8051_idata_n144), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4006) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u747 ( .A(
        oc8051_ram_top1_oc8051_idata_n143), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4007) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u746 ( .A(
        oc8051_ram_top1_oc8051_idata_n142), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4008) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u745 ( .A(
        oc8051_ram_top1_oc8051_idata_n141), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4009) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u744 ( .A(
        oc8051_ram_top1_oc8051_idata_n140), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n773), .Y(
        oc8051_ram_top1_oc8051_idata_n4010) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u743 ( .A(
        oc8051_ram_top1_oc8051_idata_n772), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n771) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u742 ( .A(
        oc8051_ram_top1_oc8051_idata_n139), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4011) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u741 ( .A(
        oc8051_ram_top1_oc8051_idata_n138), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4012) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u740 ( .A(
        oc8051_ram_top1_oc8051_idata_n137), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4013) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u739 ( .A(
        oc8051_ram_top1_oc8051_idata_n136), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4014) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u738 ( .A(
        oc8051_ram_top1_oc8051_idata_n135), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4015) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u737 ( .A(
        oc8051_ram_top1_oc8051_idata_n134), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4016) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u736 ( .A(
        oc8051_ram_top1_oc8051_idata_n133), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4017) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u735 ( .A(
        oc8051_ram_top1_oc8051_idata_n132), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n771), .Y(
        oc8051_ram_top1_oc8051_idata_n4018) );
  NOR2B_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u734 ( .AN(
        oc8051_ram_top1_oc8051_idata_n770), .B(oc8051_ram_top1_wr_addr_m_6_), 
        .Y(oc8051_ram_top1_oc8051_idata_n682) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u733 ( .A(
        oc8051_ram_top1_oc8051_idata_n769), .B(
        oc8051_ram_top1_oc8051_idata_n682), .Y(
        oc8051_ram_top1_oc8051_idata_n729) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u732 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n768) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u731 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4019) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u730 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4020) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u729 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4021) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u728 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4022) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u727 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4023) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u726 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4024) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u725 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4025) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u724 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_63__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n768), .Y(
        oc8051_ram_top1_oc8051_idata_n4026) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u723 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n767) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u722 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4027) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u721 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4028) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u720 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4029) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u719 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4030) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u718 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4031) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u717 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4032) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u716 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4033) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u715 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_62__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n767), .Y(
        oc8051_ram_top1_oc8051_idata_n4034) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u714 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n766) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u713 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4035) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u712 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4036) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u711 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4037) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u710 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4038) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u709 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4039) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u708 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4040) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u707 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4041) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u706 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_61__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n766), .Y(
        oc8051_ram_top1_oc8051_idata_n4042) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u705 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n765) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u704 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4043) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u703 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4044) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u702 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4045) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u701 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4046) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u700 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4047) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u699 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4048) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u698 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4049) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u697 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_60__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n765), .Y(
        oc8051_ram_top1_oc8051_idata_n4050) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u696 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n764) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u695 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__0_), .B(
        oc8051_ram_top1_oc8051_idata_n516), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4051) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u694 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__1_), .B(
        oc8051_ram_top1_oc8051_idata_n533), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4052) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u693 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__2_), .B(
        oc8051_ram_top1_oc8051_idata_n550), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4053) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u692 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__3_), .B(
        oc8051_ram_top1_oc8051_idata_n567), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4054) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u691 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__4_), .B(
        oc8051_ram_top1_oc8051_idata_n584), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4055) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u690 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__5_), .B(
        oc8051_ram_top1_oc8051_idata_n601), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4056) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u689 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__6_), .B(
        oc8051_ram_top1_oc8051_idata_n618), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4057) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u688 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_59__7_), .B(
        oc8051_ram_top1_oc8051_idata_n635), .S0(
        oc8051_ram_top1_oc8051_idata_n764), .Y(
        oc8051_ram_top1_oc8051_idata_n4058) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u687 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n763) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u686 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4059) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u685 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4060) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u684 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4061) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u683 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4062) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u682 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4063) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u681 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4064) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u680 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4065) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u679 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_58__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n763), .Y(
        oc8051_ram_top1_oc8051_idata_n4066) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u678 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n762) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u677 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4067) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u676 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4068) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u675 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4069) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u674 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4070) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u673 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4071) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u672 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4072) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u671 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4073) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u670 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_57__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n762), .Y(
        oc8051_ram_top1_oc8051_idata_n4074) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u669 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n761) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u668 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4075) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u667 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4076) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u666 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4077) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u665 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4078) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u664 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4079) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u663 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4080) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u662 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4081) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u661 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_56__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n761), .Y(
        oc8051_ram_top1_oc8051_idata_n4082) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u660 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n760) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u659 ( .A(
        oc8051_ram_top1_oc8051_idata_n131), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4083) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u658 ( .A(
        oc8051_ram_top1_oc8051_idata_n130), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4084) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u657 ( .A(
        oc8051_ram_top1_oc8051_idata_n129), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4085) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u656 ( .A(
        oc8051_ram_top1_oc8051_idata_n128), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4086) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u655 ( .A(
        oc8051_ram_top1_oc8051_idata_n127), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4087) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u654 ( .A(
        oc8051_ram_top1_oc8051_idata_n126), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4088) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u653 ( .A(
        oc8051_ram_top1_oc8051_idata_n125), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4089) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u652 ( .A(
        oc8051_ram_top1_oc8051_idata_n124), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n760), .Y(
        oc8051_ram_top1_oc8051_idata_n4090) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u651 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n759) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u650 ( .A(
        oc8051_ram_top1_oc8051_idata_n123), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4091) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u649 ( .A(
        oc8051_ram_top1_oc8051_idata_n122), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4092) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u648 ( .A(
        oc8051_ram_top1_oc8051_idata_n121), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4093) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u647 ( .A(
        oc8051_ram_top1_oc8051_idata_n120), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4094) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u646 ( .A(
        oc8051_ram_top1_oc8051_idata_n119), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4095) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u645 ( .A(
        oc8051_ram_top1_oc8051_idata_n118), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4096) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u644 ( .A(
        oc8051_ram_top1_oc8051_idata_n117), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4097) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u643 ( .A(
        oc8051_ram_top1_oc8051_idata_n116), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n759), .Y(
        oc8051_ram_top1_oc8051_idata_n4098) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u642 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n751) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u641 ( .A(
        oc8051_ram_top1_oc8051_idata_n758), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4099) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u640 ( .A(
        oc8051_ram_top1_oc8051_idata_n757), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4100) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u639 ( .A(
        oc8051_ram_top1_oc8051_idata_n756), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4101) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u638 ( .A(
        oc8051_ram_top1_oc8051_idata_n755), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4102) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u637 ( .A(
        oc8051_ram_top1_oc8051_idata_n754), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4103) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u636 ( .A(
        oc8051_ram_top1_oc8051_idata_n753), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4104) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u635 ( .A(
        oc8051_ram_top1_oc8051_idata_n752), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4105) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u634 ( .A(
        oc8051_ram_top1_oc8051_idata_n750), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n751), .Y(
        oc8051_ram_top1_oc8051_idata_n4106) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u633 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n742) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u632 ( .A(
        oc8051_ram_top1_oc8051_idata_n749), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4107) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u631 ( .A(
        oc8051_ram_top1_oc8051_idata_n748), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4108) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u630 ( .A(
        oc8051_ram_top1_oc8051_idata_n747), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4109) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u629 ( .A(
        oc8051_ram_top1_oc8051_idata_n746), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4110) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u628 ( .A(
        oc8051_ram_top1_oc8051_idata_n745), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4111) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u627 ( .A(
        oc8051_ram_top1_oc8051_idata_n744), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4112) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u626 ( .A(
        oc8051_ram_top1_oc8051_idata_n743), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4113) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u625 ( .A(
        oc8051_ram_top1_oc8051_idata_n741), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n742), .Y(
        oc8051_ram_top1_oc8051_idata_n4114) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u624 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n740) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u623 ( .A(
        oc8051_ram_top1_oc8051_idata_n115), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4115) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u622 ( .A(
        oc8051_ram_top1_oc8051_idata_n114), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4116) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u621 ( .A(
        oc8051_ram_top1_oc8051_idata_n113), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4117) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u620 ( .A(
        oc8051_ram_top1_oc8051_idata_n112), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4118) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u619 ( .A(
        oc8051_ram_top1_oc8051_idata_n111), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4119) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u618 ( .A(
        oc8051_ram_top1_oc8051_idata_n110), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4120) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u617 ( .A(
        oc8051_ram_top1_oc8051_idata_n109), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4121) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u616 ( .A(
        oc8051_ram_top1_oc8051_idata_n108), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n740), .Y(
        oc8051_ram_top1_oc8051_idata_n4122) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u615 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n739) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u614 ( .A(
        oc8051_ram_top1_oc8051_idata_n107), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4123) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u613 ( .A(
        oc8051_ram_top1_oc8051_idata_n106), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4124) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u612 ( .A(
        oc8051_ram_top1_oc8051_idata_n105), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4125) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u611 ( .A(
        oc8051_ram_top1_oc8051_idata_n104), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4126) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u610 ( .A(
        oc8051_ram_top1_oc8051_idata_n103), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4127) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u609 ( .A(
        oc8051_ram_top1_oc8051_idata_n102), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4128) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u608 ( .A(
        oc8051_ram_top1_oc8051_idata_n101), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4129) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u607 ( .A(
        oc8051_ram_top1_oc8051_idata_n100), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n739), .Y(
        oc8051_ram_top1_oc8051_idata_n4130) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u606 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n731) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u605 ( .A(
        oc8051_ram_top1_oc8051_idata_n738), .B(
        oc8051_ram_top1_oc8051_idata_n527), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4131) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u604 ( .A(
        oc8051_ram_top1_oc8051_idata_n737), .B(
        oc8051_ram_top1_oc8051_idata_n544), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4132) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u603 ( .A(
        oc8051_ram_top1_oc8051_idata_n736), .B(
        oc8051_ram_top1_oc8051_idata_n561), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4133) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u602 ( .A(
        oc8051_ram_top1_oc8051_idata_n735), .B(
        oc8051_ram_top1_oc8051_idata_n578), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4134) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u601 ( .A(
        oc8051_ram_top1_oc8051_idata_n734), .B(
        oc8051_ram_top1_oc8051_idata_n595), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4135) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u600 ( .A(
        oc8051_ram_top1_oc8051_idata_n733), .B(
        oc8051_ram_top1_oc8051_idata_n612), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4136) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u599 ( .A(
        oc8051_ram_top1_oc8051_idata_n732), .B(
        oc8051_ram_top1_oc8051_idata_n629), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4137) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u598 ( .A(
        oc8051_ram_top1_oc8051_idata_n730), .B(
        oc8051_ram_top1_oc8051_idata_n646), .S0(
        oc8051_ram_top1_oc8051_idata_n731), .Y(
        oc8051_ram_top1_oc8051_idata_n4138) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u597 ( .A(
        oc8051_ram_top1_oc8051_idata_n729), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n721) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u596 ( .A(
        oc8051_ram_top1_oc8051_idata_n728), .B(
        oc8051_ram_top1_oc8051_idata_n526), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4139) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u595 ( .A(
        oc8051_ram_top1_oc8051_idata_n727), .B(
        oc8051_ram_top1_oc8051_idata_n543), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4140) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u594 ( .A(
        oc8051_ram_top1_oc8051_idata_n726), .B(
        oc8051_ram_top1_oc8051_idata_n560), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4141) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u593 ( .A(
        oc8051_ram_top1_oc8051_idata_n725), .B(
        oc8051_ram_top1_oc8051_idata_n577), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4142) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u592 ( .A(
        oc8051_ram_top1_oc8051_idata_n724), .B(
        oc8051_ram_top1_oc8051_idata_n594), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4143) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u591 ( .A(
        oc8051_ram_top1_oc8051_idata_n723), .B(
        oc8051_ram_top1_oc8051_idata_n611), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4144) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u590 ( .A(
        oc8051_ram_top1_oc8051_idata_n722), .B(
        oc8051_ram_top1_oc8051_idata_n628), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4145) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u589 ( .A(
        oc8051_ram_top1_oc8051_idata_n720), .B(
        oc8051_ram_top1_oc8051_idata_n645), .S0(
        oc8051_ram_top1_oc8051_idata_n721), .Y(
        oc8051_ram_top1_oc8051_idata_n4146) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u588 ( .A(
        oc8051_ram_top1_oc8051_idata_n719), .B(
        oc8051_ram_top1_oc8051_idata_n682), .Y(
        oc8051_ram_top1_oc8051_idata_n703) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u587 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n718) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u586 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4147) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u585 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4148) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u584 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4149) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u583 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4150) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u582 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4151) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u581 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4152) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u580 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4153) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u579 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_47__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n718), .Y(
        oc8051_ram_top1_oc8051_idata_n4154) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u578 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n717) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u577 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4155) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u576 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4156) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u575 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4157) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u574 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4158) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u573 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4159) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u572 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4160) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u571 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4161) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u570 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_46__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n717), .Y(
        oc8051_ram_top1_oc8051_idata_n4162) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u569 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n716) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u568 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4163) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u567 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4164) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u566 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4165) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u565 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4166) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u564 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4167) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u563 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4168) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u562 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4169) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u561 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_45__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n716), .Y(
        oc8051_ram_top1_oc8051_idata_n4170) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u560 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n715) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u559 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4171) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u558 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4172) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u557 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4173) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u556 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4174) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u555 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4175) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u554 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4176) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u553 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4177) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u552 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_44__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n715), .Y(
        oc8051_ram_top1_oc8051_idata_n4178) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u551 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n714) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u550 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4179) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u549 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4180) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u548 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4181) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u547 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4182) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u546 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4183) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u545 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4184) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u544 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4185) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u543 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_43__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n714), .Y(
        oc8051_ram_top1_oc8051_idata_n4186) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u542 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n713) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u541 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4187) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u540 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4188) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u539 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4189) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u538 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4190) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u537 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4191) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u536 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4192) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u535 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4193) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u534 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_42__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n713), .Y(
        oc8051_ram_top1_oc8051_idata_n4194) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u533 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n712) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u532 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4195) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u531 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4196) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u530 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4197) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u529 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4198) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u528 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4199) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u527 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4200) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u526 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4201) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u525 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_41__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n712), .Y(
        oc8051_ram_top1_oc8051_idata_n4202) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u524 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n711) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u523 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4203) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u522 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4204) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u521 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4205) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u520 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4206) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u519 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4207) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u518 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4208) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u517 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4209) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u516 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_40__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n711), .Y(
        oc8051_ram_top1_oc8051_idata_n4210) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u515 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n710) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u514 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4211) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u513 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4212) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u512 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4213) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u511 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4214) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u510 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4215) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u509 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4216) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u508 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4217) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u507 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_39__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n710), .Y(
        oc8051_ram_top1_oc8051_idata_n4218) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u506 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n709) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u505 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__0_), .B(
        oc8051_ram_top1_oc8051_idata_n3), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4219) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u504 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__1_), .B(
        oc8051_ram_top1_oc8051_idata_n532), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4220) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u503 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__2_), .B(
        oc8051_ram_top1_oc8051_idata_n549), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4221) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u502 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__3_), .B(
        oc8051_ram_top1_oc8051_idata_n566), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4222) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u501 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__4_), .B(
        oc8051_ram_top1_oc8051_idata_n583), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4223) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u500 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__5_), .B(
        oc8051_ram_top1_oc8051_idata_n600), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4224) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u499 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__6_), .B(
        oc8051_ram_top1_oc8051_idata_n617), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4225) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u498 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_38__7_), .B(
        oc8051_ram_top1_oc8051_idata_n634), .S0(
        oc8051_ram_top1_oc8051_idata_n709), .Y(
        oc8051_ram_top1_oc8051_idata_n4226) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u497 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n708) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u496 ( .A(
        oc8051_ram_top1_oc8051_idata_n99), .B(
        oc8051_ram_top1_oc8051_idata_n526), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4227) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u495 ( .A(
        oc8051_ram_top1_oc8051_idata_n98), .B(
        oc8051_ram_top1_oc8051_idata_n543), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4228) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u494 ( .A(
        oc8051_ram_top1_oc8051_idata_n97), .B(
        oc8051_ram_top1_oc8051_idata_n560), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4229) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u493 ( .A(
        oc8051_ram_top1_oc8051_idata_n96), .B(
        oc8051_ram_top1_oc8051_idata_n577), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4230) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u492 ( .A(
        oc8051_ram_top1_oc8051_idata_n95), .B(
        oc8051_ram_top1_oc8051_idata_n594), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4231) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u491 ( .A(
        oc8051_ram_top1_oc8051_idata_n94), .B(
        oc8051_ram_top1_oc8051_idata_n611), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4232) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u490 ( .A(
        oc8051_ram_top1_oc8051_idata_n93), .B(
        oc8051_ram_top1_oc8051_idata_n628), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4233) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u489 ( .A(
        oc8051_ram_top1_oc8051_idata_n92), .B(
        oc8051_ram_top1_oc8051_idata_n645), .S0(
        oc8051_ram_top1_oc8051_idata_n708), .Y(
        oc8051_ram_top1_oc8051_idata_n4234) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u488 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n707) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u487 ( .A(
        oc8051_ram_top1_oc8051_idata_n91), .B(
        oc8051_ram_top1_oc8051_idata_n526), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4235) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u486 ( .A(
        oc8051_ram_top1_oc8051_idata_n90), .B(
        oc8051_ram_top1_oc8051_idata_n543), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4236) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u485 ( .A(
        oc8051_ram_top1_oc8051_idata_n89), .B(
        oc8051_ram_top1_oc8051_idata_n560), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4237) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u484 ( .A(
        oc8051_ram_top1_oc8051_idata_n88), .B(
        oc8051_ram_top1_oc8051_idata_n577), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4238) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u483 ( .A(
        oc8051_ram_top1_oc8051_idata_n87), .B(
        oc8051_ram_top1_oc8051_idata_n594), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4239) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u482 ( .A(
        oc8051_ram_top1_oc8051_idata_n86), .B(
        oc8051_ram_top1_oc8051_idata_n611), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4240) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u481 ( .A(
        oc8051_ram_top1_oc8051_idata_n85), .B(
        oc8051_ram_top1_oc8051_idata_n628), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4241) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u480 ( .A(
        oc8051_ram_top1_oc8051_idata_n84), .B(
        oc8051_ram_top1_oc8051_idata_n645), .S0(
        oc8051_ram_top1_oc8051_idata_n707), .Y(
        oc8051_ram_top1_oc8051_idata_n4242) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u479 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n706) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u478 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4243) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u477 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4244) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u476 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4245) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u475 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4246) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u474 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4247) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u473 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4248) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u472 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4249) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u471 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_35__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n706), .Y(
        oc8051_ram_top1_oc8051_idata_n4250) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u470 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n705) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u469 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4251) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u468 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4252) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u467 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4253) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u466 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4254) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u465 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4255) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u464 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4256) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u463 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4257) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u462 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_34__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n705), .Y(
        oc8051_ram_top1_oc8051_idata_n4258) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u461 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n704) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u460 ( .A(
        oc8051_ram_top1_oc8051_idata_n83), .B(
        oc8051_ram_top1_oc8051_idata_n525), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4259) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u459 ( .A(
        oc8051_ram_top1_oc8051_idata_n82), .B(
        oc8051_ram_top1_oc8051_idata_n542), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4260) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u458 ( .A(
        oc8051_ram_top1_oc8051_idata_n81), .B(
        oc8051_ram_top1_oc8051_idata_n559), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4261) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u457 ( .A(
        oc8051_ram_top1_oc8051_idata_n80), .B(
        oc8051_ram_top1_oc8051_idata_n576), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4262) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u456 ( .A(
        oc8051_ram_top1_oc8051_idata_n79), .B(
        oc8051_ram_top1_oc8051_idata_n593), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4263) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u455 ( .A(
        oc8051_ram_top1_oc8051_idata_n78), .B(
        oc8051_ram_top1_oc8051_idata_n610), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4264) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u454 ( .A(
        oc8051_ram_top1_oc8051_idata_n77), .B(
        oc8051_ram_top1_oc8051_idata_n627), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4265) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u453 ( .A(
        oc8051_ram_top1_oc8051_idata_n76), .B(
        oc8051_ram_top1_oc8051_idata_n644), .S0(
        oc8051_ram_top1_oc8051_idata_n704), .Y(
        oc8051_ram_top1_oc8051_idata_n4266) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u452 ( .A(
        oc8051_ram_top1_oc8051_idata_n703), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n702) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u451 ( .A(
        oc8051_ram_top1_oc8051_idata_n75), .B(
        oc8051_ram_top1_oc8051_idata_n525), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4267) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u450 ( .A(
        oc8051_ram_top1_oc8051_idata_n74), .B(
        oc8051_ram_top1_oc8051_idata_n542), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4268) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u449 ( .A(
        oc8051_ram_top1_oc8051_idata_n73), .B(
        oc8051_ram_top1_oc8051_idata_n559), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4269) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u448 ( .A(
        oc8051_ram_top1_oc8051_idata_n72), .B(
        oc8051_ram_top1_oc8051_idata_n576), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4270) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u447 ( .A(
        oc8051_ram_top1_oc8051_idata_n71), .B(
        oc8051_ram_top1_oc8051_idata_n593), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4271) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u446 ( .A(
        oc8051_ram_top1_oc8051_idata_n70), .B(
        oc8051_ram_top1_oc8051_idata_n610), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4272) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u445 ( .A(
        oc8051_ram_top1_oc8051_idata_n69), .B(
        oc8051_ram_top1_oc8051_idata_n627), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4273) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u444 ( .A(
        oc8051_ram_top1_oc8051_idata_n68), .B(
        oc8051_ram_top1_oc8051_idata_n644), .S0(
        oc8051_ram_top1_oc8051_idata_n702), .Y(
        oc8051_ram_top1_oc8051_idata_n4274) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u443 ( .A(
        oc8051_ram_top1_oc8051_idata_n701), .B(
        oc8051_ram_top1_oc8051_idata_n682), .Y(
        oc8051_ram_top1_oc8051_idata_n685) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u442 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n681), .Y(
        oc8051_ram_top1_oc8051_idata_n700) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u441 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4275) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u440 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4276) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u439 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4277) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u438 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4278) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u437 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4279) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u436 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4280) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u435 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4281) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u434 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_31__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n700), .Y(
        oc8051_ram_top1_oc8051_idata_n4282) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u433 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n679), .Y(
        oc8051_ram_top1_oc8051_idata_n699) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u432 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4283) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u431 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4284) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u430 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4285) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u429 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4286) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u428 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4287) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u427 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4288) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u426 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4289) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u425 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_30__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n699), .Y(
        oc8051_ram_top1_oc8051_idata_n4290) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u424 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n677), .Y(
        oc8051_ram_top1_oc8051_idata_n698) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u423 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4291) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u422 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4292) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u421 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4293) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u420 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4294) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u419 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4295) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u418 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4296) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u417 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4297) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u416 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_29__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n698), .Y(
        oc8051_ram_top1_oc8051_idata_n4298) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u415 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n675), .Y(
        oc8051_ram_top1_oc8051_idata_n697) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u414 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4299) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u413 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4300) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u412 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4301) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u411 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4302) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u410 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4303) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u409 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4304) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u408 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4305) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u407 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_28__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n697), .Y(
        oc8051_ram_top1_oc8051_idata_n4306) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u406 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n673), .Y(
        oc8051_ram_top1_oc8051_idata_n696) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u405 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4307) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u404 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4308) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u403 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4309) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u402 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4310) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u401 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4311) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u400 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4312) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u399 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4313) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u398 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_27__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n696), .Y(
        oc8051_ram_top1_oc8051_idata_n4314) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u397 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n671), .Y(
        oc8051_ram_top1_oc8051_idata_n695) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u396 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4315) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u395 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4316) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u394 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4317) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u393 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4318) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u392 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4319) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u391 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4320) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u390 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4321) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u389 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_26__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n695), .Y(
        oc8051_ram_top1_oc8051_idata_n4322) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u388 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n669), .Y(
        oc8051_ram_top1_oc8051_idata_n694) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u387 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4323) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u386 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4324) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u385 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4325) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u384 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4326) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u383 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4327) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u382 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4328) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u381 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4329) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u380 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_25__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n694), .Y(
        oc8051_ram_top1_oc8051_idata_n4330) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u379 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n667), .Y(
        oc8051_ram_top1_oc8051_idata_n693) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u378 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4331) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u377 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4332) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u376 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4333) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u375 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4334) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u374 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4335) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u373 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4336) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u372 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4337) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u371 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_24__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n693), .Y(
        oc8051_ram_top1_oc8051_idata_n4338) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u370 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n665), .Y(
        oc8051_ram_top1_oc8051_idata_n692) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u369 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4339) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u368 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4340) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u367 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4341) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u366 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4342) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u365 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4343) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u364 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4344) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u363 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4345) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u362 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_23__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n692), .Y(
        oc8051_ram_top1_oc8051_idata_n4346) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u361 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n663), .Y(
        oc8051_ram_top1_oc8051_idata_n691) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u360 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4347) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u359 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4348) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u358 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4349) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u357 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4350) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u356 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4351) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u355 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4352) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u354 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4353) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u353 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_22__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n691), .Y(
        oc8051_ram_top1_oc8051_idata_n4354) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u352 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n661), .Y(
        oc8051_ram_top1_oc8051_idata_n690) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u351 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__0_), .B(
        oc8051_ram_top1_oc8051_idata_n2), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4355) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u350 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__1_), .B(
        oc8051_ram_top1_oc8051_idata_n531), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4356) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u349 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__2_), .B(
        oc8051_ram_top1_oc8051_idata_n548), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4357) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u348 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__3_), .B(
        oc8051_ram_top1_oc8051_idata_n565), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4358) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u347 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__4_), .B(
        oc8051_ram_top1_oc8051_idata_n582), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4359) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u346 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__5_), .B(
        oc8051_ram_top1_oc8051_idata_n599), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4360) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u345 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__6_), .B(
        oc8051_ram_top1_oc8051_idata_n616), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4361) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u344 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_21__7_), .B(
        oc8051_ram_top1_oc8051_idata_n633), .S0(
        oc8051_ram_top1_oc8051_idata_n690), .Y(
        oc8051_ram_top1_oc8051_idata_n4362) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u343 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n659), .Y(
        oc8051_ram_top1_oc8051_idata_n689) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u342 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4363) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u341 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4364) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u340 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4365) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u339 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4366) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u338 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4367) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u337 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4368) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u336 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4369) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u335 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_20__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n689), .Y(
        oc8051_ram_top1_oc8051_idata_n4370) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u334 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n657), .Y(
        oc8051_ram_top1_oc8051_idata_n688) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u333 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4371) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u332 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4372) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u331 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4373) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u330 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4374) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u329 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4375) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u328 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4376) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u327 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4377) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u326 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_19__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n688), .Y(
        oc8051_ram_top1_oc8051_idata_n4378) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u325 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n655), .Y(
        oc8051_ram_top1_oc8051_idata_n687) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u324 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4379) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u323 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4380) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u322 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4381) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u321 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4382) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u320 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4383) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u319 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4384) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u318 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4385) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u317 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_18__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n687), .Y(
        oc8051_ram_top1_oc8051_idata_n4386) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u316 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n653), .Y(
        oc8051_ram_top1_oc8051_idata_n686) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u315 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4387) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u314 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4388) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u313 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4389) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u312 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4390) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u311 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4391) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u310 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4392) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u309 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4393) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u308 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_17__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n686), .Y(
        oc8051_ram_top1_oc8051_idata_n4394) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u307 ( .A(
        oc8051_ram_top1_oc8051_idata_n685), .B(
        oc8051_ram_top1_oc8051_idata_n650), .Y(
        oc8051_ram_top1_oc8051_idata_n684) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u306 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4395) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u305 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4396) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u304 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4397) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u303 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4398) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u302 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4399) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u301 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4400) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u300 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4401) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u299 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_16__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n684), .Y(
        oc8051_ram_top1_oc8051_idata_n4402) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u298 ( .A(
        oc8051_ram_top1_oc8051_idata_n682), .B(
        oc8051_ram_top1_oc8051_idata_n683), .Y(
        oc8051_ram_top1_oc8051_idata_n651) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u297 ( .A(
        oc8051_ram_top1_oc8051_idata_n681), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n680) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u296 ( .A(
        oc8051_ram_top1_oc8051_idata_n67), .B(
        oc8051_ram_top1_oc8051_idata_n525), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4403) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u295 ( .A(
        oc8051_ram_top1_oc8051_idata_n66), .B(
        oc8051_ram_top1_oc8051_idata_n542), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4404) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u294 ( .A(
        oc8051_ram_top1_oc8051_idata_n65), .B(
        oc8051_ram_top1_oc8051_idata_n559), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4405) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u293 ( .A(
        oc8051_ram_top1_oc8051_idata_n64), .B(
        oc8051_ram_top1_oc8051_idata_n576), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4406) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u292 ( .A(
        oc8051_ram_top1_oc8051_idata_n63), .B(
        oc8051_ram_top1_oc8051_idata_n593), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4407) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u291 ( .A(
        oc8051_ram_top1_oc8051_idata_n62), .B(
        oc8051_ram_top1_oc8051_idata_n610), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4408) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u290 ( .A(
        oc8051_ram_top1_oc8051_idata_n61), .B(
        oc8051_ram_top1_oc8051_idata_n627), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4409) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u289 ( .A(
        oc8051_ram_top1_oc8051_idata_n60), .B(
        oc8051_ram_top1_oc8051_idata_n644), .S0(
        oc8051_ram_top1_oc8051_idata_n680), .Y(
        oc8051_ram_top1_oc8051_idata_n4410) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u288 ( .A(
        oc8051_ram_top1_oc8051_idata_n679), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n678) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u287 ( .A(
        oc8051_ram_top1_oc8051_idata_n59), .B(
        oc8051_ram_top1_oc8051_idata_n524), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4411) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u286 ( .A(
        oc8051_ram_top1_oc8051_idata_n58), .B(
        oc8051_ram_top1_oc8051_idata_n541), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4412) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u285 ( .A(
        oc8051_ram_top1_oc8051_idata_n57), .B(
        oc8051_ram_top1_oc8051_idata_n558), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4413) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u284 ( .A(
        oc8051_ram_top1_oc8051_idata_n56), .B(
        oc8051_ram_top1_oc8051_idata_n575), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4414) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u283 ( .A(
        oc8051_ram_top1_oc8051_idata_n55), .B(
        oc8051_ram_top1_oc8051_idata_n592), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4415) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u282 ( .A(
        oc8051_ram_top1_oc8051_idata_n54), .B(
        oc8051_ram_top1_oc8051_idata_n609), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4416) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u281 ( .A(
        oc8051_ram_top1_oc8051_idata_n53), .B(
        oc8051_ram_top1_oc8051_idata_n626), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4417) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u280 ( .A(
        oc8051_ram_top1_oc8051_idata_n52), .B(
        oc8051_ram_top1_oc8051_idata_n643), .S0(
        oc8051_ram_top1_oc8051_idata_n678), .Y(
        oc8051_ram_top1_oc8051_idata_n4418) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u279 ( .A(
        oc8051_ram_top1_oc8051_idata_n677), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n676) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u278 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4419) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u277 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4420) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u276 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4421) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u275 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4422) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u274 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4423) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u273 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4424) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u272 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4425) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u271 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_13__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n676), .Y(
        oc8051_ram_top1_oc8051_idata_n4426) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u270 ( .A(
        oc8051_ram_top1_oc8051_idata_n675), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n674) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u269 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4427) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u268 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4428) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u267 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4429) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u266 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4430) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u265 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4431) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u264 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4432) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u263 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4433) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u262 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_12__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n674), .Y(
        oc8051_ram_top1_oc8051_idata_n4434) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u261 ( .A(
        oc8051_ram_top1_oc8051_idata_n673), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n672) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u260 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4435) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u259 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4436) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u258 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4437) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u257 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4438) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u256 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4439) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u255 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4440) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u254 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4441) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u253 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_11__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n672), .Y(
        oc8051_ram_top1_oc8051_idata_n4442) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u252 ( .A(
        oc8051_ram_top1_oc8051_idata_n671), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n670) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u251 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4443) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u250 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4444) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u249 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4445) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u248 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4446) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u247 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4447) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u246 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4448) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u245 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4449) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u244 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_10__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n670), .Y(
        oc8051_ram_top1_oc8051_idata_n4450) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u243 ( .A(
        oc8051_ram_top1_oc8051_idata_n669), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n668) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u242 ( .A(
        oc8051_ram_top1_oc8051_idata_n51), .B(
        oc8051_ram_top1_oc8051_idata_n524), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4451) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u241 ( .A(
        oc8051_ram_top1_oc8051_idata_n50), .B(
        oc8051_ram_top1_oc8051_idata_n541), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4452) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u240 ( .A(
        oc8051_ram_top1_oc8051_idata_n49), .B(
        oc8051_ram_top1_oc8051_idata_n558), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4453) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u239 ( .A(
        oc8051_ram_top1_oc8051_idata_n48), .B(
        oc8051_ram_top1_oc8051_idata_n575), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4454) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u238 ( .A(
        oc8051_ram_top1_oc8051_idata_n47), .B(
        oc8051_ram_top1_oc8051_idata_n592), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4455) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u237 ( .A(
        oc8051_ram_top1_oc8051_idata_n46), .B(
        oc8051_ram_top1_oc8051_idata_n609), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4456) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u236 ( .A(
        oc8051_ram_top1_oc8051_idata_n45), .B(
        oc8051_ram_top1_oc8051_idata_n626), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4457) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u235 ( .A(
        oc8051_ram_top1_oc8051_idata_n44), .B(
        oc8051_ram_top1_oc8051_idata_n643), .S0(
        oc8051_ram_top1_oc8051_idata_n668), .Y(
        oc8051_ram_top1_oc8051_idata_n4458) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u234 ( .A(
        oc8051_ram_top1_oc8051_idata_n667), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n666) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u233 ( .A(
        oc8051_ram_top1_oc8051_idata_n43), .B(
        oc8051_ram_top1_oc8051_idata_n524), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4459) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u232 ( .A(
        oc8051_ram_top1_oc8051_idata_n42), .B(
        oc8051_ram_top1_oc8051_idata_n541), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4460) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u231 ( .A(
        oc8051_ram_top1_oc8051_idata_n41), .B(
        oc8051_ram_top1_oc8051_idata_n558), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4461) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u230 ( .A(
        oc8051_ram_top1_oc8051_idata_n40), .B(
        oc8051_ram_top1_oc8051_idata_n575), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4462) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u229 ( .A(
        oc8051_ram_top1_oc8051_idata_n39), .B(
        oc8051_ram_top1_oc8051_idata_n592), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4463) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u228 ( .A(
        oc8051_ram_top1_oc8051_idata_n38), .B(
        oc8051_ram_top1_oc8051_idata_n609), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4464) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u227 ( .A(
        oc8051_ram_top1_oc8051_idata_n37), .B(
        oc8051_ram_top1_oc8051_idata_n626), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4465) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u226 ( .A(
        oc8051_ram_top1_oc8051_idata_n36), .B(
        oc8051_ram_top1_oc8051_idata_n643), .S0(
        oc8051_ram_top1_oc8051_idata_n666), .Y(
        oc8051_ram_top1_oc8051_idata_n4466) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u225 ( .A(
        oc8051_ram_top1_oc8051_idata_n665), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n664) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u224 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4467) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u223 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4468) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u222 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4469) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u221 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4470) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u220 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4471) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u219 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4472) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u218 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4473) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u217 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_7__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n664), .Y(
        oc8051_ram_top1_oc8051_idata_n4474) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u216 ( .A(
        oc8051_ram_top1_oc8051_idata_n663), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n662) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u215 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4475) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u214 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4476) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u213 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4477) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u212 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4478) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u211 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4479) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u210 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4480) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u209 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4481) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u208 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_6__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n662), .Y(
        oc8051_ram_top1_oc8051_idata_n4482) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u207 ( .A(
        oc8051_ram_top1_oc8051_idata_n661), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n660) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u206 ( .A(
        oc8051_ram_top1_oc8051_idata_n35), .B(
        oc8051_ram_top1_oc8051_idata_n523), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4483) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u205 ( .A(
        oc8051_ram_top1_oc8051_idata_n34), .B(
        oc8051_ram_top1_oc8051_idata_n540), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4484) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u204 ( .A(
        oc8051_ram_top1_oc8051_idata_n33), .B(
        oc8051_ram_top1_oc8051_idata_n557), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4485) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u203 ( .A(
        oc8051_ram_top1_oc8051_idata_n32), .B(
        oc8051_ram_top1_oc8051_idata_n574), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4486) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u202 ( .A(
        oc8051_ram_top1_oc8051_idata_n31), .B(
        oc8051_ram_top1_oc8051_idata_n591), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4487) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u201 ( .A(
        oc8051_ram_top1_oc8051_idata_n30), .B(
        oc8051_ram_top1_oc8051_idata_n608), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4488) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u200 ( .A(
        oc8051_ram_top1_oc8051_idata_n29), .B(
        oc8051_ram_top1_oc8051_idata_n625), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4489) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u199 ( .A(
        oc8051_ram_top1_oc8051_idata_n28), .B(
        oc8051_ram_top1_oc8051_idata_n642), .S0(
        oc8051_ram_top1_oc8051_idata_n660), .Y(
        oc8051_ram_top1_oc8051_idata_n4490) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u198 ( .A(
        oc8051_ram_top1_oc8051_idata_n659), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n658) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u197 ( .A(
        oc8051_ram_top1_oc8051_idata_n27), .B(
        oc8051_ram_top1_oc8051_idata_n523), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4491) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u196 ( .A(
        oc8051_ram_top1_oc8051_idata_n26), .B(
        oc8051_ram_top1_oc8051_idata_n540), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4492) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u195 ( .A(
        oc8051_ram_top1_oc8051_idata_n25), .B(
        oc8051_ram_top1_oc8051_idata_n557), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4493) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u194 ( .A(
        oc8051_ram_top1_oc8051_idata_n24), .B(
        oc8051_ram_top1_oc8051_idata_n574), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4494) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u193 ( .A(
        oc8051_ram_top1_oc8051_idata_n23), .B(
        oc8051_ram_top1_oc8051_idata_n591), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4495) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u192 ( .A(
        oc8051_ram_top1_oc8051_idata_n22), .B(
        oc8051_ram_top1_oc8051_idata_n608), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4496) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u191 ( .A(
        oc8051_ram_top1_oc8051_idata_n21), .B(
        oc8051_ram_top1_oc8051_idata_n625), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4497) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u190 ( .A(
        oc8051_ram_top1_oc8051_idata_n20), .B(
        oc8051_ram_top1_oc8051_idata_n642), .S0(
        oc8051_ram_top1_oc8051_idata_n658), .Y(
        oc8051_ram_top1_oc8051_idata_n4498) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u189 ( .A(
        oc8051_ram_top1_oc8051_idata_n657), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n656) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u188 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4499) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u187 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4500) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u186 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4501) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u185 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4502) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u184 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4503) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u183 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4504) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u182 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4505) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u181 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_3__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n656), .Y(
        oc8051_ram_top1_oc8051_idata_n4506) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u180 ( .A(
        oc8051_ram_top1_oc8051_idata_n655), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n654) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u179 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__0_), .B(
        oc8051_ram_top1_oc8051_idata_n1), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4507) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u178 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__1_), .B(
        oc8051_ram_top1_oc8051_idata_n530), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4508) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u177 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__2_), .B(
        oc8051_ram_top1_oc8051_idata_n547), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4509) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u176 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__3_), .B(
        oc8051_ram_top1_oc8051_idata_n564), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4510) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u175 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__4_), .B(
        oc8051_ram_top1_oc8051_idata_n581), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4511) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u174 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__5_), .B(
        oc8051_ram_top1_oc8051_idata_n598), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4512) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u173 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__6_), .B(
        oc8051_ram_top1_oc8051_idata_n615), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4513) );
  MXT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u172 ( .A(
        oc8051_ram_top1_oc8051_idata_buff_2__7_), .B(
        oc8051_ram_top1_oc8051_idata_n632), .S0(
        oc8051_ram_top1_oc8051_idata_n654), .Y(
        oc8051_ram_top1_oc8051_idata_n4514) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u171 ( .A(
        oc8051_ram_top1_oc8051_idata_n653), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n652) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u170 ( .A(
        oc8051_ram_top1_oc8051_idata_n19), .B(
        oc8051_ram_top1_oc8051_idata_n523), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4515) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u169 ( .A(
        oc8051_ram_top1_oc8051_idata_n18), .B(
        oc8051_ram_top1_oc8051_idata_n540), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4516) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u168 ( .A(
        oc8051_ram_top1_oc8051_idata_n17), .B(
        oc8051_ram_top1_oc8051_idata_n557), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4517) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u167 ( .A(
        oc8051_ram_top1_oc8051_idata_n16), .B(
        oc8051_ram_top1_oc8051_idata_n574), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4518) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u166 ( .A(
        oc8051_ram_top1_oc8051_idata_n15), .B(
        oc8051_ram_top1_oc8051_idata_n591), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4519) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u165 ( .A(
        oc8051_ram_top1_oc8051_idata_n14), .B(
        oc8051_ram_top1_oc8051_idata_n608), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4520) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u164 ( .A(
        oc8051_ram_top1_oc8051_idata_n13), .B(
        oc8051_ram_top1_oc8051_idata_n625), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4521) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u163 ( .A(
        oc8051_ram_top1_oc8051_idata_n12), .B(
        oc8051_ram_top1_oc8051_idata_n642), .S0(
        oc8051_ram_top1_oc8051_idata_n652), .Y(
        oc8051_ram_top1_oc8051_idata_n4522) );
  AND2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u162 ( .A(
        oc8051_ram_top1_oc8051_idata_n650), .B(
        oc8051_ram_top1_oc8051_idata_n651), .Y(
        oc8051_ram_top1_oc8051_idata_n649) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u161 ( .A(
        oc8051_ram_top1_oc8051_idata_n11), .B(
        oc8051_ram_top1_oc8051_idata_n528), .S0(
        oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4523) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u160 ( .A(
        oc8051_ram_top1_oc8051_idata_n10), .B(
        oc8051_ram_top1_oc8051_idata_n545), .S0(
        oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4524) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u159 ( .A(
        oc8051_ram_top1_oc8051_idata_n9), .B(oc8051_ram_top1_oc8051_idata_n562), .S0(oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4525) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u158 ( .A(
        oc8051_ram_top1_oc8051_idata_n8), .B(oc8051_ram_top1_oc8051_idata_n579), .S0(oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4526) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u157 ( .A(
        oc8051_ram_top1_oc8051_idata_n7), .B(oc8051_ram_top1_oc8051_idata_n596), .S0(oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4527) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u156 ( .A(
        oc8051_ram_top1_oc8051_idata_n6), .B(oc8051_ram_top1_oc8051_idata_n613), .S0(oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4528) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u155 ( .A(
        oc8051_ram_top1_oc8051_idata_n5), .B(oc8051_ram_top1_oc8051_idata_n630), .S0(oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4529) );
  MXIT2_X0P5M_A12TS oc8051_ram_top1_oc8051_idata_u154 ( .A(
        oc8051_ram_top1_oc8051_idata_n4), .B(oc8051_ram_top1_oc8051_idata_n647), .S0(oc8051_ram_top1_oc8051_idata_n649), .Y(
        oc8051_ram_top1_oc8051_idata_n4530) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u153 ( .A(oc8051_ram_top1_n3), 
        .Y(oc8051_ram_top1_oc8051_idata_n563) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u152 ( .A(oc8051_ram_top1_n1), 
        .Y(oc8051_ram_top1_oc8051_idata_n529) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u151 ( .A(oc8051_ram_top1_n2), 
        .Y(oc8051_ram_top1_oc8051_idata_n546) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u150 ( .A(oc8051_ram_top1_n7), 
        .Y(oc8051_ram_top1_oc8051_idata_n631) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u149 ( .A(oc8051_ram_top1_n6), 
        .Y(oc8051_ram_top1_oc8051_idata_n614) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u148 ( .A(oc8051_ram_top1_n5), 
        .Y(oc8051_ram_top1_oc8051_idata_n597) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u147 ( .A(oc8051_ram_top1_n4), 
        .Y(oc8051_ram_top1_oc8051_idata_n580) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u146 ( .A(oc8051_ram_top1_n8), 
        .Y(oc8051_ram_top1_oc8051_idata_n648) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u145 ( .A(
        oc8051_ram_top1_oc8051_idata_n648), .Y(
        oc8051_ram_top1_oc8051_idata_n647) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u144 ( .A(
        oc8051_ram_top1_oc8051_idata_n631), .Y(
        oc8051_ram_top1_oc8051_idata_n630) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u143 ( .A(
        oc8051_ram_top1_oc8051_idata_n614), .Y(
        oc8051_ram_top1_oc8051_idata_n613) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u142 ( .A(
        oc8051_ram_top1_oc8051_idata_n597), .Y(
        oc8051_ram_top1_oc8051_idata_n596) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u141 ( .A(
        oc8051_ram_top1_oc8051_idata_n580), .Y(
        oc8051_ram_top1_oc8051_idata_n579) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u140 ( .A(
        oc8051_ram_top1_oc8051_idata_n563), .Y(
        oc8051_ram_top1_oc8051_idata_n562) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u139 ( .A(
        oc8051_ram_top1_oc8051_idata_n546), .Y(
        oc8051_ram_top1_oc8051_idata_n545) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u138 ( .A(
        oc8051_ram_top1_oc8051_idata_n529), .Y(
        oc8051_ram_top1_oc8051_idata_n528) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u137 ( .A(
        oc8051_ram_top1_oc8051_idata_n648), .Y(
        oc8051_ram_top1_oc8051_idata_n646) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u136 ( .A(
        oc8051_ram_top1_oc8051_idata_n631), .Y(
        oc8051_ram_top1_oc8051_idata_n629) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u135 ( .A(
        oc8051_ram_top1_oc8051_idata_n614), .Y(
        oc8051_ram_top1_oc8051_idata_n612) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u134 ( .A(
        oc8051_ram_top1_oc8051_idata_n597), .Y(
        oc8051_ram_top1_oc8051_idata_n595) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u133 ( .A(
        oc8051_ram_top1_oc8051_idata_n580), .Y(
        oc8051_ram_top1_oc8051_idata_n578) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u132 ( .A(
        oc8051_ram_top1_oc8051_idata_n563), .Y(
        oc8051_ram_top1_oc8051_idata_n561) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u131 ( .A(
        oc8051_ram_top1_oc8051_idata_n546), .Y(
        oc8051_ram_top1_oc8051_idata_n544) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u130 ( .A(
        oc8051_ram_top1_oc8051_idata_n529), .Y(
        oc8051_ram_top1_oc8051_idata_n527) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u129 ( .A(
        oc8051_ram_top1_oc8051_idata_n648), .Y(
        oc8051_ram_top1_oc8051_idata_n642) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u128 ( .A(
        oc8051_ram_top1_oc8051_idata_n631), .Y(
        oc8051_ram_top1_oc8051_idata_n625) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u127 ( .A(
        oc8051_ram_top1_oc8051_idata_n614), .Y(
        oc8051_ram_top1_oc8051_idata_n608) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u126 ( .A(
        oc8051_ram_top1_oc8051_idata_n597), .Y(
        oc8051_ram_top1_oc8051_idata_n591) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u125 ( .A(
        oc8051_ram_top1_oc8051_idata_n580), .Y(
        oc8051_ram_top1_oc8051_idata_n574) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u124 ( .A(
        oc8051_ram_top1_oc8051_idata_n563), .Y(
        oc8051_ram_top1_oc8051_idata_n557) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u123 ( .A(
        oc8051_ram_top1_oc8051_idata_n546), .Y(
        oc8051_ram_top1_oc8051_idata_n540) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u122 ( .A(
        oc8051_ram_top1_oc8051_idata_n529), .Y(
        oc8051_ram_top1_oc8051_idata_n523) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u121 ( .A(
        oc8051_ram_top1_oc8051_idata_n648), .Y(
        oc8051_ram_top1_oc8051_idata_n643) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u120 ( .A(
        oc8051_ram_top1_oc8051_idata_n631), .Y(
        oc8051_ram_top1_oc8051_idata_n626) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u119 ( .A(
        oc8051_ram_top1_oc8051_idata_n614), .Y(
        oc8051_ram_top1_oc8051_idata_n609) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u118 ( .A(
        oc8051_ram_top1_oc8051_idata_n597), .Y(
        oc8051_ram_top1_oc8051_idata_n592) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u117 ( .A(
        oc8051_ram_top1_oc8051_idata_n580), .Y(
        oc8051_ram_top1_oc8051_idata_n575) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u116 ( .A(
        oc8051_ram_top1_oc8051_idata_n563), .Y(
        oc8051_ram_top1_oc8051_idata_n558) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u115 ( .A(
        oc8051_ram_top1_oc8051_idata_n546), .Y(
        oc8051_ram_top1_oc8051_idata_n541) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u114 ( .A(
        oc8051_ram_top1_oc8051_idata_n529), .Y(
        oc8051_ram_top1_oc8051_idata_n524) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u113 ( .A(
        oc8051_ram_top1_oc8051_idata_n648), .Y(
        oc8051_ram_top1_oc8051_idata_n644) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u112 ( .A(
        oc8051_ram_top1_oc8051_idata_n631), .Y(
        oc8051_ram_top1_oc8051_idata_n627) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u111 ( .A(
        oc8051_ram_top1_oc8051_idata_n614), .Y(
        oc8051_ram_top1_oc8051_idata_n610) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u110 ( .A(
        oc8051_ram_top1_oc8051_idata_n597), .Y(
        oc8051_ram_top1_oc8051_idata_n593) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u109 ( .A(
        oc8051_ram_top1_oc8051_idata_n580), .Y(
        oc8051_ram_top1_oc8051_idata_n576) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u108 ( .A(
        oc8051_ram_top1_oc8051_idata_n563), .Y(
        oc8051_ram_top1_oc8051_idata_n559) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u107 ( .A(
        oc8051_ram_top1_oc8051_idata_n546), .Y(
        oc8051_ram_top1_oc8051_idata_n542) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u106 ( .A(
        oc8051_ram_top1_oc8051_idata_n529), .Y(
        oc8051_ram_top1_oc8051_idata_n525) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u105 ( .A(
        oc8051_ram_top1_oc8051_idata_n648), .Y(
        oc8051_ram_top1_oc8051_idata_n645) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u104 ( .A(
        oc8051_ram_top1_oc8051_idata_n631), .Y(
        oc8051_ram_top1_oc8051_idata_n628) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u103 ( .A(
        oc8051_ram_top1_oc8051_idata_n614), .Y(
        oc8051_ram_top1_oc8051_idata_n611) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u102 ( .A(
        oc8051_ram_top1_oc8051_idata_n597), .Y(
        oc8051_ram_top1_oc8051_idata_n594) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u101 ( .A(
        oc8051_ram_top1_oc8051_idata_n580), .Y(
        oc8051_ram_top1_oc8051_idata_n577) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u100 ( .A(
        oc8051_ram_top1_oc8051_idata_n563), .Y(
        oc8051_ram_top1_oc8051_idata_n560) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u99 ( .A(
        oc8051_ram_top1_oc8051_idata_n546), .Y(
        oc8051_ram_top1_oc8051_idata_n543) );
  BUFH_X1M_A12TS oc8051_ram_top1_oc8051_idata_u98 ( .A(
        oc8051_ram_top1_oc8051_idata_n529), .Y(
        oc8051_ram_top1_oc8051_idata_n526) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u97 ( .A(
        oc8051_ram_top1_oc8051_idata_n646), .Y(
        oc8051_ram_top1_oc8051_idata_n632) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u96 ( .A(
        oc8051_ram_top1_oc8051_idata_n629), .Y(
        oc8051_ram_top1_oc8051_idata_n615) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u95 ( .A(
        oc8051_ram_top1_oc8051_idata_n612), .Y(
        oc8051_ram_top1_oc8051_idata_n598) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u94 ( .A(
        oc8051_ram_top1_oc8051_idata_n595), .Y(
        oc8051_ram_top1_oc8051_idata_n581) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u93 ( .A(
        oc8051_ram_top1_oc8051_idata_n578), .Y(
        oc8051_ram_top1_oc8051_idata_n564) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u92 ( .A(
        oc8051_ram_top1_oc8051_idata_n561), .Y(
        oc8051_ram_top1_oc8051_idata_n547) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u91 ( .A(
        oc8051_ram_top1_oc8051_idata_n544), .Y(
        oc8051_ram_top1_oc8051_idata_n530) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u90 ( .A(
        oc8051_ram_top1_oc8051_idata_n527), .Y(oc8051_ram_top1_oc8051_idata_n1) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u89 ( .A(
        oc8051_ram_top1_oc8051_idata_n646), .Y(
        oc8051_ram_top1_oc8051_idata_n633) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u88 ( .A(
        oc8051_ram_top1_oc8051_idata_n629), .Y(
        oc8051_ram_top1_oc8051_idata_n616) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u87 ( .A(
        oc8051_ram_top1_oc8051_idata_n612), .Y(
        oc8051_ram_top1_oc8051_idata_n599) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u86 ( .A(
        oc8051_ram_top1_oc8051_idata_n595), .Y(
        oc8051_ram_top1_oc8051_idata_n582) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u85 ( .A(
        oc8051_ram_top1_oc8051_idata_n578), .Y(
        oc8051_ram_top1_oc8051_idata_n565) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u84 ( .A(
        oc8051_ram_top1_oc8051_idata_n561), .Y(
        oc8051_ram_top1_oc8051_idata_n548) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u83 ( .A(
        oc8051_ram_top1_oc8051_idata_n544), .Y(
        oc8051_ram_top1_oc8051_idata_n531) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u82 ( .A(
        oc8051_ram_top1_oc8051_idata_n527), .Y(oc8051_ram_top1_oc8051_idata_n2) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u81 ( .A(
        oc8051_ram_top1_oc8051_idata_n645), .Y(
        oc8051_ram_top1_oc8051_idata_n634) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u80 ( .A(
        oc8051_ram_top1_oc8051_idata_n628), .Y(
        oc8051_ram_top1_oc8051_idata_n617) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u79 ( .A(
        oc8051_ram_top1_oc8051_idata_n611), .Y(
        oc8051_ram_top1_oc8051_idata_n600) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u78 ( .A(
        oc8051_ram_top1_oc8051_idata_n594), .Y(
        oc8051_ram_top1_oc8051_idata_n583) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u77 ( .A(
        oc8051_ram_top1_oc8051_idata_n577), .Y(
        oc8051_ram_top1_oc8051_idata_n566) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u76 ( .A(
        oc8051_ram_top1_oc8051_idata_n560), .Y(
        oc8051_ram_top1_oc8051_idata_n549) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u75 ( .A(
        oc8051_ram_top1_oc8051_idata_n543), .Y(
        oc8051_ram_top1_oc8051_idata_n532) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u74 ( .A(
        oc8051_ram_top1_oc8051_idata_n526), .Y(oc8051_ram_top1_oc8051_idata_n3) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u73 ( .A(
        oc8051_ram_top1_oc8051_idata_n645), .Y(
        oc8051_ram_top1_oc8051_idata_n635) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u72 ( .A(
        oc8051_ram_top1_oc8051_idata_n628), .Y(
        oc8051_ram_top1_oc8051_idata_n618) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u71 ( .A(
        oc8051_ram_top1_oc8051_idata_n611), .Y(
        oc8051_ram_top1_oc8051_idata_n601) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u70 ( .A(
        oc8051_ram_top1_oc8051_idata_n594), .Y(
        oc8051_ram_top1_oc8051_idata_n584) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u69 ( .A(
        oc8051_ram_top1_oc8051_idata_n577), .Y(
        oc8051_ram_top1_oc8051_idata_n567) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u68 ( .A(
        oc8051_ram_top1_oc8051_idata_n560), .Y(
        oc8051_ram_top1_oc8051_idata_n550) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u67 ( .A(
        oc8051_ram_top1_oc8051_idata_n543), .Y(
        oc8051_ram_top1_oc8051_idata_n533) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u66 ( .A(
        oc8051_ram_top1_oc8051_idata_n526), .Y(
        oc8051_ram_top1_oc8051_idata_n516) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u65 ( .A(
        oc8051_ram_top1_oc8051_idata_n645), .Y(
        oc8051_ram_top1_oc8051_idata_n636) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u64 ( .A(
        oc8051_ram_top1_oc8051_idata_n628), .Y(
        oc8051_ram_top1_oc8051_idata_n619) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u63 ( .A(
        oc8051_ram_top1_oc8051_idata_n611), .Y(
        oc8051_ram_top1_oc8051_idata_n602) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u62 ( .A(
        oc8051_ram_top1_oc8051_idata_n594), .Y(
        oc8051_ram_top1_oc8051_idata_n585) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u61 ( .A(
        oc8051_ram_top1_oc8051_idata_n577), .Y(
        oc8051_ram_top1_oc8051_idata_n568) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u60 ( .A(
        oc8051_ram_top1_oc8051_idata_n560), .Y(
        oc8051_ram_top1_oc8051_idata_n551) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u59 ( .A(
        oc8051_ram_top1_oc8051_idata_n543), .Y(
        oc8051_ram_top1_oc8051_idata_n534) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u58 ( .A(
        oc8051_ram_top1_oc8051_idata_n526), .Y(
        oc8051_ram_top1_oc8051_idata_n517) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u57 ( .A(
        oc8051_ram_top1_oc8051_idata_n644), .Y(
        oc8051_ram_top1_oc8051_idata_n637) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u56 ( .A(
        oc8051_ram_top1_oc8051_idata_n627), .Y(
        oc8051_ram_top1_oc8051_idata_n620) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u55 ( .A(
        oc8051_ram_top1_oc8051_idata_n610), .Y(
        oc8051_ram_top1_oc8051_idata_n603) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u54 ( .A(
        oc8051_ram_top1_oc8051_idata_n593), .Y(
        oc8051_ram_top1_oc8051_idata_n586) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u53 ( .A(
        oc8051_ram_top1_oc8051_idata_n576), .Y(
        oc8051_ram_top1_oc8051_idata_n569) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u52 ( .A(
        oc8051_ram_top1_oc8051_idata_n559), .Y(
        oc8051_ram_top1_oc8051_idata_n552) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u51 ( .A(
        oc8051_ram_top1_oc8051_idata_n542), .Y(
        oc8051_ram_top1_oc8051_idata_n535) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u50 ( .A(
        oc8051_ram_top1_oc8051_idata_n525), .Y(
        oc8051_ram_top1_oc8051_idata_n518) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u49 ( .A(
        oc8051_ram_top1_oc8051_idata_n644), .Y(
        oc8051_ram_top1_oc8051_idata_n638) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u48 ( .A(
        oc8051_ram_top1_oc8051_idata_n627), .Y(
        oc8051_ram_top1_oc8051_idata_n621) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u47 ( .A(
        oc8051_ram_top1_oc8051_idata_n610), .Y(
        oc8051_ram_top1_oc8051_idata_n604) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u46 ( .A(
        oc8051_ram_top1_oc8051_idata_n593), .Y(
        oc8051_ram_top1_oc8051_idata_n587) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u45 ( .A(
        oc8051_ram_top1_oc8051_idata_n576), .Y(
        oc8051_ram_top1_oc8051_idata_n570) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u44 ( .A(
        oc8051_ram_top1_oc8051_idata_n559), .Y(
        oc8051_ram_top1_oc8051_idata_n553) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u43 ( .A(
        oc8051_ram_top1_oc8051_idata_n542), .Y(
        oc8051_ram_top1_oc8051_idata_n536) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u42 ( .A(
        oc8051_ram_top1_oc8051_idata_n525), .Y(
        oc8051_ram_top1_oc8051_idata_n519) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u41 ( .A(
        oc8051_ram_top1_oc8051_idata_n644), .Y(
        oc8051_ram_top1_oc8051_idata_n639) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u40 ( .A(
        oc8051_ram_top1_oc8051_idata_n627), .Y(
        oc8051_ram_top1_oc8051_idata_n622) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u39 ( .A(
        oc8051_ram_top1_oc8051_idata_n610), .Y(
        oc8051_ram_top1_oc8051_idata_n605) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u38 ( .A(
        oc8051_ram_top1_oc8051_idata_n593), .Y(
        oc8051_ram_top1_oc8051_idata_n588) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u37 ( .A(
        oc8051_ram_top1_oc8051_idata_n576), .Y(
        oc8051_ram_top1_oc8051_idata_n571) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u36 ( .A(
        oc8051_ram_top1_oc8051_idata_n559), .Y(
        oc8051_ram_top1_oc8051_idata_n554) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u35 ( .A(
        oc8051_ram_top1_oc8051_idata_n542), .Y(
        oc8051_ram_top1_oc8051_idata_n537) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u34 ( .A(
        oc8051_ram_top1_oc8051_idata_n525), .Y(
        oc8051_ram_top1_oc8051_idata_n520) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u33 ( .A(
        oc8051_ram_top1_oc8051_idata_n643), .Y(
        oc8051_ram_top1_oc8051_idata_n640) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u32 ( .A(
        oc8051_ram_top1_oc8051_idata_n626), .Y(
        oc8051_ram_top1_oc8051_idata_n623) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u31 ( .A(
        oc8051_ram_top1_oc8051_idata_n609), .Y(
        oc8051_ram_top1_oc8051_idata_n606) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u30 ( .A(
        oc8051_ram_top1_oc8051_idata_n592), .Y(
        oc8051_ram_top1_oc8051_idata_n589) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u29 ( .A(
        oc8051_ram_top1_oc8051_idata_n575), .Y(
        oc8051_ram_top1_oc8051_idata_n572) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u28 ( .A(
        oc8051_ram_top1_oc8051_idata_n558), .Y(
        oc8051_ram_top1_oc8051_idata_n555) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u27 ( .A(
        oc8051_ram_top1_oc8051_idata_n541), .Y(
        oc8051_ram_top1_oc8051_idata_n538) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u26 ( .A(
        oc8051_ram_top1_oc8051_idata_n524), .Y(
        oc8051_ram_top1_oc8051_idata_n521) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u25 ( .A(
        oc8051_ram_top1_oc8051_idata_n643), .Y(
        oc8051_ram_top1_oc8051_idata_n641) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u24 ( .A(
        oc8051_ram_top1_oc8051_idata_n626), .Y(
        oc8051_ram_top1_oc8051_idata_n624) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u23 ( .A(
        oc8051_ram_top1_oc8051_idata_n609), .Y(
        oc8051_ram_top1_oc8051_idata_n607) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u22 ( .A(
        oc8051_ram_top1_oc8051_idata_n592), .Y(
        oc8051_ram_top1_oc8051_idata_n590) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u21 ( .A(
        oc8051_ram_top1_oc8051_idata_n575), .Y(
        oc8051_ram_top1_oc8051_idata_n573) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u20 ( .A(
        oc8051_ram_top1_oc8051_idata_n558), .Y(
        oc8051_ram_top1_oc8051_idata_n556) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u19 ( .A(
        oc8051_ram_top1_oc8051_idata_n541), .Y(
        oc8051_ram_top1_oc8051_idata_n539) );
  INV_X1M_A12TS oc8051_ram_top1_oc8051_idata_u18 ( .A(
        oc8051_ram_top1_oc8051_idata_n524), .Y(
        oc8051_ram_top1_oc8051_idata_n522) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u17 ( .A(
        oc8051_ram_top1_oc8051_idata_n4594), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n1124) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u16 ( .A(
        oc8051_ram_top1_oc8051_idata_n4627), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1176) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u15 ( .A(
        oc8051_ram_top1_oc8051_idata_n4593), .B(
        oc8051_ram_top1_oc8051_idata_n4588), .Y(
        oc8051_ram_top1_oc8051_idata_n1125) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u14 ( .A(
        oc8051_ram_top1_oc8051_idata_n4627), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1177) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u13 ( .A(
        oc8051_ram_top1_oc8051_idata_n4578), .B(
        oc8051_ram_top1_oc8051_idata_n4579), .Y(
        oc8051_ram_top1_oc8051_idata_n1110) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u12 ( .A(
        oc8051_ram_top1_oc8051_idata_n4615), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1158) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u11 ( .A(
        oc8051_ram_top1_oc8051_idata_n4622), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1170) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u10 ( .A(
        oc8051_ram_top1_oc8051_idata_n4586), .B(
        oc8051_ram_top1_oc8051_idata_n4580), .Y(
        oc8051_ram_top1_oc8051_idata_n1119) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u9 ( .A(
        oc8051_ram_top1_oc8051_idata_n4586), .B(
        oc8051_ram_top1_oc8051_idata_n4579), .Y(
        oc8051_ram_top1_oc8051_idata_n1120) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u8 ( .A(
        oc8051_ram_top1_oc8051_idata_n4618), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1163) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u7 ( .A(
        oc8051_ram_top1_oc8051_idata_n4580), .B(
        oc8051_ram_top1_oc8051_idata_n4578), .Y(
        oc8051_ram_top1_oc8051_idata_n1109) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u6 ( .A(
        oc8051_ram_top1_oc8051_idata_n4615), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1157) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u5 ( .A(
        oc8051_ram_top1_oc8051_idata_n4584), .B(
        oc8051_ram_top1_oc8051_idata_n4579), .Y(
        oc8051_ram_top1_oc8051_idata_n1115) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u4 ( .A(
        oc8051_ram_top1_oc8051_idata_n4618), .B(
        oc8051_ram_top1_oc8051_idata_n4589), .Y(
        oc8051_ram_top1_oc8051_idata_n1162) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u3 ( .A(
        oc8051_ram_top1_oc8051_idata_n4622), .B(
        oc8051_ram_top1_oc8051_idata_n4587), .Y(
        oc8051_ram_top1_oc8051_idata_n1169) );
  NAND2_X1M_A12TS oc8051_ram_top1_oc8051_idata_u2 ( .A(
        oc8051_ram_top1_oc8051_idata_n4584), .B(
        oc8051_ram_top1_oc8051_idata_n4580), .Y(
        oc8051_ram_top1_oc8051_idata_n1114) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2547), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n515) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2548), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n514) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2549), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n513) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2550), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n512) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2551), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n511) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2552), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n510) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2553), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n509) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_247__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2554), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n508) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2555), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n507) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2556), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n506) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2557), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n505) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2558), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n504) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2559), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n503) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2560), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n502) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2561), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n501) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_246__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2562), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n500) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2579), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n499) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2580), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n498) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2581), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n497) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2582), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n496) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2583), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n495) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2584), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n494) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2585), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n493) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_243__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2586), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n492) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2587), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n491) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2588), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n490) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2589), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n489) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2590), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n488) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2591), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n487) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2592), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n486) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2593), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n485) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_242__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2594), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n484) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3059), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n387) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3060), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n386) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3061), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n385) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3062), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n384) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3063), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n383) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3064), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n382) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3065), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n381) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_183__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3066), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n380) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3067), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n379) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3068), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n378) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3069), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n377) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3070), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n376) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3071), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n375) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3072), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n374) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3073), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n373) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_182__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3074), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n372) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3091), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n371) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3092), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n370) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3093), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n369) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3094), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n368) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3095), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n367) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3096), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n366) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3097), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n365) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_179__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3098), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n364) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3099), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n363) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3100), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n362) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3101), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n361) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3102), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n360) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3103), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n359) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3104), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n358) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3105), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n357) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_178__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3106), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n356) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3571), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n259) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3572), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n258) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3573), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n257) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3574), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n256) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3575), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n255) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3576), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n254) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3577), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n253) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_119__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3578), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n252) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3579), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n251) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3580), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n250) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3581), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n249) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3582), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n248) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3583), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n247) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3584), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n246) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3585), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n245) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_118__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3586), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n244) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3603), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n243) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3604), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n242) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3605), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n241) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3606), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n240) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3607), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n239) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3608), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n238) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3609), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n237) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_115__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3610), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n236) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3611), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n235) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3612), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n234) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3613), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n233) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3614), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n232) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3615), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n231) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3616), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n230) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3617), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n229) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_114__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3618), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n228) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4083), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n131) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4084), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n130) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4085), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n129) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4086), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n128) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4087), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n127) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4088), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n126) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4089), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n125) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_55__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4090), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n124) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4091), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n123) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4092), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n122) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4093), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n121) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4094), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n120) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4095), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n119) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4096), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n118) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4097), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n117) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_54__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4098), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n116) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4115), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n115) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4116), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n114) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4117), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n113) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4118), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n112) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4119), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n111) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4120), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n110) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4121), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n109) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_51__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4122), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n108) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4123), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n107) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4124), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n106) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4125), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n105) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4126), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n104) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4127), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n103) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4128), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n102) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4129), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n101) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_50__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4130), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n100) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2691), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n483) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2692), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n482) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2693), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n481) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2694), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n480) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2695), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n479) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2696), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n478) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2697), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n477) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_229__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2698), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n476) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2723), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n467) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2724), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n466) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2725), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n465) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2726), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n464) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2727), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n463) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2728), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n462) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2729), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n461) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_225__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2730), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n460) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2867), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n451) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2868), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n450) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2869), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n449) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2870), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n448) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2871), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n447) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2872), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n446) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2873), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n445) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_207__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2874), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n444) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2915), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n435) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2916), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n434) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2917), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n433) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2918), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n432) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2919), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n431) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2920), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n430) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2921), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n429) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_201__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2922), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n428) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2947), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n419) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2948), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n418) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2949), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n417) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2950), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n416) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2951), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n415) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2952), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n414) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2953), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n413) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_197__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2954), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n412) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2979), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n403) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2980), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n402) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2981), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n401) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2982), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n400) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2983), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n399) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2984), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n398) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2985), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n397) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_193__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2986), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n396) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3203), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n355) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3204), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n354) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3205), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n353) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3206), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n352) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3207), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n351) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3208), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n350) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3209), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n349) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_165__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3210), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n348) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3235), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n339) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3236), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n338) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3237), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n337) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3238), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n336) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3239), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n335) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3240), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n334) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3241), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n333) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_161__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3242), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n332) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3379), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n323) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3380), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n322) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3381), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n321) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3382), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n320) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3383), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n319) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3384), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n318) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3385), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n317) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_143__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3386), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n316) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3427), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n307) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3428), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n306) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3429), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n305) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3430), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n304) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3431), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n303) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3432), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n302) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3433), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n301) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_137__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3434), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n300) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3459), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n291) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3460), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n290) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3461), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n289) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3462), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n288) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3463), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n287) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3464), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n286) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3465), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n285) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_133__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3466), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n284) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3491), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n275) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3492), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n274) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3493), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n273) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3494), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n272) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3495), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n271) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3496), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n270) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3497), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n269) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_129__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3498), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n268) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3715), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n227) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3716), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n226) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3717), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n225) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3718), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n224) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3719), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n223) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3720), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n222) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3721), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n221) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_101__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3722), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n220) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3747), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n211) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3748), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n210) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3749), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n209) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3750), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n208) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3751), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n207) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3752), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n206) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3753), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n205) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_97__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3754), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n204) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3891), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n195) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3892), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n194) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3893), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n193) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3894), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n192) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3895), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n191) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3896), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n190) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3897), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n189) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_79__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3898), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n188) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3939), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n179) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3940), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n178) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3941), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n177) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3942), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n176) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3943), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n175) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3944), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n174) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3945), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n173) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_73__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3946), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n172) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3971), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n163) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3972), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n162) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3973), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n161) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3974), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n160) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3975), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n159) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3976), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n158) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3977), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n157) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_69__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3978), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n156) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4003), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n147) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4004), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n146) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4005), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n145) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4006), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n144) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4007), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n143) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4008), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n142) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4009), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n141) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_65__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4010), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n140) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4227), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n99) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4228), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n98) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4229), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n97) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4230), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n96) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4231), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n95) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4232), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n94) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4233), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n93) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_37__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4234), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n92) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4259), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n83) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4260), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n82) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4261), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n81) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4262), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n80) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4263), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n79) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4264), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n78) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4265), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n77) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_33__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4266), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n76) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4403), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n67) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4404), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n66) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4405), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n65) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4406), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n64) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4407), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n63) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4408), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n62) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4409), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n61) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_15__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4410), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n60) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4451), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n51) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4452), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n50) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4453), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n49) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4454), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n48) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4455), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n47) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4456), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n46) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4457), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n45) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_9__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4458), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n44) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4483), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n35) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4484), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n34) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4485), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n33) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4486), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n32) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4487), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n31) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4488), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n30) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4489), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n29) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_5__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4490), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n28) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4515), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n19) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4516), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n18) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4517), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n17) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4518), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n16) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4519), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n15) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4520), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n14) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4521), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n13) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_1__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4522), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n12) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2699), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n475) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2700), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n474) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2701), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n473) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2702), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n472) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2703), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n471) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2704), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n470) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2705), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n469) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_228__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2706), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n468) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2731), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n459) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2732), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n458) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2733), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n457) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2734), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n456) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2735), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n455) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2736), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n454) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2737), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n453) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_224__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2738), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n452) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2875), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n443) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2876), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n442) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2877), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n441) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2878), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n440) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2879), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n439) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2880), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n438) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2881), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n437) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_206__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2882), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n436) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2923), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n427) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2924), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n426) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2925), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n425) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2926), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n424) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2927), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n423) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2928), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n422) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2929), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n421) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_200__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2930), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n420) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2955), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n411) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2956), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n410) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2957), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n409) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2958), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n408) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2959), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n407) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2960), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n406) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2961), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n405) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_196__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2962), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n404) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2987), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n395) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2988), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n394) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2989), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n393) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2990), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n392) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2991), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n391) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2992), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n390) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2993), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n389) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_192__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2994), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n388) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3211), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n347) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3212), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n346) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3213), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n345) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3214), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n344) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3215), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n343) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3216), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n342) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3217), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n341) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_164__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3218), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n340) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3243), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n331) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3244), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n330) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3245), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n329) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3246), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n328) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3247), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n327) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3248), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n326) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3249), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n325) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_160__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3250), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n324) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3387), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n315) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3388), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n314) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3389), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n313) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3390), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n312) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3391), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n311) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3392), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n310) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3393), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n309) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_142__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3394), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n308) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3435), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n299) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3436), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n298) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3437), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n297) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3438), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n296) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3439), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n295) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3440), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n294) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3441), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n293) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_136__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3442), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n292) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3467), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n283) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3468), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n282) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3469), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n281) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3470), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n280) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3471), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n279) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3472), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n278) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3473), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n277) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_132__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3474), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n276) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3499), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n267) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3500), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n266) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3501), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n265) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3502), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n264) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3503), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n263) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3504), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n262) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3505), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n261) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_128__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3506), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n260) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3723), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n219) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3724), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n218) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3725), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n217) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3726), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n216) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3727), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n215) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3728), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n214) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3729), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n213) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_100__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3730), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n212) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3755), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n203) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3756), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n202) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3757), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n201) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3758), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n200) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3759), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n199) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3760), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n198) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3761), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n197) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_96__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3762), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n196) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3899), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n187) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3900), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n186) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3901), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n185) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3902), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n184) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3903), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n183) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3904), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n182) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3905), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n181) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_78__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3906), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n180) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3947), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n171) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3948), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n170) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3949), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n169) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3950), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n168) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3951), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n167) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3952), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n166) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3953), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n165) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_72__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3954), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n164) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3979), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n155) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3980), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n154) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3981), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n153) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3982), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n152) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3983), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n151) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3984), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n150) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3985), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n149) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_68__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3986), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n148) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4011), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n139) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4012), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n138) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4013), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n137) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4014), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n136) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4015), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n135) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4016), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n134) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4017), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n133) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_64__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4018), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n132) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4235), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n91) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4236), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n90) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4237), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n89) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4238), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n88) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4239), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n87) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4240), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n86) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4241), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n85) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_36__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4242), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n84) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4267), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n75) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4268), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n74) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4269), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n73) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4270), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n72) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4271), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n71) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4272), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n70) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4273), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n69) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_32__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4274), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n68) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4411), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n59) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4412), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n58) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4413), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n57) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4414), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n56) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4415), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n55) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4416), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n54) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4417), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n53) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_14__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4418), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n52) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4459), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n43) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4460), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n42) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4461), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n41) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4462), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n40) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4463), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n39) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4464), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n38) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4465), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n37) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_8__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4466), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n36) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4491), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n27) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4492), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n26) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4493), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n25) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4494), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n24) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4495), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n23) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4496), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n22) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4497), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n21) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_4__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4498), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n20) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4523), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n11) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4524), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n10) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4525), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n9) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4526), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n8) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4527), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n7) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4528), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n6) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4529), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n5) );
  DFFQN_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_0__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4530), .CK(wb_clk_i), .QN(
        oc8051_ram_top1_oc8051_idata_n4) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2475), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[0]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2476), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[1]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2477), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[2]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2478), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[3]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2479), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[4]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2480), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[5]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2481), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[6]) );
  DFFRPQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_rd_data_reg_7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2482), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_ram_top1_rd_data_m[7]) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2675), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2676), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2677), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2678), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2679), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2680), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2681), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_231__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2682), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_231__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2707), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2708), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2709), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2710), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2711), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2712), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2713), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_227__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2714), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_227__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2883), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2884), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2885), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2886), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2887), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2888), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2889), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_205__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2890), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_205__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2899), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2900), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2901), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2902), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2903), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2904), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2905), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_203__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2906), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_203__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2931), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2932), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2933), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2934), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2935), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2936), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2937), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_199__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2938), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_199__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2963), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2964), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2965), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2966), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2967), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2968), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2969), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_195__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2970), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_195__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3187), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3188), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3189), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3190), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3191), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3192), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3193), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_167__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3194), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_167__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3219), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3220), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3221), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3222), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3223), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3224), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3225), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_163__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3226), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_163__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3395), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3396), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3397), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3398), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3399), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3400), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3401), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_141__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3402), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_141__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3411), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3412), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3413), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3414), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3415), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3416), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3417), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_139__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3418), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_139__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3443), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3444), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3445), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3446), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3447), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3448), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3449), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_135__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3450), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_135__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3475), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3476), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3477), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3478), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3479), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3480), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3481), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_131__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3482), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_131__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3699), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3700), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3701), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3702), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3703), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3704), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3705), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_103__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3706), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_103__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3731), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3732), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3733), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3734), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3735), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3736), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3737), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_99__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3738), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_99__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3907), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3908), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3909), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3910), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3911), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3912), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3913), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_77__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3914), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_77__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3923), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3924), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3925), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3926), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3927), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3928), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3929), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_75__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3930), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_75__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3955), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3956), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3957), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3958), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3959), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3960), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3961), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_71__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3962), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_71__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3987), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3988), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3989), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3990), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3991), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3992), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3993), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_67__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3994), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_67__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4211), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4212), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4213), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4214), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4215), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4216), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4217), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_39__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4218), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_39__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4243), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4244), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4245), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4246), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4247), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4248), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4249), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_35__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4250), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_35__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4419), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4420), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4421), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4422), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4423), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4424), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4425), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_13__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4426), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_13__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4435), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4436), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4437), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4438), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4439), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4440), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4441), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_11__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4442), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_11__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4467), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4468), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4469), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4470), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4471), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4472), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4473), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_7__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4474), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_7__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4499), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4500), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4501), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4502), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4503), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4504), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4505), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_3__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4506), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_3__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2491), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2492), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2493), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2494), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2495), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2496), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2497), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_254__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2498), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_254__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2507), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2508), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2509), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2510), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2511), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2512), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2513), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_252__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2514), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_252__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2515), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2516), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2517), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2518), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2519), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2520), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2521), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_251__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2522), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_251__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2523), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2524), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2525), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2526), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2527), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2528), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2529), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_250__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2530), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_250__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2531), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2532), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2533), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2534), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2535), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2536), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2537), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_249__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2538), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_249__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2539), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2540), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2541), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2542), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2543), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2544), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2545), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_248__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2546), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_248__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2643), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2644), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2645), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2646), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2647), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2648), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2649), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_235__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2650), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_235__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2659), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2660), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2661), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2662), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2663), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2664), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2665), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_233__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2666), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_233__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2747), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2748), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2749), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2750), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2751), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2752), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2753), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_222__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2754), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_222__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2763), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2764), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2765), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2766), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2767), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2768), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2769), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_220__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2770), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_220__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2779), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2780), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2781), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2782), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2783), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2784), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2785), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_218__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2786), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_218__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2795), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2796), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2797), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2798), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2799), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2800), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2801), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_216__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2802), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_216__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2811), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2812), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2813), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2814), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2815), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2816), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2817), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_214__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2818), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_214__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2827), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2828), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2829), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2830), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2831), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2832), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2833), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_212__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2834), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_212__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2843), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2844), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2845), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2846), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2847), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2848), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2849), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_210__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2850), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_210__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2859), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2860), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2861), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2862), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2863), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2864), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2865), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_208__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2866), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_208__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3003), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3004), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3005), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3006), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3007), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3008), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3009), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_190__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3010), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_190__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3019), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3020), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3021), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3022), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3023), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3024), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3025), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_188__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3026), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_188__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3027), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3028), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3029), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3030), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3031), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3032), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3033), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_187__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3034), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_187__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3035), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3036), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3037), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3038), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3039), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3040), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3041), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_186__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3042), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_186__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3043), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3044), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3045), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3046), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3047), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3048), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3049), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_185__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3050), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_185__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3051), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3052), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3053), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3054), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3055), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3056), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3057), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_184__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3058), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_184__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3155), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3156), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3157), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3158), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3159), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3160), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3161), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_171__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3162), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_171__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3171), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3172), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3173), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3174), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3175), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3176), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3177), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_169__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3178), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_169__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3259), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3260), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3261), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3262), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3263), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3264), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3265), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_158__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3266), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_158__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3275), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3276), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3277), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3278), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3279), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3280), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3281), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_156__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3282), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_156__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3291), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3292), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3293), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3294), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3295), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3296), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3297), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_154__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3298), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_154__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3307), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3308), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3309), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3310), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3311), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3312), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3313), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_152__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3314), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_152__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3323), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3324), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3325), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3326), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3327), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3328), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3329), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_150__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3330), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_150__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3339), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3340), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3341), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3342), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3343), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3344), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3345), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_148__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3346), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_148__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3355), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3356), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3357), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3358), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3359), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3360), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3361), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_146__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3362), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_146__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3371), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3372), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3373), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3374), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3375), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3376), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3377), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_144__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3378), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_144__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3515), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3516), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3517), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3518), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3519), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3520), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3521), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_126__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3522), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_126__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3531), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3532), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3533), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3534), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3535), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3536), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3537), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_124__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3538), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_124__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3539), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3540), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3541), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3542), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3543), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3544), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3545), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_123__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3546), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_123__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3547), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3548), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3549), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3550), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3551), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3552), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3553), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_122__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3554), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_122__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3555), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3556), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3557), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3558), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3559), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3560), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3561), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_121__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3562), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_121__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3563), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3564), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3565), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3566), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3567), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3568), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3569), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_120__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3570), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_120__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3667), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3668), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3669), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3670), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3671), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3672), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3673), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_107__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3674), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_107__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3683), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3684), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3685), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3686), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3687), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3688), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3689), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_105__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3690), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_105__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3771), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3772), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3773), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3774), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3775), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3776), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3777), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_94__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3778), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_94__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3787), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3788), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3789), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3790), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3791), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3792), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3793), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_92__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3794), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_92__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3803), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3804), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3805), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3806), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3807), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3808), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3809), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_90__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3810), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_90__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3819), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3820), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3821), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3822), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3823), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3824), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3825), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_88__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3826), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_88__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3835), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3836), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3837), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3838), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3839), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3840), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3841), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_86__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3842), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_86__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3851), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3852), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3853), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3854), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3855), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3856), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3857), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_84__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3858), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_84__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3867), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3868), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3869), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3870), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3871), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3872), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3873), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_82__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3874), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_82__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3883), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3884), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3885), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3886), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3887), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3888), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3889), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_80__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3890), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_80__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4027), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4028), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4029), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4030), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4031), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4032), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4033), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_62__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4034), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_62__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4043), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4044), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4045), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4046), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4047), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4048), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4049), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_60__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4050), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_60__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4051), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4052), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4053), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4054), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4055), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4056), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4057), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_59__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4058), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_59__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4059), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4060), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4061), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4062), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4063), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4064), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4065), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_58__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4066), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_58__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4067), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4068), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4069), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4070), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4071), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4072), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4073), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_57__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4074), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_57__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4075), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4076), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4077), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4078), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4079), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4080), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4081), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_56__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4082), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_56__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4179), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4180), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4181), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4182), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4183), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4184), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4185), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_43__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4186), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_43__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4195), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4196), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4197), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4198), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4199), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4200), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4201), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_41__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4202), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_41__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4283), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4284), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4285), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4286), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4287), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4288), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4289), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_30__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4290), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_30__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4299), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4300), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4301), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4302), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4303), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4304), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4305), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_28__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4306), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_28__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4315), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4316), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4317), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4318), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4319), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4320), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4321), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_26__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4322), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_26__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4331), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4332), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4333), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4334), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4335), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4336), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4337), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_24__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4338), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_24__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4347), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4348), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4349), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4350), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4351), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4352), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4353), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_22__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4354), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_22__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4363), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4364), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4365), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4366), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4367), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4368), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4369), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_20__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4370), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_20__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4379), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4380), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4381), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4382), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4383), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4384), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4385), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_18__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4386), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_18__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4395), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4396), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4397), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4398), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4399), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4400), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4401), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_16__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4402), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_16__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2683), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2684), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2685), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2686), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2687), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2688), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2689), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_230__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2690), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_230__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2715), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2716), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2717), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2718), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2719), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2720), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2721), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_226__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2722), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_226__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2891), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2892), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2893), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2894), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2895), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2896), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2897), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_204__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2898), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_204__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2907), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2908), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2909), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2910), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2911), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2912), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2913), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_202__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2914), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_202__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2939), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2940), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2941), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2942), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2943), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2944), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2945), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_198__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2946), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_198__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2971), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2972), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2973), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2974), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2975), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2976), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2977), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_194__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2978), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_194__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3195), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3196), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3197), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3198), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3199), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3200), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3201), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_166__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3202), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_166__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3227), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3228), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3229), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3230), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3231), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3232), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3233), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_162__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3234), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_162__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3403), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3404), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3405), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3406), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3407), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3408), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3409), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_140__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3410), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_140__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3419), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3420), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3421), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3422), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3423), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3424), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3425), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_138__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3426), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_138__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3451), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3452), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3453), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3454), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3455), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3456), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3457), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_134__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3458), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_134__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3483), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3484), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3485), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3486), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3487), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3488), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3489), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_130__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3490), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_130__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3707), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3708), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3709), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3710), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3711), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3712), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3713), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_102__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3714), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_102__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3739), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3740), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3741), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3742), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3743), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3744), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3745), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_98__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3746), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_98__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3915), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3916), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3917), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3918), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3919), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3920), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3921), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_76__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3922), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_76__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3931), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3932), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3933), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3934), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3935), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3936), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3937), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_74__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3938), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_74__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3963), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3964), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3965), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3966), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3967), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3968), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3969), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_70__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3970), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_70__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3995), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3996), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3997), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3998), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3999), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4000), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4001), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_66__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4002), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_66__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4219), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4220), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4221), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4222), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4223), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4224), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4225), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_38__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4226), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_38__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4251), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4252), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4253), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4254), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4255), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4256), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4257), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_34__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4258), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_34__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4427), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4428), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4429), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4430), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4431), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4432), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4433), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_12__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4434), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_12__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4443), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4444), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4445), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4446), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4447), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4448), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4449), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_10__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4450), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_10__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4475), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4476), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4477), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4478), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4479), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4480), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4481), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_6__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4482), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_6__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4507), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4508), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4509), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4510), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4511), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4512), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4513), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_2__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4514), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_2__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2483), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2484), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2485), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2486), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2487), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2488), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2489), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_255__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2490), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_255__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2499), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2500), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2501), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2502), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2503), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2504), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2505), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_253__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2506), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_253__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2611), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2612), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2613), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2614), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2615), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2616), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2617), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_239__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2618), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_239__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2619), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2620), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2621), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2622), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2623), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2624), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2625), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_238__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2626), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_238__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2627), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2628), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2629), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2630), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2631), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2632), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2633), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_237__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2634), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_237__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2635), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2636), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2637), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2638), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2639), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2640), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2641), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_236__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2642), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_236__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2651), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2652), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2653), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2654), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2655), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2656), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2657), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_234__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2658), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_234__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2667), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2668), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2669), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2670), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2671), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2672), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2673), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_232__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2674), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_232__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2739), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2740), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2741), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2742), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2743), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2744), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2745), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_223__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2746), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_223__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2755), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2756), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2757), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2758), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2759), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2760), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2761), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_221__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2762), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_221__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2771), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2772), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2773), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2774), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2775), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2776), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2777), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_219__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2778), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_219__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2787), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2788), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2789), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2790), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2791), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2792), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2793), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_217__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2794), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_217__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2803), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2804), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2805), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2806), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2807), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2808), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2809), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_215__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2810), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_215__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2819), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2820), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2821), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2822), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2823), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2824), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2825), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_213__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2826), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_213__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2835), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2836), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2837), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2838), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2839), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2840), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2841), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_211__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2842), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_211__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2851), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2852), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2853), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2854), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2855), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2856), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2857), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_209__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2858), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_209__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2995), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2996), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2997), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2998), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2999), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3000), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3001), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_191__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3002), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_191__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3011), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3012), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3013), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3014), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3015), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3016), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3017), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_189__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3018), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_189__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3123), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3124), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3125), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3126), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3127), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3128), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3129), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_175__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3130), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_175__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3131), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3132), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3133), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3134), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3135), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3136), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3137), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_174__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3138), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_174__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3139), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3140), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3141), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3142), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3143), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3144), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3145), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_173__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3146), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_173__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3147), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3148), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3149), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3150), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3151), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3152), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3153), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_172__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3154), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_172__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3163), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3164), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3165), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3166), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3167), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3168), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3169), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_170__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3170), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_170__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3179), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3180), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3181), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3182), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3183), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3184), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3185), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_168__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3186), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_168__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3251), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3252), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3253), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3254), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3255), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3256), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3257), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_159__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3258), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_159__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3267), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3268), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3269), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3270), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3271), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3272), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3273), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_157__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3274), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_157__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3283), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3284), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3285), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3286), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3287), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3288), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3289), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_155__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3290), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_155__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3299), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3300), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3301), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3302), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3303), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3304), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3305), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_153__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3306), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_153__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3315), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3316), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3317), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3318), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3319), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3320), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3321), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_151__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3322), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_151__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3331), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3332), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3333), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3334), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3335), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3336), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3337), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_149__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3338), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_149__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3347), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3348), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3349), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3350), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3351), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3352), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3353), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_147__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3354), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_147__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3363), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3364), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3365), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3366), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3367), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3368), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3369), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_145__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3370), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_145__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3507), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3508), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3509), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3510), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3511), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3512), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3513), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_127__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3514), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_127__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3523), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3524), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3525), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3526), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3527), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3528), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3529), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_125__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3530), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_125__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3635), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3636), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3637), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3638), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3639), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3640), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3641), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_111__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3642), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_111__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3643), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3644), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3645), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3646), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3647), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3648), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3649), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_110__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3650), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_110__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3651), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3652), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3653), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3654), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3655), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3656), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3657), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_109__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3658), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_109__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3659), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3660), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3661), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3662), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3663), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3664), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3665), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_108__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3666), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_108__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3675), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3676), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3677), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3678), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3679), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3680), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3681), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_106__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3682), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_106__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3691), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3692), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3693), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3694), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3695), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3696), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3697), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_104__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3698), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_104__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3763), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3764), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3765), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3766), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3767), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3768), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3769), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_95__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3770), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_95__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3779), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3780), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3781), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3782), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3783), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3784), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3785), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_93__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3786), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_93__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3795), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3796), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3797), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3798), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3799), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3800), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3801), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_91__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3802), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_91__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3811), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3812), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3813), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3814), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3815), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3816), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3817), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_89__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3818), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_89__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3827), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3828), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3829), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3830), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3831), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3832), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3833), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_87__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3834), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_87__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3843), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3844), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3845), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3846), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3847), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3848), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3849), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_85__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3850), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_85__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3859), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3860), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3861), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3862), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3863), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3864), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3865), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_83__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3866), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_83__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3875), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3876), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3877), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3878), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3879), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3880), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3881), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_81__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3882), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_81__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4019), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4020), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4021), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4022), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4023), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4024), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4025), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_63__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4026), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_63__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4035), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4036), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4037), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4038), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4039), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4040), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4041), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_61__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4042), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_61__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4147), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4148), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4149), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4150), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4151), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4152), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4153), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_47__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4154), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_47__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4155), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4156), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4157), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4158), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4159), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4160), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4161), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_46__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4162), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_46__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4163), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4164), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4165), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4166), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4167), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4168), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4169), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_45__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4170), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_45__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4171), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4172), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4173), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4174), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4175), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4176), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4177), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_44__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4178), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_44__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4187), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4188), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4189), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4190), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4191), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4192), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4193), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_42__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4194), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_42__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4203), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4204), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4205), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4206), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4207), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4208), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4209), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_40__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4210), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_40__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4275), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4276), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4277), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4278), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4279), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4280), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4281), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_31__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4282), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_31__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4291), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4292), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4293), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4294), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4295), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4296), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4297), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_29__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4298), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_29__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4307), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4308), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4309), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4310), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4311), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4312), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4313), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_27__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4314), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_27__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4323), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4324), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4325), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4326), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4327), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4328), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4329), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_25__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4330), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_25__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4339), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4340), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4341), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4342), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4343), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4344), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4345), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_23__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4346), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_23__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4355), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4356), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4357), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4358), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4359), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4360), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4361), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_21__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4362), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_21__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4371), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4372), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4373), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4374), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4375), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4376), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4377), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_19__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4378), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_19__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4387), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4388), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4389), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4390), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4391), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4392), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4393), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_17__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4394), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_17__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2563), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2564), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2565), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2566), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2567), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2568), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2569), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_245__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2570), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_245__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2571), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2572), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2573), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2574), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2575), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2576), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2577), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_244__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2578), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_244__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2595), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2596), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2597), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2598), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2599), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2600), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2601), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_241__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2602), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_241__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2603), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2604), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2605), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2606), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2607), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2608), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2609), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_240__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n2610), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_240__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3075), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3076), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3077), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3078), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3079), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3080), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3081), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_181__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3082), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_181__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3083), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3084), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3085), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3086), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3087), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3088), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3089), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_180__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3090), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_180__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3107), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3108), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3109), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3110), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3111), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3112), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3113), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_177__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3114), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_177__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3115), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3116), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3117), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3118), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3119), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3120), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3121), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_176__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3122), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_176__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3587), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3588), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3589), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3590), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3591), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3592), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3593), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_117__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3594), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_117__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3595), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3596), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3597), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3598), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3599), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3600), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3601), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_116__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3602), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_116__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3619), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3620), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3621), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3622), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3623), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3624), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3625), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_113__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3626), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_113__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3627), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3628), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3629), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3630), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3631), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3632), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3633), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_112__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n3634), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_112__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4099), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4100), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4101), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4102), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4103), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4104), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4105), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_53__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4106), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_53__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4107), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4108), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4109), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4110), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4111), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4112), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4113), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_52__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4114), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_52__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4131), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4132), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4133), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4134), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4135), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4136), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4137), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_49__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4138), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_49__7_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__0_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4139), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__0_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__1_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4140), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__1_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__2_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4141), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__2_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__3_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4142), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__3_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__4_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4143), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__4_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__5_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4144), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__5_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__6_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4145), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__6_) );
  DFFQ_X1M_A12TS oc8051_ram_top1_oc8051_idata_buff_reg_48__7_ ( .D(
        oc8051_ram_top1_oc8051_idata_n4146), .CK(wb_clk_i), .Q(
        oc8051_ram_top1_oc8051_idata_buff_48__7_) );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u87 ( .A(src_sel1[1]), .B(src_sel1[2]), 
        .C(src_sel1[0]), .Y(oc8051_alu_src_sel1_n36) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u86 ( .A(src_sel1[2]), .Y(
        oc8051_alu_src_sel1_n60) );
  NOR2_X0P5A_A12TS oc8051_alu_src_sel1_u85 ( .A(oc8051_alu_src_sel1_n60), .B(
        src_sel1[0]), .Y(oc8051_alu_src_sel1_n37) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u84 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[0]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[8]), .Y(
        oc8051_alu_src_sel1_n56) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u83 ( .A(src_sel1[0]), .Y(
        oc8051_alu_src_sel1_n59) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u82 ( .A(src_sel1[1]), .Y(
        oc8051_alu_src_sel1_n61) );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u81 ( .A(oc8051_alu_src_sel1_n59), .B(
        src_sel1[2]), .C(oc8051_alu_src_sel1_n61), .Y(oc8051_alu_src_sel1_n34)
         );
  NOR2_X0P5A_A12TS oc8051_alu_src_sel1_u80 ( .A(oc8051_alu_src_sel1_n60), .B(
        oc8051_alu_src_sel1_n61), .Y(oc8051_alu_src_sel1_n35) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u79 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[0]), .B0(oc8051_alu_src_sel1_op1_r[0]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n57) );
  NOR2_X0P5A_A12TS oc8051_alu_src_sel1_u78 ( .A(oc8051_alu_src_sel1_n61), .B(
        src_sel1[0]), .Y(oc8051_alu_src_sel1_n31) );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u77 ( .A(oc8051_alu_src_sel1_n59), .B(
        src_sel1[1]), .C(oc8051_alu_src_sel1_n60), .Y(oc8051_alu_src_sel1_n32)
         );
  NOR3_X0P5A_A12TS oc8051_alu_src_sel1_u76 ( .A(src_sel1[1]), .B(src_sel1[2]), 
        .C(oc8051_alu_src_sel1_n59), .Y(oc8051_alu_src_sel1_n33) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u75 ( .A0(
        oc8051_alu_src_sel1_op3_r[0]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[0]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_0_), .Y(oc8051_alu_src_sel1_n58) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u74 ( .A(oc8051_alu_src_sel1_n56), .B(
        oc8051_alu_src_sel1_n57), .C(oc8051_alu_src_sel1_n58), .Y(src1[0]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u73 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[1]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[9]), .Y(
        oc8051_alu_src_sel1_n53) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u72 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[1]), .B0(oc8051_alu_src_sel1_op1_r[1]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n54) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u71 ( .A0(
        oc8051_alu_src_sel1_op3_r[1]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[1]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_1_), .Y(oc8051_alu_src_sel1_n55) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u70 ( .A(oc8051_alu_src_sel1_n53), .B(
        oc8051_alu_src_sel1_n54), .C(oc8051_alu_src_sel1_n55), .Y(src1[1]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u69 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[2]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[10]), .Y(
        oc8051_alu_src_sel1_n50) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u68 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[2]), .B0(oc8051_alu_src_sel1_op1_r[2]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n51) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u67 ( .A0(
        oc8051_alu_src_sel1_op3_r[2]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[2]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_2_), .Y(oc8051_alu_src_sel1_n52) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u66 ( .A(oc8051_alu_src_sel1_n50), .B(
        oc8051_alu_src_sel1_n51), .C(oc8051_alu_src_sel1_n52), .Y(src1[2]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u65 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[3]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[11]), .Y(
        oc8051_alu_src_sel1_n47) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u64 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[3]), .B0(oc8051_alu_src_sel1_op1_r[3]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n48) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u63 ( .A0(
        oc8051_alu_src_sel1_op3_r[3]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[3]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_3_), .Y(oc8051_alu_src_sel1_n49) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u62 ( .A(oc8051_alu_src_sel1_n47), .B(
        oc8051_alu_src_sel1_n48), .C(oc8051_alu_src_sel1_n49), .Y(src1[3]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u61 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[4]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[12]), .Y(
        oc8051_alu_src_sel1_n44) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u60 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[4]), .B0(oc8051_alu_src_sel1_op1_r[4]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n45) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u59 ( .A0(
        oc8051_alu_src_sel1_op3_r[4]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[4]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_4_), .Y(oc8051_alu_src_sel1_n46) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u58 ( .A(oc8051_alu_src_sel1_n44), .B(
        oc8051_alu_src_sel1_n45), .C(oc8051_alu_src_sel1_n46), .Y(src1[4]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u57 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[5]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[13]), .Y(
        oc8051_alu_src_sel1_n41) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u56 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[5]), .B0(oc8051_alu_src_sel1_op1_r[5]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n42) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u55 ( .A0(
        oc8051_alu_src_sel1_op3_r[5]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[5]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_5_), .Y(oc8051_alu_src_sel1_n43) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u54 ( .A(oc8051_alu_src_sel1_n41), .B(
        oc8051_alu_src_sel1_n42), .C(oc8051_alu_src_sel1_n43), .Y(src1[5]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u53 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[6]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[14]), .Y(
        oc8051_alu_src_sel1_n38) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u52 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[6]), .B0(oc8051_alu_src_sel1_op1_r[6]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n39) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u51 ( .A0(
        oc8051_alu_src_sel1_op3_r[6]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[6]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_6_), .Y(oc8051_alu_src_sel1_n40) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u50 ( .A(oc8051_alu_src_sel1_n38), .B(
        oc8051_alu_src_sel1_n39), .C(oc8051_alu_src_sel1_n40), .Y(src1[6]) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u49 ( .A0(oc8051_alu_src_sel1_n36), 
        .A1(ram_out[7]), .B0(oc8051_alu_src_sel1_n37), .B1(pc[15]), .Y(
        oc8051_alu_src_sel1_n28) );
  AOI22_X0P5M_A12TS oc8051_alu_src_sel1_u48 ( .A0(oc8051_alu_src_sel1_n34), 
        .A1(acc[7]), .B0(oc8051_alu_src_sel1_op1_r[7]), .B1(
        oc8051_alu_src_sel1_n35), .Y(oc8051_alu_src_sel1_n29) );
  AOI222_X0P5M_A12TS oc8051_alu_src_sel1_u47 ( .A0(
        oc8051_alu_src_sel1_op3_r[7]), .A1(oc8051_alu_src_sel1_n31), .B0(pc[7]), .B1(oc8051_alu_src_sel1_n32), .C0(oc8051_alu_src_sel1_n33), .C1(
        oc8051_alu_src_sel1_op2_r_7_), .Y(oc8051_alu_src_sel1_n30) );
  NAND3_X0P5A_A12TS oc8051_alu_src_sel1_u46 ( .A(oc8051_alu_src_sel1_n28), .B(
        oc8051_alu_src_sel1_n29), .C(oc8051_alu_src_sel1_n30), .Y(src1[7]) );
  NAND2_X0P5A_A12TS oc8051_alu_src_sel1_u45 ( .A(src_sel2[1]), .B(src_sel2[0]), 
        .Y(oc8051_alu_src_sel1_n1) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u44 ( .A(oc8051_alu_src_sel1_op2_r_0_), 
        .Y(oc8051_alu_src_sel1_n25) );
  NAND2B_X0P5M_A12TS oc8051_alu_src_sel1_u43 ( .AN(src_sel2[1]), .B(
        src_sel2[0]), .Y(oc8051_alu_src_sel1_n3) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u42 ( .A(acc[0]), .Y(
        oc8051_alu_src_sel1_n26) );
  OR2_X0P5M_A12TS oc8051_alu_src_sel1_u41 ( .A(src_sel2[0]), .B(src_sel2[1]), 
        .Y(oc8051_alu_src_sel1_n5) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u40 ( .A(ram_out[0]), .Y(
        oc8051_alu_src_sel1_n27) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u39 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n25), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n26), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n27), .Y(src2[0]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u38 ( .A(oc8051_alu_src_sel1_op2_r_1_), 
        .Y(oc8051_alu_src_sel1_n22) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u37 ( .A(acc[1]), .Y(
        oc8051_alu_src_sel1_n23) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u36 ( .A(ram_out[1]), .Y(
        oc8051_alu_src_sel1_n24) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u35 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n22), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n23), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n24), .Y(src2[1]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u34 ( .A(oc8051_alu_src_sel1_op2_r_2_), 
        .Y(oc8051_alu_src_sel1_n19) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u33 ( .A(acc[2]), .Y(
        oc8051_alu_src_sel1_n20) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u32 ( .A(ram_out[2]), .Y(
        oc8051_alu_src_sel1_n21) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u31 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n19), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n20), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n21), .Y(src2[2]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u30 ( .A(oc8051_alu_src_sel1_op2_r_3_), 
        .Y(oc8051_alu_src_sel1_n16) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u29 ( .A(acc[3]), .Y(
        oc8051_alu_src_sel1_n17) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u28 ( .A(ram_out[3]), .Y(
        oc8051_alu_src_sel1_n18) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u27 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n16), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n17), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n18), .Y(src2[3]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u26 ( .A(oc8051_alu_src_sel1_op2_r_4_), 
        .Y(oc8051_alu_src_sel1_n13) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u25 ( .A(acc[4]), .Y(
        oc8051_alu_src_sel1_n14) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u24 ( .A(ram_out[4]), .Y(
        oc8051_alu_src_sel1_n15) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u23 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n13), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n14), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n15), .Y(src2[4]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u22 ( .A(oc8051_alu_src_sel1_op2_r_5_), 
        .Y(oc8051_alu_src_sel1_n10) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u21 ( .A(acc[5]), .Y(
        oc8051_alu_src_sel1_n11) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u20 ( .A(ram_out[5]), .Y(
        oc8051_alu_src_sel1_n12) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u19 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n10), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n11), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n12), .Y(src2[5]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u18 ( .A(oc8051_alu_src_sel1_op2_r_6_), 
        .Y(oc8051_alu_src_sel1_n7) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u17 ( .A(acc[6]), .Y(
        oc8051_alu_src_sel1_n8) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u16 ( .A(ram_out[6]), .Y(
        oc8051_alu_src_sel1_n9) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u15 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n7), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n8), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n9), .Y(src2[6]) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u14 ( .A(oc8051_alu_src_sel1_op2_r_7_), 
        .Y(oc8051_alu_src_sel1_n2) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u13 ( .A(acc[7]), .Y(
        oc8051_alu_src_sel1_n4) );
  INV_X0P5B_A12TS oc8051_alu_src_sel1_u12 ( .A(ram_out[7]), .Y(
        oc8051_alu_src_sel1_n6) );
  OAI222_X0P5M_A12TS oc8051_alu_src_sel1_u11 ( .A0(oc8051_alu_src_sel1_n1), 
        .A1(oc8051_alu_src_sel1_n2), .B0(oc8051_alu_src_sel1_n3), .B1(
        oc8051_alu_src_sel1_n4), .C0(oc8051_alu_src_sel1_n5), .C1(
        oc8051_alu_src_sel1_n6), .Y(src2[7]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u10 ( .A(dptr_hi[0]), .B(pc[8]), .S0(
        src_sel3), .Y(src3[0]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u9 ( .A(dptr_hi[1]), .B(pc[9]), .S0(
        src_sel3), .Y(src3[1]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u8 ( .A(dptr_hi[2]), .B(pc[10]), .S0(
        src_sel3), .Y(src3[2]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u7 ( .A(dptr_hi[3]), .B(pc[11]), .S0(
        src_sel3), .Y(src3[3]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u6 ( .A(dptr_hi[4]), .B(pc[12]), .S0(
        src_sel3), .Y(src3[4]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u5 ( .A(dptr_hi[5]), .B(pc[13]), .S0(
        src_sel3), .Y(src3[5]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u4 ( .A(dptr_hi[6]), .B(pc[14]), .S0(
        src_sel3), .Y(src3[6]) );
  MXT2_X0P5M_A12TS oc8051_alu_src_sel1_u3 ( .A(dptr_hi[7]), .B(pc[15]), .S0(
        src_sel3), .Y(src3[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_0_ ( .D(op2_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_0_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_1_ ( .D(op2_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_1_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_2_ ( .D(op2_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_2_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_3_ ( .D(op2_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_3_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_4_ ( .D(op2_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_4_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_5_ ( .D(op2_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_5_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_6_ ( .D(op2_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_6_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op2_r_reg_7_ ( .D(op2_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op2_r_7_) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_0_ ( .D(op1_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_1_ ( .D(op1_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_2_ ( .D(op1_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_3_ ( .D(op1_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_4_ ( .D(op1_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_5_ ( .D(op1_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_6_ ( .D(op1_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op1_r_reg_7_ ( .D(op1_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op1_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_0_ ( .D(op3_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_1_ ( .D(op3_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_2_ ( .D(op3_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_3_ ( .D(op3_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_4_ ( .D(op3_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_5_ ( .D(op3_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_6_ ( .D(op3_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_alu_src_sel1_op3_r_reg_7_ ( .D(op3_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_alu_src_sel1_op3_r[7]) );
  NOR2_X0P5A_A12TS oc8051_comp1_u11 ( .A(acc[1]), .B(acc[0]), .Y(
        oc8051_comp1_n7) );
  NOR2_X0P5A_A12TS oc8051_comp1_u10 ( .A(acc[3]), .B(acc[2]), .Y(
        oc8051_comp1_n8) );
  NOR2_X0P5A_A12TS oc8051_comp1_u9 ( .A(acc[5]), .B(acc[4]), .Y(
        oc8051_comp1_n9) );
  NOR2_X0P5A_A12TS oc8051_comp1_u8 ( .A(acc[7]), .B(acc[6]), .Y(
        oc8051_comp1_n10) );
  AND4_X0P5M_A12TS oc8051_comp1_u7 ( .A(oc8051_comp1_n7), .B(oc8051_comp1_n8), 
        .C(oc8051_comp1_n9), .D(oc8051_comp1_n10), .Y(oc8051_comp1_n1) );
  NOR2_X0P5A_A12TS oc8051_comp1_u6 ( .A(sub_result[1]), .B(sub_result[0]), .Y(
        oc8051_comp1_n3) );
  NOR2_X0P5A_A12TS oc8051_comp1_u5 ( .A(sub_result[3]), .B(sub_result[2]), .Y(
        oc8051_comp1_n4) );
  NOR2_X0P5A_A12TS oc8051_comp1_u4 ( .A(sub_result[5]), .B(sub_result[4]), .Y(
        oc8051_comp1_n5) );
  NOR2_X0P5A_A12TS oc8051_comp1_u3 ( .A(sub_result[7]), .B(sub_result[6]), .Y(
        oc8051_comp1_n6) );
  AND4_X0P5M_A12TS oc8051_comp1_u2 ( .A(oc8051_comp1_n3), .B(oc8051_comp1_n4), 
        .C(oc8051_comp1_n5), .D(oc8051_comp1_n6), .Y(oc8051_comp1_n2) );
  MXT4_X0P5M_A12TS oc8051_comp1_u1 ( .A(oc8051_comp1_n1), .B(cy), .C(
        oc8051_comp1_n2), .D(bit_out), .S0(comp_sel[1]), .S1(comp_sel[0]), .Y(
        eq) );
  TIEHI_X1M_A12TS oc8051_rom1_u4 ( .Y(oc8051_rom1_ea_int) );
  TIELO_X1M_A12TS oc8051_rom1_u3 ( .Y(oc8051_rom1_data_o_0_) );
  OAI21_X0P5M_A12TS oc8051_cy_select1_u4 ( .A0(cy_sel[0]), .A1(bit_out), .B0(
        cy_sel[1]), .Y(oc8051_cy_select1_n1) );
  AO1B2_X0P5M_A12TS oc8051_cy_select1_u3 ( .B0(cy_sel[0]), .B1(cy), .A0N(
        oc8051_cy_select1_n1), .Y(alu_cy) );
  INV_X0P5B_A12TS oc8051_indi_addr1_u116 ( .A(wr_addr[0]), .Y(
        oc8051_indi_addr1_n26) );
  INV_X0P5B_A12TS oc8051_indi_addr1_u115 ( .A(wr_addr[3]), .Y(
        oc8051_indi_addr1_n92) );
  NOR2B_X0P5M_A12TS oc8051_indi_addr1_u114 ( .AN(wr_o), .B(
        oc8051_indi_addr1_wr_bit_r), .Y(oc8051_indi_addr1_n22) );
  NOR2B_X0P5M_A12TS oc8051_indi_addr1_u113 ( .AN(oc8051_indi_addr1_n22), .B(
        wr_addr[4]), .Y(oc8051_indi_addr1_n95) );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u112 ( .A(oc8051_indi_addr1_n26), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n95), .Y(
        oc8051_indi_addr1_n98) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u111 ( .A(oc8051_indi_addr1_buff_0__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n28)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u110 ( .A(oc8051_indi_addr1_buff_0__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n29)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u109 ( .A(oc8051_indi_addr1_buff_0__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n30)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u108 ( .A(oc8051_indi_addr1_buff_0__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n31)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u107 ( .A(oc8051_indi_addr1_buff_0__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n32)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u106 ( .A(oc8051_indi_addr1_buff_0__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n33)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u105 ( .A(oc8051_indi_addr1_buff_0__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n34)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u104 ( .A(oc8051_indi_addr1_buff_0__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n98), .Y(oc8051_indi_addr1_n35)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u103 ( .A(wr_addr[0]), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n95), .Y(
        oc8051_indi_addr1_n97) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u102 ( .A(oc8051_indi_addr1_buff_1__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n36)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u101 ( .A(oc8051_indi_addr1_buff_1__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n37)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u100 ( .A(oc8051_indi_addr1_buff_1__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n38)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u99 ( .A(oc8051_indi_addr1_buff_1__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n39)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u98 ( .A(oc8051_indi_addr1_buff_1__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n40)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u97 ( .A(oc8051_indi_addr1_buff_1__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n41)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u96 ( .A(oc8051_indi_addr1_buff_1__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n42)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u95 ( .A(oc8051_indi_addr1_buff_1__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n97), .Y(oc8051_indi_addr1_n43)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u94 ( .A(wr_addr[3]), .B(
        oc8051_indi_addr1_n26), .C(oc8051_indi_addr1_n95), .Y(
        oc8051_indi_addr1_n96) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u93 ( .A(oc8051_indi_addr1_buff_2__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n44)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u92 ( .A(oc8051_indi_addr1_buff_2__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n45)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u91 ( .A(oc8051_indi_addr1_buff_2__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n46)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u90 ( .A(oc8051_indi_addr1_buff_2__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n47)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u89 ( .A(oc8051_indi_addr1_buff_2__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n48)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u88 ( .A(oc8051_indi_addr1_buff_2__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n49)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u87 ( .A(oc8051_indi_addr1_buff_2__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n50)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u86 ( .A(oc8051_indi_addr1_buff_2__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n96), .Y(oc8051_indi_addr1_n51)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u85 ( .A(wr_addr[3]), .B(wr_addr[0]), .C(
        oc8051_indi_addr1_n95), .Y(oc8051_indi_addr1_n94) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u84 ( .A(oc8051_indi_addr1_buff_3__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n52)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u83 ( .A(oc8051_indi_addr1_buff_3__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n53)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u82 ( .A(oc8051_indi_addr1_buff_3__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n54)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u81 ( .A(oc8051_indi_addr1_buff_3__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n55)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u80 ( .A(oc8051_indi_addr1_buff_3__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n56)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u79 ( .A(oc8051_indi_addr1_buff_3__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n57)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u78 ( .A(oc8051_indi_addr1_buff_3__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n58)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u77 ( .A(oc8051_indi_addr1_buff_3__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n94), .Y(oc8051_indi_addr1_n59)
         );
  AND2_X0P5M_A12TS oc8051_indi_addr1_u76 ( .A(oc8051_indi_addr1_n22), .B(
        wr_addr[4]), .Y(oc8051_indi_addr1_n24) );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u75 ( .A(oc8051_indi_addr1_n26), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n24), .Y(
        oc8051_indi_addr1_n93) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u74 ( .A(oc8051_indi_addr1_buff_4__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n60)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u73 ( .A(oc8051_indi_addr1_buff_4__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n61)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u72 ( .A(oc8051_indi_addr1_buff_4__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n62)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u71 ( .A(oc8051_indi_addr1_buff_4__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n63)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u70 ( .A(oc8051_indi_addr1_buff_4__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n64)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u69 ( .A(oc8051_indi_addr1_buff_4__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n65)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u68 ( .A(oc8051_indi_addr1_buff_4__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n66)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u67 ( .A(oc8051_indi_addr1_buff_4__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n93), .Y(oc8051_indi_addr1_n67)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u66 ( .A(wr_addr[0]), .B(
        oc8051_indi_addr1_n92), .C(oc8051_indi_addr1_n24), .Y(
        oc8051_indi_addr1_n27) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u65 ( .A(oc8051_indi_addr1_buff_5__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n68)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u64 ( .A(oc8051_indi_addr1_buff_5__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n69)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u63 ( .A(oc8051_indi_addr1_buff_5__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n70)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u62 ( .A(oc8051_indi_addr1_buff_5__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n71)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u61 ( .A(oc8051_indi_addr1_buff_5__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n72)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u60 ( .A(oc8051_indi_addr1_buff_5__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n73)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u59 ( .A(oc8051_indi_addr1_buff_5__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n74)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u58 ( .A(oc8051_indi_addr1_buff_5__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n27), .Y(oc8051_indi_addr1_n75)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u57 ( .A(wr_addr[3]), .B(
        oc8051_indi_addr1_n26), .C(oc8051_indi_addr1_n24), .Y(
        oc8051_indi_addr1_n25) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u56 ( .A(oc8051_indi_addr1_buff_6__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n76)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u55 ( .A(oc8051_indi_addr1_buff_6__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n77)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u54 ( .A(oc8051_indi_addr1_buff_6__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n78)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u53 ( .A(oc8051_indi_addr1_buff_6__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n79)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u52 ( .A(oc8051_indi_addr1_buff_6__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n80)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u51 ( .A(oc8051_indi_addr1_buff_6__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n81)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u50 ( .A(oc8051_indi_addr1_buff_6__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n82)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u49 ( .A(oc8051_indi_addr1_buff_6__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n25), .Y(oc8051_indi_addr1_n83)
         );
  AND3_X0P5M_A12TS oc8051_indi_addr1_u48 ( .A(wr_addr[3]), .B(wr_addr[0]), .C(
        oc8051_indi_addr1_n24), .Y(oc8051_indi_addr1_n23) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u47 ( .A(oc8051_indi_addr1_buff_7__7_), 
        .B(wr_dat[7]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n84)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u46 ( .A(oc8051_indi_addr1_buff_7__6_), 
        .B(wr_dat[6]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n85)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u45 ( .A(oc8051_indi_addr1_buff_7__5_), 
        .B(wr_dat[5]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n86)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u44 ( .A(oc8051_indi_addr1_buff_7__4_), 
        .B(wr_dat[4]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n87)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u43 ( .A(oc8051_indi_addr1_buff_7__3_), 
        .B(wr_dat[3]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n88)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u42 ( .A(oc8051_indi_addr1_buff_7__2_), 
        .B(wr_dat[2]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n89)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u41 ( .A(oc8051_indi_addr1_buff_7__1_), 
        .B(wr_dat[1]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n90)
         );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u40 ( .A(oc8051_indi_addr1_buff_7__0_), 
        .B(wr_dat[0]), .S0(oc8051_indi_addr1_n23), .Y(oc8051_indi_addr1_n91)
         );
  XNOR2_X0P5M_A12TS oc8051_indi_addr1_u39 ( .A(wr_addr[4]), .B(bank_sel[1]), 
        .Y(oc8051_indi_addr1_n19) );
  XNOR2_X0P5M_A12TS oc8051_indi_addr1_u38 ( .A(wr_addr[3]), .B(bank_sel[0]), 
        .Y(oc8051_indi_addr1_n20) );
  XNOR2_X0P5M_A12TS oc8051_indi_addr1_u37 ( .A(wr_addr[0]), .B(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n21) );
  NAND4_X0P5A_A12TS oc8051_indi_addr1_u36 ( .A(oc8051_indi_addr1_n19), .B(
        oc8051_indi_addr1_n20), .C(oc8051_indi_addr1_n21), .D(
        oc8051_indi_addr1_n22), .Y(oc8051_indi_addr1_n18) );
  OR6_X0P5M_A12TS oc8051_indi_addr1_u35 ( .A(wr_addr[7]), .B(wr_addr[6]), .C(
        wr_addr[5]), .D(wr_addr[2]), .E(wr_addr[1]), .F(oc8051_indi_addr1_n18), 
        .Y(oc8051_indi_addr1_n17) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u34 ( .A(wr_dat[0]), .B(
        oc8051_indi_addr1_n106), .S0(oc8051_indi_addr1_n17), .Y(ri[0]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u33 ( .A(wr_dat[1]), .B(
        oc8051_indi_addr1_n105), .S0(oc8051_indi_addr1_n17), .Y(ri[1]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u32 ( .A(wr_dat[2]), .B(
        oc8051_indi_addr1_n104), .S0(oc8051_indi_addr1_n17), .Y(ri[2]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u31 ( .A(wr_dat[3]), .B(
        oc8051_indi_addr1_n103), .S0(oc8051_indi_addr1_n17), .Y(ri[3]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u30 ( .A(wr_dat[4]), .B(
        oc8051_indi_addr1_n102), .S0(oc8051_indi_addr1_n17), .Y(ri[4]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u29 ( .A(wr_dat[5]), .B(
        oc8051_indi_addr1_n101), .S0(oc8051_indi_addr1_n17), .Y(ri[5]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u28 ( .A(wr_dat[6]), .B(
        oc8051_indi_addr1_n100), .S0(oc8051_indi_addr1_n17), .Y(ri[6]) );
  MXT2_X0P5M_A12TS oc8051_indi_addr1_u27 ( .A(wr_dat[7]), .B(
        oc8051_indi_addr1_n99), .S0(oc8051_indi_addr1_n17), .Y(ri[7]) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u26 ( .A(oc8051_indi_addr1_n15), .B(
        oc8051_indi_addr1_n16), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n106)
         );
  MXT2_X1M_A12TS oc8051_indi_addr1_u25 ( .A(oc8051_indi_addr1_n13), .B(
        oc8051_indi_addr1_n14), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n104)
         );
  MXT2_X1M_A12TS oc8051_indi_addr1_u24 ( .A(oc8051_indi_addr1_n11), .B(
        oc8051_indi_addr1_n12), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n105)
         );
  MXT2_X1M_A12TS oc8051_indi_addr1_u23 ( .A(oc8051_indi_addr1_n9), .B(
        oc8051_indi_addr1_n10), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n100)
         );
  MXT2_X1M_A12TS oc8051_indi_addr1_u22 ( .A(oc8051_indi_addr1_n7), .B(
        oc8051_indi_addr1_n8), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n101) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u21 ( .A(oc8051_indi_addr1_n5), .B(
        oc8051_indi_addr1_n6), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n102) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u20 ( .A(oc8051_indi_addr1_n3), .B(
        oc8051_indi_addr1_n4), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n99) );
  MXT2_X1M_A12TS oc8051_indi_addr1_u19 ( .A(oc8051_indi_addr1_n1), .B(
        oc8051_indi_addr1_n2), .S0(bank_sel[1]), .Y(oc8051_indi_addr1_n103) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u18 ( .A(oc8051_indi_addr1_buff_0__0_), 
        .B(oc8051_indi_addr1_buff_2__0_), .C(oc8051_indi_addr1_buff_1__0_), 
        .D(oc8051_indi_addr1_buff_3__0_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n15) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u17 ( .A(oc8051_indi_addr1_buff_4__0_), 
        .B(oc8051_indi_addr1_buff_6__0_), .C(oc8051_indi_addr1_buff_5__0_), 
        .D(oc8051_indi_addr1_buff_7__0_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n16) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u16 ( .A(oc8051_indi_addr1_buff_0__2_), 
        .B(oc8051_indi_addr1_buff_2__2_), .C(oc8051_indi_addr1_buff_1__2_), 
        .D(oc8051_indi_addr1_buff_3__2_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n13) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u15 ( .A(oc8051_indi_addr1_buff_4__2_), 
        .B(oc8051_indi_addr1_buff_6__2_), .C(oc8051_indi_addr1_buff_5__2_), 
        .D(oc8051_indi_addr1_buff_7__2_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n14) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u14 ( .A(oc8051_indi_addr1_buff_0__1_), 
        .B(oc8051_indi_addr1_buff_2__1_), .C(oc8051_indi_addr1_buff_1__1_), 
        .D(oc8051_indi_addr1_buff_3__1_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n11) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u13 ( .A(oc8051_indi_addr1_buff_4__1_), 
        .B(oc8051_indi_addr1_buff_6__1_), .C(oc8051_indi_addr1_buff_5__1_), 
        .D(oc8051_indi_addr1_buff_7__1_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n12) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u12 ( .A(oc8051_indi_addr1_buff_0__6_), 
        .B(oc8051_indi_addr1_buff_2__6_), .C(oc8051_indi_addr1_buff_1__6_), 
        .D(oc8051_indi_addr1_buff_3__6_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n9) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u11 ( .A(oc8051_indi_addr1_buff_4__6_), 
        .B(oc8051_indi_addr1_buff_6__6_), .C(oc8051_indi_addr1_buff_5__6_), 
        .D(oc8051_indi_addr1_buff_7__6_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n10) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u10 ( .A(oc8051_indi_addr1_buff_0__5_), 
        .B(oc8051_indi_addr1_buff_2__5_), .C(oc8051_indi_addr1_buff_1__5_), 
        .D(oc8051_indi_addr1_buff_3__5_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n7) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u9 ( .A(oc8051_indi_addr1_buff_4__5_), 
        .B(oc8051_indi_addr1_buff_6__5_), .C(oc8051_indi_addr1_buff_5__5_), 
        .D(oc8051_indi_addr1_buff_7__5_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n8) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u8 ( .A(oc8051_indi_addr1_buff_0__4_), 
        .B(oc8051_indi_addr1_buff_2__4_), .C(oc8051_indi_addr1_buff_1__4_), 
        .D(oc8051_indi_addr1_buff_3__4_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n5) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u7 ( .A(oc8051_indi_addr1_buff_4__4_), 
        .B(oc8051_indi_addr1_buff_6__4_), .C(oc8051_indi_addr1_buff_5__4_), 
        .D(oc8051_indi_addr1_buff_7__4_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n6) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u6 ( .A(oc8051_indi_addr1_buff_0__7_), 
        .B(oc8051_indi_addr1_buff_2__7_), .C(oc8051_indi_addr1_buff_1__7_), 
        .D(oc8051_indi_addr1_buff_3__7_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n3) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u5 ( .A(oc8051_indi_addr1_buff_4__7_), 
        .B(oc8051_indi_addr1_buff_6__7_), .C(oc8051_indi_addr1_buff_5__7_), 
        .D(oc8051_indi_addr1_buff_7__7_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n4) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u4 ( .A(oc8051_indi_addr1_buff_0__3_), 
        .B(oc8051_indi_addr1_buff_2__3_), .C(oc8051_indi_addr1_buff_1__3_), 
        .D(oc8051_indi_addr1_buff_3__3_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n1) );
  MXT4_X0P5M_A12TS oc8051_indi_addr1_u3 ( .A(oc8051_indi_addr1_buff_4__3_), 
        .B(oc8051_indi_addr1_buff_6__3_), .C(oc8051_indi_addr1_buff_5__3_), 
        .D(oc8051_indi_addr1_buff_7__3_), .S0(bank_sel[0]), .S1(op1_cur[0]), 
        .Y(oc8051_indi_addr1_n2) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__0_ ( .D(oc8051_indi_addr1_n83), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__1_ ( .D(oc8051_indi_addr1_n82), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__2_ ( .D(oc8051_indi_addr1_n81), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__3_ ( .D(oc8051_indi_addr1_n80), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__4_ ( .D(oc8051_indi_addr1_n79), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__5_ ( .D(oc8051_indi_addr1_n78), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__6_ ( .D(oc8051_indi_addr1_n77), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_6__7_ ( .D(oc8051_indi_addr1_n76), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_6__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__0_ ( .D(oc8051_indi_addr1_n51), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__1_ ( .D(oc8051_indi_addr1_n50), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__2_ ( .D(oc8051_indi_addr1_n49), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__3_ ( .D(oc8051_indi_addr1_n48), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__4_ ( .D(oc8051_indi_addr1_n47), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__5_ ( .D(oc8051_indi_addr1_n46), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__6_ ( .D(oc8051_indi_addr1_n45), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_2__7_ ( .D(oc8051_indi_addr1_n44), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_2__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__0_ ( .D(oc8051_indi_addr1_n67), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__1_ ( .D(oc8051_indi_addr1_n66), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__2_ ( .D(oc8051_indi_addr1_n65), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__3_ ( .D(oc8051_indi_addr1_n64), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__4_ ( .D(oc8051_indi_addr1_n63), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__5_ ( .D(oc8051_indi_addr1_n62), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__6_ ( .D(oc8051_indi_addr1_n61), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_4__7_ ( .D(oc8051_indi_addr1_n60), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_4__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__0_ ( .D(oc8051_indi_addr1_n35), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__1_ ( .D(oc8051_indi_addr1_n34), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__2_ ( .D(oc8051_indi_addr1_n33), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__3_ ( .D(oc8051_indi_addr1_n32), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__4_ ( .D(oc8051_indi_addr1_n31), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__5_ ( .D(oc8051_indi_addr1_n30), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__6_ ( .D(oc8051_indi_addr1_n29), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_0__7_ ( .D(oc8051_indi_addr1_n28), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_0__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__0_ ( .D(oc8051_indi_addr1_n75), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__1_ ( .D(oc8051_indi_addr1_n74), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__2_ ( .D(oc8051_indi_addr1_n73), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__3_ ( .D(oc8051_indi_addr1_n72), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__4_ ( .D(oc8051_indi_addr1_n71), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__5_ ( .D(oc8051_indi_addr1_n70), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__6_ ( .D(oc8051_indi_addr1_n69), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_5__7_ ( .D(oc8051_indi_addr1_n68), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_5__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__0_ ( .D(oc8051_indi_addr1_n43), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__1_ ( .D(oc8051_indi_addr1_n42), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__2_ ( .D(oc8051_indi_addr1_n41), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__3_ ( .D(oc8051_indi_addr1_n40), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__4_ ( .D(oc8051_indi_addr1_n39), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__5_ ( .D(oc8051_indi_addr1_n38), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__6_ ( .D(oc8051_indi_addr1_n37), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_1__7_ ( .D(oc8051_indi_addr1_n36), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_1__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__0_ ( .D(oc8051_indi_addr1_n91), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__1_ ( .D(oc8051_indi_addr1_n90), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__2_ ( .D(oc8051_indi_addr1_n89), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__3_ ( .D(oc8051_indi_addr1_n88), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__4_ ( .D(oc8051_indi_addr1_n87), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__5_ ( .D(oc8051_indi_addr1_n86), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__6_ ( .D(oc8051_indi_addr1_n85), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_7__7_ ( .D(oc8051_indi_addr1_n84), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_7__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__0_ ( .D(oc8051_indi_addr1_n59), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__0_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__1_ ( .D(oc8051_indi_addr1_n58), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__1_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__2_ ( .D(oc8051_indi_addr1_n57), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__2_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__3_ ( .D(oc8051_indi_addr1_n56), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__3_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__4_ ( .D(oc8051_indi_addr1_n55), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__4_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__5_ ( .D(oc8051_indi_addr1_n54), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__5_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__6_ ( .D(oc8051_indi_addr1_n53), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__6_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_buff_reg_3__7_ ( .D(oc8051_indi_addr1_n52), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_buff_3__7_) );
  DFFRPQ_X1M_A12TS oc8051_indi_addr1_wr_bit_r_reg ( .D(bit_addr_o), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_indi_addr1_wr_bit_r) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u888 ( .AN(mem_act[0]), .B(
        wbd_ack_i), .Y(oc8051_memory_interface1_n1310) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u887 ( .A(
        oc8051_memory_interface1_op1_5_), .Y(oc8051_memory_interface1_n772) );
  OR3_X0P5M_A12TS oc8051_memory_interface1_u886 ( .A(
        oc8051_memory_interface1_dmem_wait), .B(
        oc8051_memory_interface1_pc_wr_r2), .C(
        oc8051_memory_interface1_imem_wait), .Y(mem_wait) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u885 ( .A(rd), .Y(
        oc8051_memory_interface1_n186) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u884 ( .A(
        oc8051_memory_interface1_int_ack_t), .Y(oc8051_memory_interface1_n185)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u883 ( .A(wbi_cyc_o), .B(ea_in), 
        .Y(oc8051_memory_interface1_n167) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u882 ( .A(
        oc8051_memory_interface1_n167), .Y(oc8051_memory_interface1_n168) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u881 ( .A(wbi_ack_i), .B(
        oc8051_memory_interface1_n168), .Y(oc8051_memory_interface1_n187) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u880 ( .A(
        oc8051_memory_interface1_n185), .B(oc8051_memory_interface1_n187), .Y(
        oc8051_memory_interface1_n387) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u879 ( .A(
        oc8051_memory_interface1_n186), .B(oc8051_memory_interface1_n387), .Y(
        oc8051_memory_interface1_n718) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u878 ( .A(
        oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n716) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u877 ( .A(
        oc8051_memory_interface1_n772), .B(mem_wait), .C(
        oc8051_memory_interface1_n716), .Y(oc8051_memory_interface1_n769) );
  OR3_X0P5M_A12TS oc8051_memory_interface1_u876 ( .A(
        oc8051_memory_interface1_op1_6_), .B(oc8051_memory_interface1_op1_7_), 
        .C(oc8051_memory_interface1_op1_3_), .Y(oc8051_memory_interface1_n771)
         );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u875 ( .A(
        oc8051_memory_interface1_n771), .B(oc8051_memory_interface1_op1_2_), 
        .C(oc8051_memory_interface1_op1_0_), .Y(oc8051_memory_interface1_n770)
         );
  AND4_X0P5M_A12TS oc8051_memory_interface1_u874 ( .A(
        oc8051_memory_interface1_op1_4_), .B(oc8051_memory_interface1_op1_1_), 
        .C(oc8051_memory_interface1_n769), .D(oc8051_memory_interface1_n770), 
        .Y(oc8051_memory_interface1_n2000) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u873 ( .AN(
        oc8051_memory_interface1_int_ack_buff), .B(
        oc8051_memory_interface1_int_ack_t), .Y(oc8051_memory_interface1_n3720) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u872 ( .A(pc_wr_sel[2]), .Y(
        oc8051_memory_interface1_n652) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u871 ( .A(pc_wr_sel[1]), .Y(
        oc8051_memory_interface1_n653) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u870 ( .A(
        oc8051_memory_interface1_n652), .B(oc8051_memory_interface1_n653), .Y(
        oc8051_memory_interface1_n614) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u869 ( .A(
        oc8051_memory_interface1_n614), .Y(oc8051_memory_interface1_n667) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u868 ( .A(n_3_net_), .Y(
        oc8051_memory_interface1_n601) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u867 ( .A(pc_wr_sel[0]), .Y(
        oc8051_memory_interface1_n603) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u866 ( .A(n_3_net_), .B(
        oc8051_memory_interface1_n603), .Y(oc8051_memory_interface1_n655) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u865 ( .A0(
        oc8051_memory_interface1_n667), .A1(oc8051_memory_interface1_n601), 
        .B0(oc8051_memory_interface1_n655), .Y(oc8051_memory_interface1_n5530)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u864 ( .A(ram_rd_sel[0]), .Y(
        oc8051_memory_interface1_n113) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u863 ( .A(
        oc8051_memory_interface1_n113), .B(ram_rd_sel[2]), .Y(
        oc8051_memory_interface1_n830) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u862 ( .A(ram_wr_sel[1]), .Y(
        oc8051_memory_interface1_n86) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u861 ( .A(
        oc8051_memory_interface1_n86), .B(ram_wr_sel[2]), .Y(wr_ind) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u860 ( .AN(
        oc8051_memory_interface1_rd_addr_r), .B(
        oc8051_memory_interface1_rd_ind), .Y(oc8051_memory_interface1_n736) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u859 ( .A(bit_data), .B(sfr_bit), 
        .S0(oc8051_memory_interface1_n736), .Y(bit_out) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u858 ( .A(
        oc8051_memory_interface1_istb_t), .Y(oc8051_memory_interface1_n172) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u857 ( .A(
        oc8051_memory_interface1_iadr_t_0_), .Y(oc8051_memory_interface1_n734)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u856 ( .A(
        oc8051_memory_interface1_pc_wr_r2), .Y(oc8051_memory_interface1_n197)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u855 ( .A0(
        oc8051_memory_interface1_op_pos_1_), .A1(
        oc8051_memory_interface1_op_pos_0_), .B0(
        oc8051_memory_interface1_op_pos_2_), .C0(rd), .Y(
        oc8051_memory_interface1_n768) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u854 ( .A(
        oc8051_memory_interface1_n197), .B(oc8051_memory_interface1_n768), .Y(
        oc8051_memory_interface1_n194) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u853 ( .A(
        oc8051_memory_interface1_n200), .B(oc8051_memory_interface1_n172), .Y(
        oc8051_memory_interface1_n744) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u852 ( .A(
        oc8051_memory_interface1_n744), .Y(oc8051_memory_interface1_n738) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u851 ( .A(
        oc8051_memory_interface1_n172), .B(oc8051_memory_interface1_n194), .Y(
        oc8051_memory_interface1_n745) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u850 ( .A(
        oc8051_memory_interface1_n745), .Y(oc8051_memory_interface1_n739) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u849 ( .A(
        oc8051_memory_interface1_n738), .B(oc8051_memory_interface1_n739), .Y(
        oc8051_memory_interface1_n755) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u848 ( .A(
        oc8051_memory_interface1_pc_buf_0_), .Y(oc8051_memory_interface1_n239)
         );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u847 ( .A0(
        oc8051_memory_interface1_n172), .A1(oc8051_memory_interface1_n734), 
        .B0(oc8051_memory_interface1_n755), .B1(oc8051_memory_interface1_n239), 
        .Y(wbi_adr_o[0]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u846 ( .A(
        oc8051_memory_interface1_pc_buf_10_), .Y(oc8051_memory_interface1_n292) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u845 ( .A(
        oc8051_memory_interface1_pc_buf_9_), .Y(oc8051_memory_interface1_n287)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u844 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .Y(oc8051_memory_interface1_n254)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u843 ( .A(
        oc8051_memory_interface1_pc_buf_2_), .Y(oc8051_memory_interface1_n249)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u842 ( .A(
        oc8051_memory_interface1_pc_buf_4_), .Y(oc8051_memory_interface1_n259)
         );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u841 ( .A(
        oc8051_memory_interface1_n254), .B(oc8051_memory_interface1_n249), .C(
        oc8051_memory_interface1_n259), .Y(oc8051_memory_interface1_n749) );
  AND3_X0P5M_A12TS oc8051_memory_interface1_u840 ( .A(
        oc8051_memory_interface1_pc_buf_6_), .B(
        oc8051_memory_interface1_pc_buf_5_), .C(oc8051_memory_interface1_n749), 
        .Y(oc8051_memory_interface1_n743) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u839 ( .A(
        oc8051_memory_interface1_pc_buf_8_), .B(
        oc8051_memory_interface1_pc_buf_7_), .C(oc8051_memory_interface1_n743), 
        .Y(oc8051_memory_interface1_n740) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u838 ( .A(
        oc8051_memory_interface1_n287), .B(oc8051_memory_interface1_n740), .Y(
        oc8051_memory_interface1_n767) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u837 ( .A(
        oc8051_memory_interface1_n292), .B(oc8051_memory_interface1_n767), .Y(
        oc8051_memory_interface1_n643) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u836 ( .A0(
        oc8051_memory_interface1_pc_buf_10_), .A1(
        oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n643), 
        .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_10_), .Y(oc8051_memory_interface1_n766) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u835 ( .A(
        oc8051_memory_interface1_n766), .Y(wbi_adr_o[10]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u834 ( .A(
        oc8051_memory_interface1_pc_buf_11_), .Y(oc8051_memory_interface1_n297) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u833 ( .A(
        oc8051_memory_interface1_n292), .B(oc8051_memory_interface1_n287), .C(
        oc8051_memory_interface1_n740), .Y(oc8051_memory_interface1_n762) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u832 ( .A(
        oc8051_memory_interface1_n297), .B(oc8051_memory_interface1_n762), .Y(
        oc8051_memory_interface1_n660) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u831 ( .A0(
        oc8051_memory_interface1_pc_buf_11_), .A1(
        oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n660), 
        .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_11_), .Y(oc8051_memory_interface1_n765) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u830 ( .A(
        oc8051_memory_interface1_n765), .Y(wbi_adr_o[11]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u829 ( .A(
        oc8051_memory_interface1_pc_buf_12_), .Y(oc8051_memory_interface1_n302) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u828 ( .A(
        oc8051_memory_interface1_n762), .B(oc8051_memory_interface1_pc_buf_11_), .Y(oc8051_memory_interface1_n764) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u827 ( .A(
        oc8051_memory_interface1_n764), .B(oc8051_memory_interface1_pc_buf_12_), .Y(oc8051_memory_interface1_n669) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u826 ( .A(
        oc8051_memory_interface1_iadr_t_12_), .Y(oc8051_memory_interface1_n763) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u825 ( .A0(
        oc8051_memory_interface1_n302), .A1(oc8051_memory_interface1_n744), 
        .B0(oc8051_memory_interface1_n669), .B1(oc8051_memory_interface1_n745), 
        .C0(oc8051_memory_interface1_n172), .C1(oc8051_memory_interface1_n763), 
        .Y(wbi_adr_o[12]) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u824 ( .A(
        oc8051_memory_interface1_pc_buf_12_), .B(
        oc8051_memory_interface1_pc_buf_11_), .C(oc8051_memory_interface1_n762), .Y(oc8051_memory_interface1_n760) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u823 ( .A(
        oc8051_memory_interface1_pc_buf_13_), .Y(oc8051_memory_interface1_n307) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u822 ( .A(
        oc8051_memory_interface1_n760), .B(oc8051_memory_interface1_n307), .Y(
        oc8051_memory_interface1_n681) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u821 ( .A0(
        oc8051_memory_interface1_pc_buf_13_), .A1(
        oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n681), 
        .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_13_), .Y(oc8051_memory_interface1_n761) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u820 ( .A(
        oc8051_memory_interface1_n761), .Y(wbi_adr_o[13]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u819 ( .A(
        oc8051_memory_interface1_pc_buf_14_), .Y(oc8051_memory_interface1_n313) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u818 ( .A(
        oc8051_memory_interface1_n760), .B(oc8051_memory_interface1_n307), .Y(
        oc8051_memory_interface1_n758) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u817 ( .A(
        oc8051_memory_interface1_n313), .B(oc8051_memory_interface1_n758), .Y(
        oc8051_memory_interface1_n692) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u816 ( .A0(
        oc8051_memory_interface1_pc_buf_14_), .A1(
        oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n692), 
        .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_14_), .Y(oc8051_memory_interface1_n759) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u815 ( .A(
        oc8051_memory_interface1_n759), .Y(wbi_adr_o[14]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u814 ( .A(
        oc8051_memory_interface1_n758), .B(oc8051_memory_interface1_pc_buf_14_), .Y(oc8051_memory_interface1_n757) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u813 ( .A(
        oc8051_memory_interface1_n757), .B(oc8051_memory_interface1_pc_buf_15_), .Y(oc8051_memory_interface1_n701) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u812 ( .A0(
        oc8051_memory_interface1_pc_buf_15_), .A1(
        oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n701), 
        .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_15_), .Y(oc8051_memory_interface1_n756) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u811 ( .A(
        oc8051_memory_interface1_n756), .Y(wbi_adr_o[15]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u810 ( .A(
        oc8051_memory_interface1_iadr_t_1_), .Y(oc8051_memory_interface1_n733)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u809 ( .A(
        oc8051_memory_interface1_pc_buf_1_), .Y(oc8051_memory_interface1_n243)
         );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u808 ( .A0(
        oc8051_memory_interface1_n172), .A1(oc8051_memory_interface1_n733), 
        .B0(oc8051_memory_interface1_n755), .B1(oc8051_memory_interface1_n243), 
        .Y(wbi_adr_o[1]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u807 ( .A(
        oc8051_memory_interface1_iadr_t_2_), .Y(oc8051_memory_interface1_n732)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u806 ( .A(
        oc8051_memory_interface1_n739), .B(oc8051_memory_interface1_n738), 
        .S0(oc8051_memory_interface1_pc_buf_2_), .Y(
        oc8051_memory_interface1_n754) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u805 ( .A0(
        oc8051_memory_interface1_n172), .A1(oc8051_memory_interface1_n732), 
        .B0(oc8051_memory_interface1_n754), .Y(wbi_adr_o[2]) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u804 ( .A(
        oc8051_memory_interface1_n249), .B(oc8051_memory_interface1_n254), .Y(
        oc8051_memory_interface1_n439) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u803 ( .A0(
        oc8051_memory_interface1_pc_buf_3_), .A1(oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n439), .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_3_), .Y(oc8051_memory_interface1_n753)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u802 ( .A(
        oc8051_memory_interface1_n753), .Y(wbi_adr_o[3]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u801 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .B(
        oc8051_memory_interface1_pc_buf_2_), .Y(oc8051_memory_interface1_n752)
         );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u800 ( .A(
        oc8051_memory_interface1_n752), .B(oc8051_memory_interface1_pc_buf_4_), 
        .Y(oc8051_memory_interface1_n546) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u799 ( .A0(
        oc8051_memory_interface1_pc_buf_4_), .A1(oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n546), .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_4_), .Y(oc8051_memory_interface1_n751)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u798 ( .A(
        oc8051_memory_interface1_n751), .Y(wbi_adr_o[4]) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u797 ( .A(
        oc8051_memory_interface1_n749), .B(oc8051_memory_interface1_pc_buf_5_), 
        .Y(oc8051_memory_interface1_n587) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u796 ( .A0(
        oc8051_memory_interface1_pc_buf_5_), .A1(oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n587), .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_5_), .Y(oc8051_memory_interface1_n750)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u795 ( .A(
        oc8051_memory_interface1_n750), .Y(wbi_adr_o[5]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u794 ( .A(
        oc8051_memory_interface1_pc_buf_6_), .Y(oc8051_memory_interface1_n271)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u793 ( .A(
        oc8051_memory_interface1_pc_buf_5_), .Y(oc8051_memory_interface1_n265)
         );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u792 ( .AN(
        oc8051_memory_interface1_n749), .B(oc8051_memory_interface1_n265), .Y(
        oc8051_memory_interface1_n748) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u791 ( .A(
        oc8051_memory_interface1_n271), .B(oc8051_memory_interface1_n748), .Y(
        oc8051_memory_interface1_n594) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u790 ( .A0(
        oc8051_memory_interface1_pc_buf_6_), .A1(oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n594), .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_6_), .Y(oc8051_memory_interface1_n747)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u789 ( .A(
        oc8051_memory_interface1_n747), .Y(wbi_adr_o[6]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u788 ( .A(
        oc8051_memory_interface1_pc_buf_7_), .Y(oc8051_memory_interface1_n277)
         );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u787 ( .A(
        oc8051_memory_interface1_n277), .B(oc8051_memory_interface1_n743), .Y(
        oc8051_memory_interface1_n599) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u786 ( .A(
        oc8051_memory_interface1_iadr_t_7_), .Y(oc8051_memory_interface1_n746)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u785 ( .A0(
        oc8051_memory_interface1_n277), .A1(oc8051_memory_interface1_n744), 
        .B0(oc8051_memory_interface1_n599), .B1(oc8051_memory_interface1_n745), 
        .C0(oc8051_memory_interface1_n172), .C1(oc8051_memory_interface1_n746), 
        .Y(wbi_adr_o[7]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u784 ( .A(
        oc8051_memory_interface1_n743), .B(oc8051_memory_interface1_pc_buf_7_), 
        .Y(oc8051_memory_interface1_n742) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u783 ( .A(
        oc8051_memory_interface1_n742), .B(oc8051_memory_interface1_pc_buf_8_), 
        .Y(oc8051_memory_interface1_n619) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u782 ( .A0(
        oc8051_memory_interface1_pc_buf_8_), .A1(oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n619), .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_8_), .Y(oc8051_memory_interface1_n741)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u781 ( .A(
        oc8051_memory_interface1_n741), .Y(wbi_adr_o[8]) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u780 ( .A(
        oc8051_memory_interface1_n740), .B(oc8051_memory_interface1_n287), .Y(
        oc8051_memory_interface1_n632) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u779 ( .A0(
        oc8051_memory_interface1_pc_buf_9_), .A1(oc8051_memory_interface1_n738), .B0(oc8051_memory_interface1_n632), .B1(oc8051_memory_interface1_n739), .C0(
        oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_iadr_t_9_), .Y(oc8051_memory_interface1_n737)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u778 ( .A(
        oc8051_memory_interface1_n737), .Y(wbi_adr_o[9]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u777 ( .A(ram_data[0]), .B(
        sfr_out[0]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[0]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u776 ( .A(ram_data[1]), .B(
        sfr_out[1]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[1]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u775 ( .A(ram_data[2]), .B(
        sfr_out[2]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[2]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u774 ( .A(ram_data[3]), .B(
        sfr_out[3]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[3]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u773 ( .A(ram_data[4]), .B(
        sfr_out[4]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[4]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u772 ( .A(ram_data[5]), .B(
        sfr_out[5]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[5]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u771 ( .A(ram_data[6]), .B(
        sfr_out[6]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[6]) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u770 ( .A(ram_data[7]), .B(
        sfr_out[7]), .S0(oc8051_memory_interface1_n736), .Y(ram_out[7]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u769 ( .A(
        oc8051_memory_interface1_n187), .Y(oc8051_memory_interface1_n169) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u768 ( .A(istb), .B(
        oc8051_memory_interface1_n167), .Y(oc8051_memory_interface1_n735) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u767 ( .A0(
        oc8051_memory_interface1_n172), .A1(oc8051_memory_interface1_n169), 
        .B0(oc8051_memory_interface1_n735), .C0(wbd_cyc_o), .Y(
        oc8051_memory_interface1_istb_o) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u766 ( .A(
        oc8051_memory_interface1_ddat_ir_0_), .B(wbd_dat_i[0]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n416) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u765 ( .A(
        oc8051_memory_interface1_ddat_ir_1_), .B(wbd_dat_i[1]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n417) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u764 ( .A(
        oc8051_memory_interface1_ddat_ir_2_), .B(wbd_dat_i[2]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n418) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u763 ( .A(
        oc8051_memory_interface1_ddat_ir_3_), .B(wbd_dat_i[3]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n419) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u762 ( .A(
        oc8051_memory_interface1_ddat_ir_4_), .B(wbd_dat_i[4]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n420) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u761 ( .A(
        oc8051_memory_interface1_ddat_ir_5_), .B(wbd_dat_i[5]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n421) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u760 ( .A(
        oc8051_memory_interface1_ddat_ir_6_), .B(wbd_dat_i[6]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n422) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u759 ( .A(
        oc8051_memory_interface1_ddat_ir_7_), .B(wbd_dat_i[7]), .S0(wbd_ack_i), 
        .Y(oc8051_memory_interface1_n423) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u758 ( .A(
        oc8051_memory_interface1_int_vec_buff_0_), .B(int_src[0]), .S0(intr), 
        .Y(oc8051_memory_interface1_n424) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u757 ( .A(
        oc8051_memory_interface1_int_vec_buff_1_), .B(int_src[1]), .S0(intr), 
        .Y(oc8051_memory_interface1_n425) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u756 ( .A(
        oc8051_memory_interface1_int_vec_buff_2_), .B(n2), .S0(intr), .Y(
        oc8051_memory_interface1_n426) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u755 ( .A(
        oc8051_memory_interface1_int_vec_buff_3_), .B(int_src[3]), .S0(intr), 
        .Y(oc8051_memory_interface1_n427) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u754 ( .A(
        oc8051_memory_interface1_int_vec_buff_4_), .B(int_src[4]), .S0(intr), 
        .Y(oc8051_memory_interface1_n428) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u753 ( .A(
        oc8051_memory_interface1_int_vec_buff_5_), .B(int_src[5]), .S0(intr), 
        .Y(oc8051_memory_interface1_n429) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u752 ( .A(
        oc8051_memory_interface1_int_vec_buff_6_), .B(n2), .S0(intr), .Y(
        oc8051_memory_interface1_n430) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u751 ( .A(
        oc8051_memory_interface1_int_vec_buff_7_), .B(n2), .S0(intr), .Y(
        oc8051_memory_interface1_n431) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u750 ( .A(des_acc[0]), .Y(
        oc8051_memory_interface1_n623) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u749 ( .A(mem_act[1]), .Y(
        oc8051_memory_interface1_n183) );
  NAND3B_X0P5M_A12TS oc8051_memory_interface1_u748 ( .AN(mem_act[0]), .B(
        oc8051_memory_interface1_n183), .C(mem_act[2]), .Y(
        oc8051_memory_interface1_n171) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u747 ( .A(
        oc8051_memory_interface1_n623), .B(oc8051_memory_interface1_n734), 
        .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n440)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u746 ( .A(des_acc[1]), .Y(
        oc8051_memory_interface1_n635) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u745 ( .A(
        oc8051_memory_interface1_n635), .B(oc8051_memory_interface1_n733), 
        .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n441)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u744 ( .A(des_acc[2]), .Y(
        oc8051_memory_interface1_n646) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u743 ( .A(
        oc8051_memory_interface1_n646), .B(oc8051_memory_interface1_n732), 
        .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n442)
         );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u742 ( .A(des_acc[3]), .B(
        oc8051_memory_interface1_iadr_t_3_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n443) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u741 ( .A(des_acc[4]), .B(
        oc8051_memory_interface1_iadr_t_4_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n444) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u740 ( .A(des_acc[5]), .B(
        oc8051_memory_interface1_iadr_t_5_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n445) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u739 ( .A(des_acc[6]), .B(
        oc8051_memory_interface1_iadr_t_6_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n446) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u738 ( .A(des_acc[7]), .B(
        oc8051_memory_interface1_iadr_t_7_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n447) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u737 ( .A(des2[0]), .B(
        oc8051_memory_interface1_iadr_t_8_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n448) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u736 ( .A(des2[1]), .B(
        oc8051_memory_interface1_iadr_t_9_), .S0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n449) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u735 ( .A(des2[2]), .B(
        oc8051_memory_interface1_iadr_t_10_), .S0(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n450) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u734 ( .A(des2[3]), .B(
        oc8051_memory_interface1_iadr_t_11_), .S0(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n451) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u733 ( .A(des2[4]), .B(
        oc8051_memory_interface1_iadr_t_12_), .S0(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n452) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u732 ( .A(des2[5]), .B(
        oc8051_memory_interface1_iadr_t_13_), .S0(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n453) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u731 ( .A(des2[6]), .B(
        oc8051_memory_interface1_iadr_t_14_), .S0(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n454) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u730 ( .A(des2[7]), .B(
        oc8051_memory_interface1_iadr_t_15_), .S0(
        oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n455) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u729 ( .A(
        oc8051_memory_interface1_n399), .Y(pc[15]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u728 ( .A(
        oc8051_memory_interface1_n655), .B(pc_wr_sel[1]), .Y(
        oc8051_memory_interface1_n621) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u727 ( .A(
        oc8051_memory_interface1_n601), .B(oc8051_memory_interface1_n621), .Y(
        oc8051_memory_interface1_n687) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u726 ( .A(
        oc8051_memory_interface1_n653), .B(pc_wr_sel[2]), .Y(
        oc8051_memory_interface1_n597) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u725 ( .A0(
        oc8051_memory_interface1_op2_buff[7]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[7]), 
        .B1(oc8051_memory_interface1_n718), .Y(op2_n[7]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u724 ( .A(
        oc8051_memory_interface1_n387), .B(rd), .Y(
        oc8051_memory_interface1_n717) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u723 ( .A0(
        oc8051_memory_interface1_op3[7]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_7_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[7]), .Y(
        oc8051_memory_interface1_n731) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u722 ( .A(
        oc8051_memory_interface1_n731), .Y(op3_n[7]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u721 ( .A(op2_n[7]), .B(op3_n[7]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n708) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u720 ( .A(
        oc8051_memory_interface1_n708), .Y(oc8051_memory_interface1_n710) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u719 ( .A(
        oc8051_memory_interface1_n597), .B(oc8051_memory_interface1_n710), .Y(
        oc8051_memory_interface1_n628) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u718 ( .A(
        oc8051_memory_interface1_n628), .Y(oc8051_memory_interface1_n608) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u717 ( .A(
        oc8051_memory_interface1_n687), .B(oc8051_memory_interface1_n608), .Y(
        oc8051_memory_interface1_n665) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u716 ( .A(
        oc8051_memory_interface1_n665), .Y(oc8051_memory_interface1_n677) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u715 ( .A0(
        oc8051_memory_interface1_op2_buff[1]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[1]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n641)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u714 ( .A0(
        oc8051_memory_interface1_op3[1]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_1_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[1]), .Y(
        oc8051_memory_interface1_n414) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u713 ( .A(
        oc8051_memory_interface1_n641), .B(oc8051_memory_interface1_n414), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n729) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u712 ( .A0(
        oc8051_memory_interface1_op2_buff[0]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[0]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n127)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u711 ( .A(
        oc8051_memory_interface1_n127), .Y(op2_n[0]) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u710 ( .A0(
        oc8051_memory_interface1_op3[0]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_0_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[0]), .Y(
        oc8051_memory_interface1_n730) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u709 ( .A(
        oc8051_memory_interface1_n730), .Y(op3_n[0]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u708 ( .A(op2_n[0]), .B(op3_n[0]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n404) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u707 ( .A(pc[0]), .Y(
        oc8051_memory_interface1_n236) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u706 ( .A(
        oc8051_memory_interface1_n404), .B(oc8051_memory_interface1_n236), .Y(
        oc8051_memory_interface1_n412) );
  CGENI_X1M_A12TS oc8051_memory_interface1_u705 ( .A(
        oc8051_memory_interface1_n729), .B(pc[1]), .CI(
        oc8051_memory_interface1_n412), .CON(oc8051_memory_interface1_n434) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u704 ( .A0(
        oc8051_memory_interface1_op2_buff[2]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[2]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n121)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u703 ( .A(
        oc8051_memory_interface1_n121), .Y(op2_n[2]) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u702 ( .A0(
        oc8051_memory_interface1_op3[2]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_2_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[2]), .Y(
        oc8051_memory_interface1_n728) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u701 ( .A(
        oc8051_memory_interface1_n728), .Y(op3_n[2]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u700 ( .A(op2_n[2]), .B(op3_n[2]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n435) );
  AND2_X0P5M_A12TS oc8051_memory_interface1_u699 ( .A(
        oc8051_memory_interface1_n434), .B(oc8051_memory_interface1_n435), .Y(
        oc8051_memory_interface1_n727) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u698 ( .A(pc[2]), .Y(
        oc8051_memory_interface1_n247) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u697 ( .A0(
        oc8051_memory_interface1_n434), .A1(oc8051_memory_interface1_n435), 
        .B0(oc8051_memory_interface1_n727), .B1(oc8051_memory_interface1_n247), 
        .Y(oc8051_memory_interface1_n725) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u696 ( .A(
        oc8051_memory_interface1_n725), .Y(oc8051_memory_interface1_n456) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u695 ( .A0(
        oc8051_memory_interface1_op2_buff[3]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[3]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n118)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u694 ( .A(
        oc8051_memory_interface1_n118), .Y(op2_n[3]) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u693 ( .A0(
        oc8051_memory_interface1_op3[3]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_3_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[3]), .Y(
        oc8051_memory_interface1_n726) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u692 ( .A(
        oc8051_memory_interface1_n726), .Y(op3_n[3]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u691 ( .A(op2_n[3]), .B(op3_n[3]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n457) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u690 ( .AN(
        oc8051_memory_interface1_n457), .B(oc8051_memory_interface1_n725), .Y(
        oc8051_memory_interface1_n724) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u689 ( .A(pc[3]), .Y(
        oc8051_memory_interface1_n252) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u688 ( .A0(
        oc8051_memory_interface1_n456), .A1(oc8051_memory_interface1_n457), 
        .B0(oc8051_memory_interface1_n724), .B1(oc8051_memory_interface1_n252), 
        .Y(oc8051_memory_interface1_n548) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u687 ( .A0(
        oc8051_memory_interface1_op2_buff[4]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[4]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n114)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u686 ( .A(
        oc8051_memory_interface1_n114), .Y(op2_n[4]) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u685 ( .A0(
        oc8051_memory_interface1_op3[4]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_4_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[4]), .Y(
        oc8051_memory_interface1_n723) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u684 ( .A(
        oc8051_memory_interface1_n723), .Y(op3_n[4]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u683 ( .A(op2_n[4]), .B(op3_n[4]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n550) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u682 ( .A(
        oc8051_memory_interface1_n550), .Y(oc8051_memory_interface1_n721) );
  OR2_X0P5M_A12TS oc8051_memory_interface1_u681 ( .A(
        oc8051_memory_interface1_n548), .B(oc8051_memory_interface1_n721), .Y(
        oc8051_memory_interface1_n722) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u680 ( .A0(
        oc8051_memory_interface1_n548), .A1(oc8051_memory_interface1_n721), 
        .B0(oc8051_memory_interface1_n722), .B1(pc[4]), .Y(
        oc8051_memory_interface1_n589) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u679 ( .A0(
        oc8051_memory_interface1_op2_buff[5]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[5]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n109)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u678 ( .A(
        oc8051_memory_interface1_n109), .Y(op2_n[5]) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u677 ( .A0(
        oc8051_memory_interface1_op3[5]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_5_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[5]), .Y(
        oc8051_memory_interface1_n720) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u676 ( .A(
        oc8051_memory_interface1_n720), .Y(op3_n[5]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u675 ( .A(op2_n[5]), .B(op3_n[5]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n590) );
  AND2_X0P5M_A12TS oc8051_memory_interface1_u674 ( .A(
        oc8051_memory_interface1_n589), .B(oc8051_memory_interface1_n590), .Y(
        oc8051_memory_interface1_n719) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u673 ( .A(pc[5]), .Y(
        oc8051_memory_interface1_n263) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u672 ( .A0(
        oc8051_memory_interface1_n589), .A1(oc8051_memory_interface1_n590), 
        .B0(oc8051_memory_interface1_n719), .B1(oc8051_memory_interface1_n263), 
        .Y(oc8051_memory_interface1_n610) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u671 ( .A(
        oc8051_memory_interface1_n610), .Y(oc8051_memory_interface1_n595) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u670 ( .A0(
        oc8051_memory_interface1_op2_buff[6]), .A1(
        oc8051_memory_interface1_n186), .B0(oc8051_memory_interface1_op2[6]), 
        .B1(oc8051_memory_interface1_n718), .Y(oc8051_memory_interface1_n103)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u669 ( .A(
        oc8051_memory_interface1_n103), .Y(op2_n[6]) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u668 ( .A0(
        oc8051_memory_interface1_op3[6]), .A1(oc8051_memory_interface1_n716), 
        .B0(oc8051_memory_interface1_int_vec_buff_6_), .B1(
        oc8051_memory_interface1_n717), .C0(rd), .C1(
        oc8051_memory_interface1_op3_buff[6]), .Y(
        oc8051_memory_interface1_n715) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u667 ( .A(
        oc8051_memory_interface1_n715), .Y(op3_n[6]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u666 ( .A(op2_n[6]), .B(op3_n[6]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n612) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u665 ( .A(
        oc8051_memory_interface1_n612), .Y(oc8051_memory_interface1_n596) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u664 ( .A(
        oc8051_memory_interface1_n610), .B(oc8051_memory_interface1_n596), .Y(
        oc8051_memory_interface1_n714) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u663 ( .A(pc[6]), .Y(
        oc8051_memory_interface1_n269) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u662 ( .A0(
        oc8051_memory_interface1_n595), .A1(oc8051_memory_interface1_n612), 
        .B0(oc8051_memory_interface1_n714), .B1(oc8051_memory_interface1_n269), 
        .Y(oc8051_memory_interface1_n713) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u661 ( .A(
        oc8051_memory_interface1_n713), .Y(oc8051_memory_interface1_n711) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u660 ( .A(
        oc8051_memory_interface1_n710), .B(oc8051_memory_interface1_n713), .Y(
        oc8051_memory_interface1_n712) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u659 ( .A(pc[7]), .Y(
        oc8051_memory_interface1_n275) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u658 ( .A0(
        oc8051_memory_interface1_n711), .A1(oc8051_memory_interface1_n708), 
        .B0(oc8051_memory_interface1_n712), .B1(oc8051_memory_interface1_n275), 
        .Y(oc8051_memory_interface1_n707) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u657 ( .A(
        oc8051_memory_interface1_n398), .B(oc8051_memory_interface1_n710), .Y(
        oc8051_memory_interface1_n709) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u656 ( .A(
        oc8051_memory_interface1_n707), .B(oc8051_memory_interface1_n709), .Y(
        oc8051_memory_interface1_n630) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u655 ( .A(
        oc8051_memory_interface1_n398), .Y(pc[8]) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u654 ( .AN(
        oc8051_memory_interface1_n630), .B(pc[8]), .Y(
        oc8051_memory_interface1_n625) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u653 ( .A(
        oc8051_memory_interface1_n625), .B(oc8051_memory_interface1_n397), .Y(
        oc8051_memory_interface1_n639) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u652 ( .A(
        oc8051_memory_interface1_n396), .Y(pc[10]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u651 ( .A(
        oc8051_memory_interface1_n639), .B(pc[10]), .Y(
        oc8051_memory_interface1_n650) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u650 ( .A(
        oc8051_memory_interface1_n650), .B(oc8051_memory_interface1_n395), .Y(
        oc8051_memory_interface1_n664) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u649 ( .A(
        oc8051_memory_interface1_n394), .Y(pc[12]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u648 ( .A(
        oc8051_memory_interface1_n664), .B(pc[12]), .Y(
        oc8051_memory_interface1_n676) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u647 ( .A(
        oc8051_memory_interface1_n676), .B(oc8051_memory_interface1_n393), .Y(
        oc8051_memory_interface1_n684) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u646 ( .A(
        oc8051_memory_interface1_n684), .Y(oc8051_memory_interface1_n695) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u645 ( .A(
        oc8051_memory_interface1_n677), .B(oc8051_memory_interface1_n392), .C(
        oc8051_memory_interface1_n695), .Y(oc8051_memory_interface1_n696) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u644 ( .A(
        oc8051_memory_interface1_n708), .B(oc8051_memory_interface1_n597), .Y(
        oc8051_memory_interface1_n629) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u643 ( .A(
        oc8051_memory_interface1_n629), .Y(oc8051_memory_interface1_n607) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u642 ( .A(
        oc8051_memory_interface1_n687), .B(oc8051_memory_interface1_n607), .Y(
        oc8051_memory_interface1_n673) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u641 ( .A(
        oc8051_memory_interface1_n673), .Y(oc8051_memory_interface1_n661) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u640 ( .A(
        oc8051_memory_interface1_n707), .B(pc[8]), .Y(
        oc8051_memory_interface1_n640) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u639 ( .A(
        oc8051_memory_interface1_n640), .B(oc8051_memory_interface1_n397), .Y(
        oc8051_memory_interface1_n651) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u638 ( .A(
        oc8051_memory_interface1_n651), .B(pc[10]), .Y(
        oc8051_memory_interface1_n666) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u637 ( .A(
        oc8051_memory_interface1_n666), .B(oc8051_memory_interface1_n395), .Y(
        oc8051_memory_interface1_n678) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u636 ( .A(
        oc8051_memory_interface1_n678), .B(pc[12]), .Y(
        oc8051_memory_interface1_n685) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u635 ( .A(
        oc8051_memory_interface1_n685), .B(oc8051_memory_interface1_n393), .Y(
        oc8051_memory_interface1_n697) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u634 ( .A(
        oc8051_memory_interface1_n392), .Y(pc[14]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u633 ( .A(
        oc8051_memory_interface1_n697), .B(pc[14]), .Y(
        oc8051_memory_interface1_n705) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u632 ( .A(
        oc8051_memory_interface1_n661), .B(oc8051_memory_interface1_n705), .Y(
        oc8051_memory_interface1_n706) );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u631 ( .A0(
        oc8051_memory_interface1_n695), .A1(oc8051_memory_interface1_n392), 
        .B0(oc8051_memory_interface1_n665), .C0(oc8051_memory_interface1_n706), 
        .Y(oc8051_memory_interface1_n703) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u630 ( .A(
        oc8051_memory_interface1_n673), .B(oc8051_memory_interface1_n705), .Y(
        oc8051_memory_interface1_n704) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u629 ( .A(
        oc8051_memory_interface1_n703), .B(oc8051_memory_interface1_n704), 
        .S0(oc8051_memory_interface1_n399), .Y(oc8051_memory_interface1_n698)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u628 ( .A(
        oc8051_memory_interface1_n200), .B(oc8051_memory_interface1_n601), .Y(
        oc8051_memory_interface1_n604) );
  NAND2B_X0P5M_A12TS oc8051_memory_interface1_u627 ( .AN(
        oc8051_memory_interface1_n621), .B(oc8051_memory_interface1_n604), .Y(
        oc8051_memory_interface1_n686) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u626 ( .A(pc_wr_sel[2]), .B(
        pc_wr_sel[1]), .Y(oc8051_memory_interface1_n615) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u625 ( .A(
        oc8051_memory_interface1_n615), .Y(oc8051_memory_interface1_n668) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u624 ( .A(
        oc8051_memory_interface1_n652), .B(pc_wr_sel[1]), .Y(
        oc8051_memory_interface1_n613) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u623 ( .A0(
        oc8051_memory_interface1_n668), .A1(des2[7]), .B0(op2_n[7]), .B1(
        oc8051_memory_interface1_n613), .C0(des_acc[7]), .C1(
        oc8051_memory_interface1_n667), .Y(oc8051_memory_interface1_n702) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u622 ( .A(
        oc8051_memory_interface1_n702), .Y(oc8051_memory_interface1_n700) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u621 ( .A(
        oc8051_memory_interface1_n601), .B(oc8051_memory_interface1_n194), .Y(
        oc8051_memory_interface1_n600) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u620 ( .A(
        oc8051_memory_interface1_n600), .Y(oc8051_memory_interface1_n411) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u619 ( .A0(
        oc8051_memory_interface1_pc_buf_15_), .A1(
        oc8051_memory_interface1_n686), .B0(oc8051_memory_interface1_n687), 
        .B1(oc8051_memory_interface1_n700), .C0(oc8051_memory_interface1_n411), 
        .C1(oc8051_memory_interface1_n701), .Y(oc8051_memory_interface1_n699)
         );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u618 ( .A0(pc[15]), .A1(
        oc8051_memory_interface1_n696), .B0(oc8051_memory_interface1_n698), 
        .C0(oc8051_memory_interface1_n699), .Y(oc8051_memory_interface1_n459)
         );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u617 ( .A(
        oc8051_memory_interface1_n392), .B(oc8051_memory_interface1_n697), .Y(
        oc8051_memory_interface1_n688) );
  OAI31_X0P5M_A12TS oc8051_memory_interface1_u616 ( .A0(
        oc8051_memory_interface1_n695), .A1(oc8051_memory_interface1_n392), 
        .A2(oc8051_memory_interface1_n665), .B0(oc8051_memory_interface1_n696), 
        .Y(oc8051_memory_interface1_n694) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u615 ( .A(
        oc8051_memory_interface1_n694), .Y(oc8051_memory_interface1_n689) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u614 ( .A0(
        oc8051_memory_interface1_n668), .A1(des2[6]), .B0(op2_n[6]), .B1(
        oc8051_memory_interface1_n613), .C0(des_acc[6]), .C1(
        oc8051_memory_interface1_n667), .Y(oc8051_memory_interface1_n693) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u613 ( .A(
        oc8051_memory_interface1_n693), .Y(oc8051_memory_interface1_n691) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u612 ( .A0(
        oc8051_memory_interface1_pc_buf_14_), .A1(
        oc8051_memory_interface1_n686), .B0(oc8051_memory_interface1_n687), 
        .B1(oc8051_memory_interface1_n691), .C0(oc8051_memory_interface1_n411), 
        .C1(oc8051_memory_interface1_n692), .Y(oc8051_memory_interface1_n690)
         );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u611 ( .A0(
        oc8051_memory_interface1_n688), .A1(oc8051_memory_interface1_n673), 
        .B0(oc8051_memory_interface1_n689), .C0(oc8051_memory_interface1_n690), 
        .Y(oc8051_memory_interface1_n460) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u610 ( .A0(
        oc8051_memory_interface1_n667), .A1(des_acc[5]), .B0(
        oc8051_memory_interface1_n613), .B1(op2_n[5]), .C0(des2[5]), .C1(
        oc8051_memory_interface1_n668), .Y(oc8051_memory_interface1_n679) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u609 ( .A(
        oc8051_memory_interface1_n687), .Y(oc8051_memory_interface1_n657) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u608 ( .A(
        oc8051_memory_interface1_n686), .Y(oc8051_memory_interface1_n658) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u607 ( .A(
        oc8051_memory_interface1_n685), .B(oc8051_memory_interface1_n393), .Y(
        oc8051_memory_interface1_n682) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u606 ( .A0(
        oc8051_memory_interface1_n393), .A1(oc8051_memory_interface1_n676), 
        .B0(oc8051_memory_interface1_n684), .C0(oc8051_memory_interface1_n665), 
        .Y(oc8051_memory_interface1_n683) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u605 ( .A0(
        oc8051_memory_interface1_n411), .A1(oc8051_memory_interface1_n681), 
        .B0(oc8051_memory_interface1_n661), .B1(oc8051_memory_interface1_n682), 
        .C0(oc8051_memory_interface1_n683), .Y(oc8051_memory_interface1_n680)
         );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u604 ( .A0(
        oc8051_memory_interface1_n679), .A1(oc8051_memory_interface1_n657), 
        .B0(oc8051_memory_interface1_n658), .B1(oc8051_memory_interface1_n307), 
        .C0(oc8051_memory_interface1_n680), .Y(oc8051_memory_interface1_n461)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u603 ( .A0(
        oc8051_memory_interface1_n668), .A1(des2[4]), .B0(op2_n[4]), .B1(
        oc8051_memory_interface1_n613), .C0(des_acc[4]), .C1(
        oc8051_memory_interface1_n667), .Y(oc8051_memory_interface1_n672) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u602 ( .A(
        oc8051_memory_interface1_n678), .B(oc8051_memory_interface1_n394), .Y(
        oc8051_memory_interface1_n674) );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u601 ( .A0(pc[12]), .A1(
        oc8051_memory_interface1_n664), .B0(oc8051_memory_interface1_n676), 
        .C0(oc8051_memory_interface1_n677), .Y(oc8051_memory_interface1_n675)
         );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u600 ( .A0(
        oc8051_memory_interface1_n657), .A1(oc8051_memory_interface1_n672), 
        .B0(oc8051_memory_interface1_n673), .B1(oc8051_memory_interface1_n674), 
        .C0(oc8051_memory_interface1_n675), .Y(oc8051_memory_interface1_n671)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u599 ( .A(
        oc8051_memory_interface1_n671), .Y(oc8051_memory_interface1_n670) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u598 ( .A0(
        oc8051_memory_interface1_n669), .A1(oc8051_memory_interface1_n600), 
        .B0(oc8051_memory_interface1_n658), .B1(oc8051_memory_interface1_n302), 
        .C0(oc8051_memory_interface1_n670), .Y(oc8051_memory_interface1_n462)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u597 ( .A0(
        oc8051_memory_interface1_n667), .A1(des_acc[3]), .B0(
        oc8051_memory_interface1_n613), .B1(op2_n[3]), .C0(des2[3]), .C1(
        oc8051_memory_interface1_n668), .Y(oc8051_memory_interface1_n656) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u596 ( .A(
        oc8051_memory_interface1_n666), .B(oc8051_memory_interface1_n395), .Y(
        oc8051_memory_interface1_n662) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u595 ( .A0(
        oc8051_memory_interface1_n395), .A1(oc8051_memory_interface1_n650), 
        .B0(oc8051_memory_interface1_n664), .C0(oc8051_memory_interface1_n665), 
        .Y(oc8051_memory_interface1_n663) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u594 ( .A0(
        oc8051_memory_interface1_n411), .A1(oc8051_memory_interface1_n660), 
        .B0(oc8051_memory_interface1_n661), .B1(oc8051_memory_interface1_n662), 
        .C0(oc8051_memory_interface1_n663), .Y(oc8051_memory_interface1_n659)
         );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u593 ( .A0(
        oc8051_memory_interface1_n656), .A1(oc8051_memory_interface1_n657), 
        .B0(oc8051_memory_interface1_n658), .B1(oc8051_memory_interface1_n297), 
        .C0(oc8051_memory_interface1_n659), .Y(oc8051_memory_interface1_n463)
         );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u592 ( .A0(
        oc8051_memory_interface1_n652), .A1(oc8051_memory_interface1_n601), 
        .B0(oc8051_memory_interface1_n655), .C0(oc8051_memory_interface1_n613), 
        .Y(oc8051_memory_interface1_n654) );
  OA21_X0P5M_A12TS oc8051_memory_interface1_u591 ( .A0(pc_wr_sel[0]), .A1(
        oc8051_memory_interface1_n653), .B0(oc8051_memory_interface1_n654), 
        .Y(oc8051_memory_interface1_n617) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u590 ( .AN(
        oc8051_memory_interface1_n604), .B(oc8051_memory_interface1_n617), .Y(
        oc8051_memory_interface1_n616) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u589 ( .A(
        oc8051_memory_interface1_cdone), .B(oc8051_memory_interface1_dack_ir), 
        .Y(oc8051_memory_interface1_n388) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u588 ( .AN(
        oc8051_memory_interface1_n388), .B(oc8051_memory_interface1_n387), .Y(
        oc8051_memory_interface1_n383) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u587 ( .AN(
        oc8051_memory_interface1_cdone), .B(oc8051_memory_interface1_dack_ir), 
        .Y(oc8051_memory_interface1_n384) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u586 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_7_), .B0(
        oc8051_memory_interface1_n383), .B1(oc8051_memory_interface1_op1_7_), 
        .C0(oc8051_memory_interface1_cdata_7_), .C1(
        oc8051_memory_interface1_n384), .Y(oc8051_memory_interface1_n353) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u585 ( .A(
        oc8051_memory_interface1_n353), .Y(op1_n[7]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u584 ( .A(des2[2]), .Y(
        oc8051_memory_interface1_n645) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u583 ( .A(
        oc8051_memory_interface1_n603), .B(oc8051_memory_interface1_n652), .Y(
        oc8051_memory_interface1_n626) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u582 ( .A(
        oc8051_memory_interface1_n651), .B(pc[10]), .Y(
        oc8051_memory_interface1_n648) );
  AO21_X0P5M_A12TS oc8051_memory_interface1_u581 ( .A0(pc[10]), .A1(
        oc8051_memory_interface1_n639), .B0(oc8051_memory_interface1_n650), 
        .Y(oc8051_memory_interface1_n649) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u580 ( .A0(
        oc8051_memory_interface1_n626), .A1(op2_n[2]), .B0(
        oc8051_memory_interface1_n607), .B1(oc8051_memory_interface1_n648), 
        .C0(oc8051_memory_interface1_n608), .C1(oc8051_memory_interface1_n649), 
        .Y(oc8051_memory_interface1_n647) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u579 ( .A0(
        oc8051_memory_interface1_n615), .A1(oc8051_memory_interface1_n645), 
        .B0(oc8051_memory_interface1_n646), .B1(oc8051_memory_interface1_n614), 
        .C0(oc8051_memory_interface1_n647), .Y(oc8051_memory_interface1_n644)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u578 ( .A0(
        oc8051_memory_interface1_n411), .A1(oc8051_memory_interface1_n643), 
        .B0(oc8051_memory_interface1_n621), .B1(op1_n[7]), .C0(n_3_net_), .C1(
        oc8051_memory_interface1_n644), .Y(oc8051_memory_interface1_n642) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u577 ( .A0(
        oc8051_memory_interface1_n616), .A1(oc8051_memory_interface1_n292), 
        .B0(oc8051_memory_interface1_n617), .B1(oc8051_memory_interface1_n642), 
        .Y(oc8051_memory_interface1_n464) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u576 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_6_), .B0(
        oc8051_memory_interface1_n383), .B1(oc8051_memory_interface1_op1_6_), 
        .C0(oc8051_memory_interface1_cdata_6_), .C1(
        oc8051_memory_interface1_n384), .Y(oc8051_memory_interface1_n341) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u575 ( .A(
        oc8051_memory_interface1_n341), .Y(op1_n[6]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u574 ( .A(des2[1]), .Y(
        oc8051_memory_interface1_n634) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u573 ( .A(
        oc8051_memory_interface1_n641), .Y(op2_n[1]) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u572 ( .A(
        oc8051_memory_interface1_n640), .B(oc8051_memory_interface1_n397), .Y(
        oc8051_memory_interface1_n637) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u571 ( .A0(
        oc8051_memory_interface1_n397), .A1(oc8051_memory_interface1_n625), 
        .B0(oc8051_memory_interface1_n639), .Y(oc8051_memory_interface1_n638)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u570 ( .A0(
        oc8051_memory_interface1_n626), .A1(op2_n[1]), .B0(
        oc8051_memory_interface1_n607), .B1(oc8051_memory_interface1_n637), 
        .C0(oc8051_memory_interface1_n608), .C1(oc8051_memory_interface1_n638), 
        .Y(oc8051_memory_interface1_n636) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u569 ( .A0(
        oc8051_memory_interface1_n615), .A1(oc8051_memory_interface1_n634), 
        .B0(oc8051_memory_interface1_n635), .B1(oc8051_memory_interface1_n614), 
        .C0(oc8051_memory_interface1_n636), .Y(oc8051_memory_interface1_n633)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u568 ( .A0(
        oc8051_memory_interface1_n411), .A1(oc8051_memory_interface1_n632), 
        .B0(oc8051_memory_interface1_n621), .B1(op1_n[6]), .C0(n_3_net_), .C1(
        oc8051_memory_interface1_n633), .Y(oc8051_memory_interface1_n631) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u567 ( .A0(
        oc8051_memory_interface1_n616), .A1(oc8051_memory_interface1_n287), 
        .B0(oc8051_memory_interface1_n617), .B1(oc8051_memory_interface1_n631), 
        .Y(oc8051_memory_interface1_n465) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u566 ( .A(
        oc8051_memory_interface1_pc_buf_8_), .Y(oc8051_memory_interface1_n281)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u565 ( .A(des2[0]), .Y(
        oc8051_memory_interface1_n622) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u564 ( .A0(
        oc8051_memory_interface1_n398), .A1(oc8051_memory_interface1_n628), 
        .B0(oc8051_memory_interface1_n629), .C0(oc8051_memory_interface1_n630), 
        .Y(oc8051_memory_interface1_n627) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u563 ( .A0(
        oc8051_memory_interface1_n625), .A1(oc8051_memory_interface1_n608), 
        .B0(oc8051_memory_interface1_n626), .B1(op2_n[0]), .C0(
        oc8051_memory_interface1_n627), .Y(oc8051_memory_interface1_n624) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u562 ( .A0(
        oc8051_memory_interface1_n615), .A1(oc8051_memory_interface1_n622), 
        .B0(oc8051_memory_interface1_n623), .B1(oc8051_memory_interface1_n614), 
        .C0(oc8051_memory_interface1_n624), .Y(oc8051_memory_interface1_n620)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u561 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_5_), .B0(
        oc8051_memory_interface1_n383), .B1(oc8051_memory_interface1_op1_5_), 
        .C0(oc8051_memory_interface1_cdata_5_), .C1(
        oc8051_memory_interface1_n384), .Y(oc8051_memory_interface1_n349) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u560 ( .A(
        oc8051_memory_interface1_n349), .Y(op1_n[5]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u559 ( .A0(
        oc8051_memory_interface1_n411), .A1(oc8051_memory_interface1_n619), 
        .B0(n_3_net_), .B1(oc8051_memory_interface1_n620), .C0(
        oc8051_memory_interface1_n621), .C1(op1_n[5]), .Y(
        oc8051_memory_interface1_n618) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u558 ( .A0(
        oc8051_memory_interface1_n616), .A1(oc8051_memory_interface1_n281), 
        .B0(oc8051_memory_interface1_n617), .B1(oc8051_memory_interface1_n618), 
        .Y(oc8051_memory_interface1_n466) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u557 ( .A(
        oc8051_memory_interface1_n614), .B(oc8051_memory_interface1_n615), .Y(
        oc8051_memory_interface1_n405) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u556 ( .AN(
        oc8051_memory_interface1_n613), .B(pc_wr_sel[0]), .Y(
        oc8051_memory_interface1_n407) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u555 ( .A(
        oc8051_memory_interface1_n603), .B(pc_wr_sel[1]), .Y(
        oc8051_memory_interface1_n406) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u554 ( .A0(op2_n[7]), .A1(
        oc8051_memory_interface1_n407), .B0(oc8051_memory_interface1_n406), 
        .B1(op3_n[7]), .Y(oc8051_memory_interface1_n605) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u553 ( .A0(
        oc8051_memory_interface1_n612), .A1(oc8051_memory_interface1_n595), 
        .B0(oc8051_memory_interface1_n269), .Y(oc8051_memory_interface1_n611)
         );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u552 ( .A0(
        oc8051_memory_interface1_n596), .A1(oc8051_memory_interface1_n610), 
        .B0(oc8051_memory_interface1_n611), .Y(oc8051_memory_interface1_n609)
         );
  MXT4_X0P5M_A12TS oc8051_memory_interface1_u551 ( .A(
        oc8051_memory_interface1_n607), .B(oc8051_memory_interface1_n608), .C(
        oc8051_memory_interface1_n608), .D(oc8051_memory_interface1_n607), 
        .S0(pc[7]), .S1(oc8051_memory_interface1_n609), .Y(
        oc8051_memory_interface1_n606) );
  AOI211_X0P5M_A12TS oc8051_memory_interface1_u550 ( .A0(des_acc[7]), .A1(
        oc8051_memory_interface1_n405), .B0(oc8051_memory_interface1_n605), 
        .C0(oc8051_memory_interface1_n606), .Y(oc8051_memory_interface1_n598)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u549 ( .A(
        oc8051_memory_interface1_n405), .Y(oc8051_memory_interface1_n602) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u548 ( .A0(
        oc8051_memory_interface1_n602), .A1(oc8051_memory_interface1_n603), 
        .B0(n_3_net_), .Y(oc8051_memory_interface1_n400) );
  OAI31_X0P5M_A12TS oc8051_memory_interface1_u547 ( .A0(
        oc8051_memory_interface1_n601), .A1(oc8051_memory_interface1_n602), 
        .A2(oc8051_memory_interface1_n603), .B0(oc8051_memory_interface1_n604), 
        .Y(oc8051_memory_interface1_n410) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u546 ( .A(
        oc8051_memory_interface1_n410), .Y(oc8051_memory_interface1_n554) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u545 ( .A0(
        oc8051_memory_interface1_n598), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n599), .B1(oc8051_memory_interface1_n600), 
        .C0(oc8051_memory_interface1_n554), .C1(oc8051_memory_interface1_n277), 
        .Y(oc8051_memory_interface1_n467) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u544 ( .A0(des_acc[6]), .A1(
        oc8051_memory_interface1_n405), .B0(op3_n[6]), .B1(
        oc8051_memory_interface1_n406), .C0(oc8051_memory_interface1_n407), 
        .C1(op2_n[6]), .Y(oc8051_memory_interface1_n591) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u543 ( .A(
        oc8051_memory_interface1_n400), .Y(oc8051_memory_interface1_n585) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u542 ( .A(
        oc8051_memory_interface1_n597), .B(oc8051_memory_interface1_n585), .Y(
        oc8051_memory_interface1_n402) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u541 ( .A(
        oc8051_memory_interface1_n595), .B(oc8051_memory_interface1_n596), .C(
        oc8051_memory_interface1_n269), .Y(oc8051_memory_interface1_n592) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u540 ( .A0(
        oc8051_memory_interface1_pc_buf_6_), .A1(oc8051_memory_interface1_n410), .B0(oc8051_memory_interface1_n411), .B1(oc8051_memory_interface1_n594), .Y(
        oc8051_memory_interface1_n593) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u539 ( .A0(
        oc8051_memory_interface1_n591), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n402), .B1(oc8051_memory_interface1_n592), 
        .C0(oc8051_memory_interface1_n593), .Y(oc8051_memory_interface1_n468)
         );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u538 ( .A(
        oc8051_memory_interface1_n589), .B(pc[5]), .C(
        oc8051_memory_interface1_n590), .Y(oc8051_memory_interface1_n552) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u537 ( .A0(op2_n[5]), .A1(
        oc8051_memory_interface1_n407), .B0(oc8051_memory_interface1_n406), 
        .B1(op3_n[5]), .C0(oc8051_memory_interface1_n405), .C1(des_acc[5]), 
        .Y(oc8051_memory_interface1_n588) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u536 ( .A(
        oc8051_memory_interface1_n588), .Y(oc8051_memory_interface1_n586) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u535 ( .A0(
        oc8051_memory_interface1_n585), .A1(oc8051_memory_interface1_n586), 
        .B0(oc8051_memory_interface1_n411), .B1(oc8051_memory_interface1_n587), 
        .Y(oc8051_memory_interface1_n556) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u534 ( .A0(
        oc8051_memory_interface1_n402), .A1(oc8051_memory_interface1_n552), 
        .B0(oc8051_memory_interface1_n554), .B1(oc8051_memory_interface1_n265), 
        .C0(oc8051_memory_interface1_n556), .Y(oc8051_memory_interface1_n469)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u533 ( .A0(des_acc[4]), .A1(
        oc8051_memory_interface1_n405), .B0(op3_n[4]), .B1(
        oc8051_memory_interface1_n406), .C0(oc8051_memory_interface1_n407), 
        .C1(op2_n[4]), .Y(oc8051_memory_interface1_n458) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u532 ( .A(pc[4]), .Y(
        oc8051_memory_interface1_n257) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u531 ( .A(
        oc8051_memory_interface1_n548), .B(oc8051_memory_interface1_n257), .C(
        oc8051_memory_interface1_n550), .Y(oc8051_memory_interface1_n542) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u530 ( .A0(
        oc8051_memory_interface1_pc_buf_4_), .A1(oc8051_memory_interface1_n410), .B0(oc8051_memory_interface1_n411), .B1(oc8051_memory_interface1_n546), .Y(
        oc8051_memory_interface1_n544) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u529 ( .A0(
        oc8051_memory_interface1_n458), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n402), .B1(oc8051_memory_interface1_n542), 
        .C0(oc8051_memory_interface1_n544), .Y(oc8051_memory_interface1_n470)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u528 ( .A0(des_acc[3]), .A1(
        oc8051_memory_interface1_n405), .B0(op3_n[3]), .B1(
        oc8051_memory_interface1_n406), .C0(oc8051_memory_interface1_n407), 
        .C1(op2_n[3]), .Y(oc8051_memory_interface1_n436) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u527 ( .A(
        oc8051_memory_interface1_n456), .B(oc8051_memory_interface1_n457), .C(
        pc[3]), .Y(oc8051_memory_interface1_n437) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u526 ( .A0(
        oc8051_memory_interface1_n411), .A1(oc8051_memory_interface1_n439), 
        .B0(oc8051_memory_interface1_pc_buf_3_), .B1(
        oc8051_memory_interface1_n410), .Y(oc8051_memory_interface1_n438) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u525 ( .A0(
        oc8051_memory_interface1_n436), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n402), .B1(oc8051_memory_interface1_n437), 
        .C0(oc8051_memory_interface1_n438), .Y(oc8051_memory_interface1_n471)
         );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u524 ( .A0(des_acc[2]), .A1(
        oc8051_memory_interface1_n405), .B0(op3_n[2]), .B1(
        oc8051_memory_interface1_n406), .C0(oc8051_memory_interface1_n407), 
        .C1(op2_n[2]), .Y(oc8051_memory_interface1_n415) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u523 ( .A(
        oc8051_memory_interface1_n434), .B(oc8051_memory_interface1_n435), .C(
        pc[2]), .Y(oc8051_memory_interface1_n432) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u522 ( .A(
        oc8051_memory_interface1_n411), .B(oc8051_memory_interface1_n410), 
        .S0(oc8051_memory_interface1_pc_buf_2_), .Y(
        oc8051_memory_interface1_n433) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u521 ( .A0(
        oc8051_memory_interface1_n415), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n402), .B1(oc8051_memory_interface1_n432), 
        .C0(oc8051_memory_interface1_n433), .Y(oc8051_memory_interface1_n472)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u520 ( .A(pc[1]), .Y(
        oc8051_memory_interface1_n241) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u519 ( .A(
        oc8051_memory_interface1_n414), .Y(op3_n[1]) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u518 ( .A(op2_n[1]), .B(op3_n[1]), 
        .S0(pc_wr_sel[0]), .Y(oc8051_memory_interface1_n413) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u517 ( .A(
        oc8051_memory_interface1_n412), .B(oc8051_memory_interface1_n241), .C(
        oc8051_memory_interface1_n413), .Y(oc8051_memory_interface1_n408) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u516 ( .A0(des_acc[1]), .A1(
        oc8051_memory_interface1_n405), .B0(op3_n[1]), .B1(
        oc8051_memory_interface1_n406), .C0(oc8051_memory_interface1_n407), 
        .C1(op2_n[1]), .Y(oc8051_memory_interface1_n409) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u515 ( .A(
        oc8051_memory_interface1_n410), .B(oc8051_memory_interface1_n411), .Y(
        oc8051_memory_interface1_n403) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u514 ( .A0(
        oc8051_memory_interface1_n408), .A1(oc8051_memory_interface1_n402), 
        .B0(oc8051_memory_interface1_n409), .B1(oc8051_memory_interface1_n400), 
        .C0(oc8051_memory_interface1_n403), .C1(oc8051_memory_interface1_n243), 
        .Y(oc8051_memory_interface1_n473) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u513 ( .A0(des_acc[0]), .A1(
        oc8051_memory_interface1_n405), .B0(oc8051_memory_interface1_n406), 
        .B1(op3_n[0]), .C0(oc8051_memory_interface1_n407), .C1(op2_n[0]), .Y(
        oc8051_memory_interface1_n391) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u512 ( .A(
        oc8051_memory_interface1_n404), .B(pc[0]), .Y(
        oc8051_memory_interface1_n401) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u511 ( .A0(
        oc8051_memory_interface1_n391), .A1(oc8051_memory_interface1_n400), 
        .B0(oc8051_memory_interface1_n401), .B1(oc8051_memory_interface1_n402), 
        .C0(oc8051_memory_interface1_n403), .C1(oc8051_memory_interface1_n239), 
        .Y(oc8051_memory_interface1_n474) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u510 ( .A(
        oc8051_memory_interface1_n185), .B(oc8051_memory_interface1_n197), .C(
        rd), .Y(oc8051_memory_interface1_n237) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u509 ( .A(
        oc8051_memory_interface1_n237), .B(oc8051_memory_interface1_n197), .Y(
        oc8051_memory_interface1_n235) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u508 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_3_), .B0(
        oc8051_memory_interface1_n383), .B1(oc8051_memory_interface1_op1_3_), 
        .C0(oc8051_memory_interface1_cdata_3_), .C1(
        oc8051_memory_interface1_n384), .Y(oc8051_memory_interface1_n343) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u507 ( .A0(
        oc8051_memory_interface1_ddat_ir_1_), .A1(
        oc8051_memory_interface1_dack_ir), .B0(oc8051_memory_interface1_n384), 
        .B1(oc8051_memory_interface1_cdata_1_), .Y(
        oc8051_memory_interface1_n390) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u506 ( .A0(
        oc8051_memory_interface1_n387), .A1(oc8051_memory_interface1_op1_1_), 
        .B0(oc8051_memory_interface1_n388), .C0(oc8051_memory_interface1_n390), 
        .Y(oc8051_memory_interface1_n346) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u505 ( .A0(
        oc8051_memory_interface1_ddat_ir_4_), .A1(
        oc8051_memory_interface1_dack_ir), .B0(oc8051_memory_interface1_n384), 
        .B1(oc8051_memory_interface1_cdata_4_), .Y(
        oc8051_memory_interface1_n389) );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u504 ( .A0(
        oc8051_memory_interface1_n387), .A1(oc8051_memory_interface1_op1_4_), 
        .B0(oc8051_memory_interface1_n388), .C0(oc8051_memory_interface1_n389), 
        .Y(oc8051_memory_interface1_n344) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u503 ( .A(op1_n[7]), .B(
        oc8051_memory_interface1_n341), .Y(oc8051_memory_interface1_n381) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u502 ( .A0(op1_n[6]), .A1(
        op1_n[5]), .B0(oc8051_memory_interface1_n353), .Y(
        oc8051_memory_interface1_n385) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u501 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_0_), .B0(
        oc8051_memory_interface1_n383), .B1(oc8051_memory_interface1_op1_0_), 
        .C0(oc8051_memory_interface1_cdata_0_), .C1(
        oc8051_memory_interface1_n384), .Y(oc8051_memory_interface1_n359) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u500 ( .A(
        oc8051_memory_interface1_n359), .Y(op1_n[0]) );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u499 ( .A0(op1_n[6]), .A1(
        oc8051_memory_interface1_n349), .B0(op1_n[0]), .Y(
        oc8051_memory_interface1_n386) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u498 ( .A0(
        oc8051_memory_interface1_n344), .A1(oc8051_memory_interface1_n381), 
        .B0(oc8051_memory_interface1_n385), .C0(oc8051_memory_interface1_n386), 
        .Y(oc8051_memory_interface1_n377) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u497 ( .A0(
        oc8051_memory_interface1_dack_ir), .A1(
        oc8051_memory_interface1_ddat_ir_2_), .B0(
        oc8051_memory_interface1_n383), .B1(oc8051_memory_interface1_op1_2_), 
        .C0(oc8051_memory_interface1_cdata_2_), .C1(
        oc8051_memory_interface1_n384), .Y(oc8051_memory_interface1_n345) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u496 ( .A(
        oc8051_memory_interface1_n345), .Y(op1_n[2]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u495 ( .A(
        oc8051_memory_interface1_n343), .Y(op1_n[3]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u494 ( .A(op1_n[2]), .B(op1_n[3]), 
        .Y(oc8051_memory_interface1_n355) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u493 ( .A(
        oc8051_memory_interface1_n346), .Y(op1_n[1]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u492 ( .A(
        oc8051_memory_interface1_n344), .Y(op1_n[4]) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u491 ( .A(op1_n[6]), .B(op1_n[1]), 
        .C(op1_n[4]), .Y(oc8051_memory_interface1_n368) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u490 ( .A(
        oc8051_memory_interface1_n359), .B(oc8051_memory_interface1_n349), .Y(
        oc8051_memory_interface1_n361) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u489 ( .A(op1_n[4]), .B(op1_n[5]), 
        .C(op1_n[0]), .Y(oc8051_memory_interface1_n382) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u488 ( .A(op1_n[6]), .B(
        oc8051_memory_interface1_n353), .C(oc8051_memory_interface1_n382), .Y(
        oc8051_memory_interface1_n379) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u487 ( .A(
        oc8051_memory_interface1_n381), .Y(oc8051_memory_interface1_n372) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u486 ( .A(
        oc8051_memory_interface1_n346), .B(oc8051_memory_interface1_n372), 
        .S0(oc8051_memory_interface1_n359), .Y(oc8051_memory_interface1_n380)
         );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u485 ( .A0(
        oc8051_memory_interface1_n368), .A1(oc8051_memory_interface1_n361), 
        .B0(oc8051_memory_interface1_n379), .C0(oc8051_memory_interface1_n380), 
        .Y(oc8051_memory_interface1_n378) );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u484 ( .A0(
        oc8051_memory_interface1_n343), .A1(oc8051_memory_interface1_n346), 
        .A2(oc8051_memory_interface1_n377), .B0(oc8051_memory_interface1_n355), 
        .B1(oc8051_memory_interface1_n378), .Y(oc8051_memory_interface1_n370)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u483 ( .A0(
        oc8051_memory_interface1_n346), .A1(oc8051_memory_interface1_n345), 
        .B0(oc8051_memory_interface1_n343), .Y(oc8051_memory_interface1_n362)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u482 ( .A(op1_n[4]), .B(
        oc8051_memory_interface1_n349), .Y(oc8051_memory_interface1_n369) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u481 ( .A(
        oc8051_memory_interface1_n341), .B(oc8051_memory_interface1_n344), .Y(
        oc8051_memory_interface1_n373) );
  OR2_X0P5M_A12TS oc8051_memory_interface1_u480 ( .A(
        oc8051_memory_interface1_n355), .B(op1_n[7]), .Y(
        oc8051_memory_interface1_n375) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u479 ( .A(op1_n[3]), .B(op1_n[7]), 
        .Y(oc8051_memory_interface1_n376) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u478 ( .A(
        oc8051_memory_interface1_n375), .B(oc8051_memory_interface1_n376), 
        .S0(oc8051_memory_interface1_n349), .Y(oc8051_memory_interface1_n374)
         );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u477 ( .A0(
        oc8051_memory_interface1_n362), .A1(oc8051_memory_interface1_n369), 
        .A2(oc8051_memory_interface1_n372), .B0(oc8051_memory_interface1_n373), 
        .B1(oc8051_memory_interface1_n374), .Y(oc8051_memory_interface1_n371)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u476 ( .A(
        oc8051_memory_interface1_n370), .B(oc8051_memory_interface1_n371), .Y(
        oc8051_memory_interface1_n245) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u475 ( .A(
        oc8051_memory_interface1_n245), .Y(oc8051_memory_interface1_n195) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u474 ( .A(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n188)
         );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u473 ( .A(
        oc8051_memory_interface1_n239), .B(oc8051_memory_interface1_n188), .Y(
        oc8051_memory_interface1_n240) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u472 ( .A(
        oc8051_memory_interface1_n369), .Y(oc8051_memory_interface1_n367) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u471 ( .A0(op1_n[4]), .A1(
        op1_n[1]), .B0(oc8051_memory_interface1_n367), .B1(op1_n[6]), .C0(
        oc8051_memory_interface1_n368), .Y(oc8051_memory_interface1_n363) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u470 ( .A(
        oc8051_memory_interface1_n349), .B(op1_n[6]), .Y(
        oc8051_memory_interface1_n365) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u469 ( .A(
        oc8051_memory_interface1_n341), .B(op1_n[0]), .Y(
        oc8051_memory_interface1_n366) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u468 ( .A(
        oc8051_memory_interface1_n365), .B(oc8051_memory_interface1_n366), 
        .S0(oc8051_memory_interface1_n344), .Y(oc8051_memory_interface1_n364)
         );
  OA21A1OI2_X0P5M_A12TS oc8051_memory_interface1_u467 ( .A0(op1_n[3]), .A1(
        oc8051_memory_interface1_n363), .B0(oc8051_memory_interface1_n364), 
        .C0(oc8051_memory_interface1_n345), .Y(oc8051_memory_interface1_n356)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u466 ( .A(
        oc8051_memory_interface1_n362), .Y(oc8051_memory_interface1_n348) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u465 ( .A(
        oc8051_memory_interface1_n343), .B(oc8051_memory_interface1_n346), .Y(
        oc8051_memory_interface1_n360) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u464 ( .A(
        oc8051_memory_interface1_n361), .Y(oc8051_memory_interface1_n347) );
  AOI211_X0P5M_A12TS oc8051_memory_interface1_u463 ( .A0(
        oc8051_memory_interface1_n345), .A1(oc8051_memory_interface1_n359), 
        .B0(oc8051_memory_interface1_n360), .C0(oc8051_memory_interface1_n347), 
        .Y(oc8051_memory_interface1_n358) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u462 ( .A0(op1_n[5]), .A1(
        oc8051_memory_interface1_n348), .B0(op1_n[6]), .B1(
        oc8051_memory_interface1_n358), .Y(oc8051_memory_interface1_n357) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u461 ( .A(
        oc8051_memory_interface1_n356), .B(oc8051_memory_interface1_n357), 
        .S0(oc8051_memory_interface1_n353), .Y(oc8051_memory_interface1_n336)
         );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u460 ( .A(op1_n[0]), .B(op1_n[1]), 
        .C(oc8051_memory_interface1_n355), .Y(oc8051_memory_interface1_n337)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u459 ( .A(op1_n[0]), .B(
        oc8051_memory_interface1_n343), .Y(oc8051_memory_interface1_n351) );
  NAND4B_X0P5M_A12TS oc8051_memory_interface1_u458 ( .AN(
        oc8051_memory_interface1_n351), .B(op1_n[2]), .C(op1_n[4]), .D(
        oc8051_memory_interface1_n346), .Y(oc8051_memory_interface1_n354) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u457 ( .A(
        oc8051_memory_interface1_n354), .Y(oc8051_memory_interface1_n352) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u456 ( .A(
        oc8051_memory_interface1_n351), .B(oc8051_memory_interface1_n352), 
        .S0(oc8051_memory_interface1_n353), .Y(oc8051_memory_interface1_n350)
         );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u455 ( .A0(op1_n[4]), .A1(
        oc8051_memory_interface1_n348), .B0(oc8051_memory_interface1_n349), 
        .B1(oc8051_memory_interface1_n350), .Y(oc8051_memory_interface1_n339)
         );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u454 ( .A(
        oc8051_memory_interface1_n345), .B(oc8051_memory_interface1_n346), .C(
        oc8051_memory_interface1_n347), .Y(oc8051_memory_interface1_n342) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u453 ( .A0(
        oc8051_memory_interface1_n342), .A1(oc8051_memory_interface1_n343), 
        .B0(oc8051_memory_interface1_n344), .Y(oc8051_memory_interface1_n340)
         );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u452 ( .A(
        oc8051_memory_interface1_n339), .B(oc8051_memory_interface1_n340), 
        .S0(oc8051_memory_interface1_n341), .Y(oc8051_memory_interface1_n338)
         );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u451 ( .A(
        oc8051_memory_interface1_n336), .B(oc8051_memory_interface1_n337), .C(
        oc8051_memory_interface1_n338), .Y(oc8051_memory_interface1_n234) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u450 ( .A(
        oc8051_memory_interface1_n240), .B(oc8051_memory_interface1_n234), .Y(
        oc8051_memory_interface1_n244) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u449 ( .AN(
        oc8051_memory_interface1_n244), .B(oc8051_memory_interface1_n245), .Y(
        oc8051_memory_interface1_n334) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u448 ( .A(
        oc8051_memory_interface1_op_pos_1_), .Y(oc8051_memory_interface1_n196)
         );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u447 ( .A(
        oc8051_memory_interface1_pc_buf_0_), .B(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n335)
         );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u446 ( .A(
        oc8051_memory_interface1_pc_buf_1_), .B(oc8051_memory_interface1_n196), 
        .C(oc8051_memory_interface1_n335), .Y(oc8051_memory_interface1_n246)
         );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u445 ( .A0(
        oc8051_memory_interface1_n195), .A1(oc8051_memory_interface1_n244), 
        .B0(oc8051_memory_interface1_n334), .B1(oc8051_memory_interface1_n246), 
        .Y(oc8051_memory_interface1_n250) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u444 ( .A(
        oc8051_memory_interface1_n188), .B(oc8051_memory_interface1_n239), .Y(
        oc8051_memory_interface1_n333) );
  CGENI_X1M_A12TS oc8051_memory_interface1_u443 ( .A(
        oc8051_memory_interface1_op_pos_1_), .B(
        oc8051_memory_interface1_pc_buf_1_), .CI(oc8051_memory_interface1_n333), .CON(oc8051_memory_interface1_n331) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u442 ( .A(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n202)
         );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u441 ( .A(
        oc8051_memory_interface1_n331), .B(oc8051_memory_interface1_n249), .C(
        oc8051_memory_interface1_n202), .Y(oc8051_memory_interface1_n251) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u440 ( .AN(
        oc8051_memory_interface1_n331), .B(oc8051_memory_interface1_op_pos_2_), 
        .Y(oc8051_memory_interface1_n332) );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u439 ( .A0(
        oc8051_memory_interface1_n331), .A1(oc8051_memory_interface1_n202), 
        .B0(oc8051_memory_interface1_n332), .B1(oc8051_memory_interface1_n249), 
        .Y(oc8051_memory_interface1_n329) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u438 ( .A(
        oc8051_memory_interface1_n329), .B(oc8051_memory_interface1_n254), .Y(
        oc8051_memory_interface1_n255) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u437 ( .A0(
        oc8051_memory_interface1_n250), .A1(oc8051_memory_interface1_n251), 
        .B0(oc8051_memory_interface1_n255), .Y(oc8051_memory_interface1_n256)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u436 ( .A(
        oc8051_memory_interface1_n256), .Y(oc8051_memory_interface1_n261) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u435 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .B(oc8051_memory_interface1_n329), 
        .Y(oc8051_memory_interface1_n330) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u434 ( .A(
        oc8051_memory_interface1_n330), .B(oc8051_memory_interface1_pc_buf_4_), 
        .Y(oc8051_memory_interface1_n260) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u433 ( .A(
        oc8051_memory_interface1_n261), .B(oc8051_memory_interface1_n260), .Y(
        oc8051_memory_interface1_n262) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u432 ( .A(
        oc8051_memory_interface1_n262), .Y(oc8051_memory_interface1_n267) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u431 ( .A(
        oc8051_memory_interface1_pc_buf_3_), .B(oc8051_memory_interface1_n329), 
        .C(oc8051_memory_interface1_pc_buf_4_), .Y(
        oc8051_memory_interface1_n327) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u430 ( .A(
        oc8051_memory_interface1_n327), .B(oc8051_memory_interface1_n265), .Y(
        oc8051_memory_interface1_n266) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u429 ( .A(
        oc8051_memory_interface1_n267), .B(oc8051_memory_interface1_n266), .Y(
        oc8051_memory_interface1_n268) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u428 ( .A(
        oc8051_memory_interface1_n268), .Y(oc8051_memory_interface1_n273) );
  NAND2B_X0P5M_A12TS oc8051_memory_interface1_u427 ( .AN(
        oc8051_memory_interface1_n327), .B(oc8051_memory_interface1_pc_buf_5_), 
        .Y(oc8051_memory_interface1_n328) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u426 ( .A(
        oc8051_memory_interface1_n328), .B(oc8051_memory_interface1_pc_buf_6_), 
        .Y(oc8051_memory_interface1_n272) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u425 ( .A(
        oc8051_memory_interface1_n273), .B(oc8051_memory_interface1_n272), .Y(
        oc8051_memory_interface1_n274) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u424 ( .A(
        oc8051_memory_interface1_n274), .Y(oc8051_memory_interface1_n279) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u423 ( .A(
        oc8051_memory_interface1_n327), .B(oc8051_memory_interface1_n265), .C(
        oc8051_memory_interface1_n271), .Y(oc8051_memory_interface1_n325) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u422 ( .A(
        oc8051_memory_interface1_n325), .B(oc8051_memory_interface1_pc_buf_7_), 
        .Y(oc8051_memory_interface1_n278) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u421 ( .A(
        oc8051_memory_interface1_n279), .B(oc8051_memory_interface1_n278), .Y(
        oc8051_memory_interface1_n280) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u420 ( .A(
        oc8051_memory_interface1_n280), .Y(oc8051_memory_interface1_n284) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u419 ( .A(
        oc8051_memory_interface1_n325), .B(oc8051_memory_interface1_pc_buf_7_), 
        .Y(oc8051_memory_interface1_n326) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u418 ( .A(
        oc8051_memory_interface1_n326), .B(oc8051_memory_interface1_pc_buf_8_), 
        .Y(oc8051_memory_interface1_n283) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u417 ( .A(
        oc8051_memory_interface1_n284), .B(oc8051_memory_interface1_n283), .Y(
        oc8051_memory_interface1_n285) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u416 ( .A(
        oc8051_memory_interface1_n285), .Y(oc8051_memory_interface1_n290) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u415 ( .A(
        oc8051_memory_interface1_n325), .B(oc8051_memory_interface1_pc_buf_7_), 
        .C(oc8051_memory_interface1_pc_buf_8_), .Y(
        oc8051_memory_interface1_n323) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u414 ( .A(
        oc8051_memory_interface1_n323), .B(oc8051_memory_interface1_n287), .Y(
        oc8051_memory_interface1_n289) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u413 ( .A(
        oc8051_memory_interface1_n290), .B(oc8051_memory_interface1_n289), .Y(
        oc8051_memory_interface1_n291) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u412 ( .A(
        oc8051_memory_interface1_n291), .Y(oc8051_memory_interface1_n295) );
  NAND2B_X0P5M_A12TS oc8051_memory_interface1_u411 ( .AN(
        oc8051_memory_interface1_n323), .B(oc8051_memory_interface1_pc_buf_9_), 
        .Y(oc8051_memory_interface1_n324) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u410 ( .A(
        oc8051_memory_interface1_n324), .B(oc8051_memory_interface1_pc_buf_10_), .Y(oc8051_memory_interface1_n294) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u409 ( .A(
        oc8051_memory_interface1_n295), .B(oc8051_memory_interface1_n294), .Y(
        oc8051_memory_interface1_n296) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u408 ( .A(
        oc8051_memory_interface1_n296), .Y(oc8051_memory_interface1_n300) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u407 ( .A(
        oc8051_memory_interface1_n323), .B(oc8051_memory_interface1_n287), .C(
        oc8051_memory_interface1_n292), .Y(oc8051_memory_interface1_n321) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u406 ( .A(
        oc8051_memory_interface1_n321), .B(oc8051_memory_interface1_pc_buf_11_), .Y(oc8051_memory_interface1_n299) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u405 ( .A(
        oc8051_memory_interface1_n300), .B(oc8051_memory_interface1_n299), .Y(
        oc8051_memory_interface1_n301) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u404 ( .A(
        oc8051_memory_interface1_n301), .Y(oc8051_memory_interface1_n305) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u403 ( .A(
        oc8051_memory_interface1_n321), .B(oc8051_memory_interface1_pc_buf_11_), .Y(oc8051_memory_interface1_n322) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u402 ( .A(
        oc8051_memory_interface1_n322), .B(oc8051_memory_interface1_pc_buf_12_), .Y(oc8051_memory_interface1_n304) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u401 ( .A(
        oc8051_memory_interface1_n305), .B(oc8051_memory_interface1_n304), .Y(
        oc8051_memory_interface1_n306) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u400 ( .A(
        oc8051_memory_interface1_n306), .Y(oc8051_memory_interface1_n310) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u399 ( .A(
        oc8051_memory_interface1_n321), .B(oc8051_memory_interface1_pc_buf_11_), .C(oc8051_memory_interface1_pc_buf_12_), .Y(oc8051_memory_interface1_n320)
         );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u398 ( .A(
        oc8051_memory_interface1_n320), .B(oc8051_memory_interface1_n307), .Y(
        oc8051_memory_interface1_n309) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u397 ( .A(
        oc8051_memory_interface1_n310), .B(oc8051_memory_interface1_n309), .Y(
        oc8051_memory_interface1_n311) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u396 ( .A(
        oc8051_memory_interface1_n320), .B(oc8051_memory_interface1_n307), .Y(
        oc8051_memory_interface1_n319) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u395 ( .A(
        oc8051_memory_interface1_n319), .B(oc8051_memory_interface1_n313), .Y(
        oc8051_memory_interface1_n314) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u394 ( .AN(
        oc8051_memory_interface1_n311), .B(oc8051_memory_interface1_n314), .Y(
        oc8051_memory_interface1_n317) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u393 ( .A(
        oc8051_memory_interface1_pc_buf_15_), .Y(oc8051_memory_interface1_n316) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u392 ( .A(
        oc8051_memory_interface1_n319), .B(oc8051_memory_interface1_pc_buf_14_), .Y(oc8051_memory_interface1_n318) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u391 ( .A(
        oc8051_memory_interface1_n317), .B(oc8051_memory_interface1_n316), .C(
        oc8051_memory_interface1_n318), .Y(oc8051_memory_interface1_n315) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u390 ( .A0(
        oc8051_memory_interface1_n399), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n315), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n316), 
        .Y(oc8051_memory_interface1_n475) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u389 ( .A(
        oc8051_memory_interface1_n311), .B(oc8051_memory_interface1_n314), .Y(
        oc8051_memory_interface1_n312) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u388 ( .A0(
        oc8051_memory_interface1_n392), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n312), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n313), 
        .Y(oc8051_memory_interface1_n476) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u387 ( .A(
        oc8051_memory_interface1_n237), .Y(oc8051_memory_interface1_n286) );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u386 ( .A0(
        oc8051_memory_interface1_n309), .A1(oc8051_memory_interface1_n310), 
        .B0(oc8051_memory_interface1_n311), .C0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n308) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u385 ( .A0(
        oc8051_memory_interface1_n393), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n307), 
        .C0(oc8051_memory_interface1_n308), .Y(oc8051_memory_interface1_n477)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u384 ( .A0(
        oc8051_memory_interface1_n304), .A1(oc8051_memory_interface1_n305), 
        .B0(oc8051_memory_interface1_n306), .C0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n303) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u383 ( .A0(
        oc8051_memory_interface1_n394), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n302), 
        .C0(oc8051_memory_interface1_n303), .Y(oc8051_memory_interface1_n478)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u382 ( .A0(
        oc8051_memory_interface1_n299), .A1(oc8051_memory_interface1_n300), 
        .B0(oc8051_memory_interface1_n301), .C0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n298) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u381 ( .A0(
        oc8051_memory_interface1_n395), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n297), 
        .C0(oc8051_memory_interface1_n298), .Y(oc8051_memory_interface1_n479)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u380 ( .A0(
        oc8051_memory_interface1_n294), .A1(oc8051_memory_interface1_n295), 
        .B0(oc8051_memory_interface1_n296), .C0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n293) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u379 ( .A0(
        oc8051_memory_interface1_n396), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n292), 
        .C0(oc8051_memory_interface1_n293), .Y(oc8051_memory_interface1_n480)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u378 ( .A0(
        oc8051_memory_interface1_n289), .A1(oc8051_memory_interface1_n290), 
        .B0(oc8051_memory_interface1_n291), .C0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n288) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u377 ( .A0(
        oc8051_memory_interface1_n397), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n287), 
        .C0(oc8051_memory_interface1_n288), .Y(oc8051_memory_interface1_n481)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_memory_interface1_u376 ( .A0(
        oc8051_memory_interface1_n283), .A1(oc8051_memory_interface1_n284), 
        .B0(oc8051_memory_interface1_n285), .C0(oc8051_memory_interface1_n286), 
        .Y(oc8051_memory_interface1_n282) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u375 ( .A0(
        oc8051_memory_interface1_n398), .A1(oc8051_memory_interface1_n235), 
        .B0(oc8051_memory_interface1_n197), .B1(oc8051_memory_interface1_n281), 
        .C0(oc8051_memory_interface1_n282), .Y(oc8051_memory_interface1_n482)
         );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u374 ( .A0(
        oc8051_memory_interface1_n278), .A1(oc8051_memory_interface1_n279), 
        .B0(oc8051_memory_interface1_n280), .Y(oc8051_memory_interface1_n276)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u373 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n275), 
        .B0(oc8051_memory_interface1_n276), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n277), 
        .Y(oc8051_memory_interface1_n483) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u372 ( .A0(
        oc8051_memory_interface1_n272), .A1(oc8051_memory_interface1_n273), 
        .B0(oc8051_memory_interface1_n274), .Y(oc8051_memory_interface1_n270)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u371 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n269), 
        .B0(oc8051_memory_interface1_n270), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n271), 
        .Y(oc8051_memory_interface1_n484) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u370 ( .A0(
        oc8051_memory_interface1_n266), .A1(oc8051_memory_interface1_n267), 
        .B0(oc8051_memory_interface1_n268), .Y(oc8051_memory_interface1_n264)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u369 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n263), 
        .B0(oc8051_memory_interface1_n264), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n265), 
        .Y(oc8051_memory_interface1_n485) );
  AOI21_X0P5M_A12TS oc8051_memory_interface1_u368 ( .A0(
        oc8051_memory_interface1_n260), .A1(oc8051_memory_interface1_n261), 
        .B0(oc8051_memory_interface1_n262), .Y(oc8051_memory_interface1_n258)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u367 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n257), 
        .B0(oc8051_memory_interface1_n258), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n259), 
        .Y(oc8051_memory_interface1_n486) );
  AOI31_X0P5M_A12TS oc8051_memory_interface1_u366 ( .A0(
        oc8051_memory_interface1_n251), .A1(oc8051_memory_interface1_n250), 
        .A2(oc8051_memory_interface1_n255), .B0(oc8051_memory_interface1_n256), 
        .Y(oc8051_memory_interface1_n253) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u365 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n252), 
        .B0(oc8051_memory_interface1_n253), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n254), 
        .Y(oc8051_memory_interface1_n487) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u364 ( .A(
        oc8051_memory_interface1_n250), .B(oc8051_memory_interface1_n251), .Y(
        oc8051_memory_interface1_n248) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u363 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n247), 
        .B0(oc8051_memory_interface1_n248), .B1(oc8051_memory_interface1_n237), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n249), 
        .Y(oc8051_memory_interface1_n488) );
  XNOR3_X0P5M_A12TS oc8051_memory_interface1_u362 ( .A(
        oc8051_memory_interface1_n244), .B(oc8051_memory_interface1_n245), .C(
        oc8051_memory_interface1_n246), .Y(oc8051_memory_interface1_n242) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u361 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n241), 
        .B0(oc8051_memory_interface1_n237), .B1(oc8051_memory_interface1_n242), 
        .C0(oc8051_memory_interface1_n197), .C1(oc8051_memory_interface1_n243), 
        .Y(oc8051_memory_interface1_n489) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u360 ( .A(
        oc8051_memory_interface1_n234), .Y(oc8051_memory_interface1_n189) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u359 ( .A(
        oc8051_memory_interface1_n189), .B(oc8051_memory_interface1_n240), .Y(
        oc8051_memory_interface1_n238) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u358 ( .A0(
        oc8051_memory_interface1_n235), .A1(oc8051_memory_interface1_n236), 
        .B0(oc8051_memory_interface1_n237), .B1(oc8051_memory_interface1_n238), 
        .C0(oc8051_memory_interface1_n239), .C1(oc8051_memory_interface1_n197), 
        .Y(oc8051_memory_interface1_n490) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u357 ( .A(
        oc8051_memory_interface1_op_pos_0_), .B(oc8051_memory_interface1_n234), 
        .Y(oc8051_memory_interface1_n233) );
  XOR2_X0P5M_A12TS oc8051_memory_interface1_u356 ( .A(
        oc8051_memory_interface1_n195), .B(oc8051_memory_interface1_n196), .Y(
        oc8051_memory_interface1_n198) );
  XNOR2_X0P5M_A12TS oc8051_memory_interface1_u355 ( .A(
        oc8051_memory_interface1_n233), .B(oc8051_memory_interface1_n198), .Y(
        oc8051_memory_interface1_n232) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u354 ( .A(
        oc8051_memory_interface1_n232), .B(oc8051_memory_interface1_n197), .Y(
        oc8051_memory_interface1_n231) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u353 ( .A(
        oc8051_memory_interface1_n186), .B(oc8051_memory_interface1_n197), .Y(
        oc8051_memory_interface1_n199) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u352 ( .A(
        oc8051_memory_interface1_n199), .Y(oc8051_memory_interface1_n193) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u351 ( .A(
        oc8051_memory_interface1_n231), .B(oc8051_memory_interface1_n196), 
        .S0(oc8051_memory_interface1_n193), .Y(oc8051_memory_interface1_n491)
         );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u350 ( .A(
        oc8051_memory_interface1_op_pos_0_), .B(oc8051_memory_interface1_n193), 
        .Y(oc8051_memory_interface1_n230) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u349 ( .A(
        oc8051_memory_interface1_n230), .B(oc8051_memory_interface1_op_pos_0_), 
        .S0(oc8051_memory_interface1_n189), .Y(oc8051_memory_interface1_n229)
         );
  OAI22_X0P5M_A12TS oc8051_memory_interface1_u348 ( .A0(
        oc8051_memory_interface1_n188), .A1(oc8051_memory_interface1_n199), 
        .B0(oc8051_memory_interface1_pc_wr_r2), .B1(
        oc8051_memory_interface1_n229), .Y(oc8051_memory_interface1_n492) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u347 ( .A(
        oc8051_memory_interface1_idat_old_31_), .B(
        oc8051_memory_interface1_idat_cur_31_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n493) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u346 ( .A(
        oc8051_memory_interface1_n132), .Y(oc8051_memory_interface1_n204) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u345 ( .A(
        oc8051_memory_interface1_n168), .B(oc8051_memory_interface1_n134), .Y(
        oc8051_memory_interface1_n130) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u344 ( .A(
        oc8051_memory_interface1_n130), .Y(oc8051_memory_interface1_n205) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u343 ( .A0(wbi_dat_i[31]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n228) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u342 ( .A1N(
        oc8051_memory_interface1_idat_cur_31_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n228), 
        .Y(oc8051_memory_interface1_n494) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u341 ( .A(
        oc8051_memory_interface1_idat_old_30_), .B(
        oc8051_memory_interface1_idat_cur_30_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n495) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u340 ( .A0(wbi_dat_i[30]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n227) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u339 ( .A1N(
        oc8051_memory_interface1_idat_cur_30_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n227), 
        .Y(oc8051_memory_interface1_n496) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u338 ( .A(
        oc8051_memory_interface1_idat_old_29_), .B(
        oc8051_memory_interface1_idat_cur_29_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n497) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u337 ( .A0(wbi_dat_i[29]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n226) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u336 ( .A1N(
        oc8051_memory_interface1_idat_cur_29_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n226), 
        .Y(oc8051_memory_interface1_n498) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u335 ( .A(
        oc8051_memory_interface1_idat_old_28_), .B(
        oc8051_memory_interface1_idat_cur_28_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n499) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u334 ( .A0(wbi_dat_i[28]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n225) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u333 ( .A1N(
        oc8051_memory_interface1_idat_cur_28_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n225), 
        .Y(oc8051_memory_interface1_n500) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u332 ( .A(
        oc8051_memory_interface1_idat_old_27_), .B(
        oc8051_memory_interface1_idat_cur_27_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n501) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u331 ( .A0(wbi_dat_i[27]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n224) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u330 ( .A1N(
        oc8051_memory_interface1_idat_cur_27_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n224), 
        .Y(oc8051_memory_interface1_n502) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u329 ( .A(
        oc8051_memory_interface1_idat_old_26_), .B(
        oc8051_memory_interface1_idat_cur_26_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n503) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u328 ( .A0(wbi_dat_i[26]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n223) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u327 ( .A1N(
        oc8051_memory_interface1_idat_cur_26_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n223), 
        .Y(oc8051_memory_interface1_n504) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u326 ( .A(
        oc8051_memory_interface1_idat_old_25_), .B(
        oc8051_memory_interface1_idat_cur_25_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n505) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u325 ( .A0(wbi_dat_i[25]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n222) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u324 ( .A1N(
        oc8051_memory_interface1_idat_cur_25_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n222), 
        .Y(oc8051_memory_interface1_n506) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u323 ( .A(
        oc8051_memory_interface1_idat_old_24_), .B(
        oc8051_memory_interface1_idat_cur_24_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n507) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u322 ( .A0(wbi_dat_i[24]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n221) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u321 ( .A1N(
        oc8051_memory_interface1_idat_cur_24_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n221), 
        .Y(oc8051_memory_interface1_n508) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u320 ( .A(
        oc8051_memory_interface1_idat_old_23_), .B(
        oc8051_memory_interface1_idat_cur_23_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n509) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u319 ( .A0(wbi_dat_i[23]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n220) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u318 ( .A1N(
        oc8051_memory_interface1_idat_cur_23_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n220), 
        .Y(oc8051_memory_interface1_n510) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u317 ( .A(
        oc8051_memory_interface1_idat_old_22_), .B(
        oc8051_memory_interface1_idat_cur_22_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n511) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u316 ( .A0(wbi_dat_i[22]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n219) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u315 ( .A1N(
        oc8051_memory_interface1_idat_cur_22_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n219), 
        .Y(oc8051_memory_interface1_n512) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u314 ( .A(
        oc8051_memory_interface1_idat_old_21_), .B(
        oc8051_memory_interface1_idat_cur_21_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n513) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u313 ( .A0(wbi_dat_i[21]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n218) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u312 ( .A1N(
        oc8051_memory_interface1_idat_cur_21_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n218), 
        .Y(oc8051_memory_interface1_n514) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u311 ( .A(
        oc8051_memory_interface1_idat_old_20_), .B(
        oc8051_memory_interface1_idat_cur_20_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n515) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u310 ( .A0(wbi_dat_i[20]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n217) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u309 ( .A1N(
        oc8051_memory_interface1_idat_cur_20_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n217), 
        .Y(oc8051_memory_interface1_n516) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u308 ( .A(
        oc8051_memory_interface1_idat_old_19_), .B(
        oc8051_memory_interface1_idat_cur_19_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n517) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u307 ( .A0(wbi_dat_i[19]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n216) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u306 ( .A1N(
        oc8051_memory_interface1_idat_cur_19_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n216), 
        .Y(oc8051_memory_interface1_n518) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u305 ( .A(
        oc8051_memory_interface1_idat_old_18_), .B(
        oc8051_memory_interface1_idat_cur_18_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n519) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u304 ( .A0(wbi_dat_i[18]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n215) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u303 ( .A1N(
        oc8051_memory_interface1_idat_cur_18_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n215), 
        .Y(oc8051_memory_interface1_n520) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u302 ( .A(
        oc8051_memory_interface1_idat_old_17_), .B(
        oc8051_memory_interface1_idat_cur_17_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n521) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u301 ( .A0(wbi_dat_i[17]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n214) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u300 ( .A1N(
        oc8051_memory_interface1_idat_cur_17_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n214), 
        .Y(oc8051_memory_interface1_n522) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u299 ( .A(
        oc8051_memory_interface1_idat_old_16_), .B(
        oc8051_memory_interface1_idat_cur_16_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n523) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u298 ( .A0(wbi_dat_i[16]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n213) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u297 ( .A1N(
        oc8051_memory_interface1_idat_cur_16_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n213), 
        .Y(oc8051_memory_interface1_n524) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u296 ( .A(
        oc8051_memory_interface1_idat_old_15_), .B(
        oc8051_memory_interface1_idat_cur_15_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n525) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u295 ( .A0(wbi_dat_i[15]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n212) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u294 ( .A1N(
        oc8051_memory_interface1_idat_cur_15_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n212), 
        .Y(oc8051_memory_interface1_n526) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u293 ( .A(
        oc8051_memory_interface1_idat_old_14_), .B(
        oc8051_memory_interface1_idat_cur_14_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n527) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u292 ( .A0(wbi_dat_i[14]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n211) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u291 ( .A1N(
        oc8051_memory_interface1_idat_cur_14_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n211), 
        .Y(oc8051_memory_interface1_n528) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u290 ( .A(
        oc8051_memory_interface1_idat_old_13_), .B(
        oc8051_memory_interface1_idat_cur_13_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n529) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u289 ( .A0(wbi_dat_i[13]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n210) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u288 ( .A1N(
        oc8051_memory_interface1_idat_cur_13_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n210), 
        .Y(oc8051_memory_interface1_n530) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u287 ( .A(
        oc8051_memory_interface1_idat_old_12_), .B(
        oc8051_memory_interface1_idat_cur_12_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n531) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u286 ( .A0(wbi_dat_i[12]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n209) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u285 ( .A1N(
        oc8051_memory_interface1_idat_cur_12_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n209), 
        .Y(oc8051_memory_interface1_n532) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u284 ( .A(
        oc8051_memory_interface1_idat_old_11_), .B(
        oc8051_memory_interface1_idat_cur_11_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n533) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u283 ( .A0(wbi_dat_i[11]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n208) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u282 ( .A1N(
        oc8051_memory_interface1_idat_cur_11_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n208), 
        .Y(oc8051_memory_interface1_n534) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u281 ( .A(
        oc8051_memory_interface1_idat_old_10_), .B(
        oc8051_memory_interface1_idat_cur_10_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n535) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u280 ( .A0(wbi_dat_i[10]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n207) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u279 ( .A1N(
        oc8051_memory_interface1_idat_cur_10_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n207), 
        .Y(oc8051_memory_interface1_n536) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u278 ( .A(
        oc8051_memory_interface1_idat_old_9_), .B(
        oc8051_memory_interface1_idat_cur_9_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n537) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u277 ( .A0(wbi_dat_i[9]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n206) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u276 ( .A1N(
        oc8051_memory_interface1_idat_cur_9_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n206), 
        .Y(oc8051_memory_interface1_n538) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u275 ( .A(
        oc8051_memory_interface1_idat_old_8_), .B(
        oc8051_memory_interface1_idat_cur_8_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n539) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u274 ( .A0(wbi_dat_i[8]), .A1(
        oc8051_memory_interface1_n204), .B0(n2), .B1(
        oc8051_memory_interface1_n205), .Y(oc8051_memory_interface1_n203) );
  OAI2XB1_X0P5M_A12TS oc8051_memory_interface1_u273 ( .A1N(
        oc8051_memory_interface1_idat_cur_8_), .A0(
        oc8051_memory_interface1_n134), .B0(oc8051_memory_interface1_n203), 
        .Y(oc8051_memory_interface1_n540) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u272 ( .A(
        oc8051_memory_interface1_idat_old_7_), .B(
        oc8051_memory_interface1_idat_cur_7_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n541) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u271 ( .A(
        oc8051_memory_interface1_idat_old_6_), .B(
        oc8051_memory_interface1_idat_cur_6_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n543) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u270 ( .A(
        oc8051_memory_interface1_idat_old_5_), .B(
        oc8051_memory_interface1_idat_cur_5_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n545) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u269 ( .A(
        oc8051_memory_interface1_idat_old_4_), .B(
        oc8051_memory_interface1_idat_cur_4_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n547) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u268 ( .A(
        oc8051_memory_interface1_idat_old_3_), .B(
        oc8051_memory_interface1_idat_cur_3_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n549) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u267 ( .A(
        oc8051_memory_interface1_idat_old_2_), .B(
        oc8051_memory_interface1_idat_cur_2_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n551) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u266 ( .A(
        oc8051_memory_interface1_idat_old_1_), .B(
        oc8051_memory_interface1_idat_cur_1_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n553) );
  MXT2_X0P5M_A12TS oc8051_memory_interface1_u265 ( .A(
        oc8051_memory_interface1_idat_old_0_), .B(
        oc8051_memory_interface1_idat_cur_0_), .S0(
        oc8051_memory_interface1_n134), .Y(oc8051_memory_interface1_n555) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u264 ( .A(
        oc8051_memory_interface1_n202), .B(oc8051_memory_interface1_op_pos_1_), 
        .C(oc8051_memory_interface1_n195), .Y(oc8051_memory_interface1_n201)
         );
  AOI31_X0P5M_A12TS oc8051_memory_interface1_u263 ( .A0(
        oc8051_memory_interface1_n198), .A1(oc8051_memory_interface1_n199), 
        .A2(oc8051_memory_interface1_n200), .B0(oc8051_memory_interface1_n201), 
        .Y(oc8051_memory_interface1_n190) );
  OAI31_X0P5M_A12TS oc8051_memory_interface1_u262 ( .A0(
        oc8051_memory_interface1_n194), .A1(oc8051_memory_interface1_n195), 
        .A2(oc8051_memory_interface1_n196), .B0(oc8051_memory_interface1_n197), 
        .Y(oc8051_memory_interface1_n192) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u261 ( .A(
        oc8051_memory_interface1_n192), .B(oc8051_memory_interface1_op_pos_2_), 
        .S0(oc8051_memory_interface1_n193), .Y(oc8051_memory_interface1_n191)
         );
  OAI31_X0P5M_A12TS oc8051_memory_interface1_u260 ( .A0(
        oc8051_memory_interface1_n188), .A1(oc8051_memory_interface1_n189), 
        .A2(oc8051_memory_interface1_n190), .B0(oc8051_memory_interface1_n191), 
        .Y(oc8051_memory_interface1_n557) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u259 ( .A(
        oc8051_memory_interface1_n186), .B(oc8051_memory_interface1_pc_wr_r2), 
        .C(oc8051_memory_interface1_n187), .Y(oc8051_memory_interface1_n184)
         );
  OAI21B_X0P5M_A12TS oc8051_memory_interface1_u258 ( .A0(
        oc8051_memory_interface1_n184), .A1(oc8051_memory_interface1_n185), 
        .B0N(intr), .Y(oc8051_memory_interface1_n558) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u257 ( .A(wbd_ack_i), .B(
        mem_act[1]), .Y(oc8051_memory_interface1_n173) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u256 ( .A(
        oc8051_memory_interface1_n183), .B(wbd_ack_i), .Y(
        oc8051_memory_interface1_n175) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u255 ( .A0(dptr_lo[0]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[0]), .Y(oc8051_memory_interface1_n182) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u254 ( .B0(wbd_adr_o[0]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n182), .Y(
        oc8051_memory_interface1_n559) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u253 ( .A0(dptr_lo[1]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[1]), .Y(oc8051_memory_interface1_n181) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u252 ( .B0(wbd_adr_o[1]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n181), .Y(
        oc8051_memory_interface1_n560) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u251 ( .A0(dptr_lo[2]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[2]), .Y(oc8051_memory_interface1_n180) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u250 ( .B0(wbd_adr_o[2]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n180), .Y(
        oc8051_memory_interface1_n561) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u249 ( .A0(dptr_lo[3]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[3]), .Y(oc8051_memory_interface1_n179) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u248 ( .B0(wbd_adr_o[3]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n179), .Y(
        oc8051_memory_interface1_n562) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u247 ( .A0(dptr_lo[4]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[4]), .Y(oc8051_memory_interface1_n178) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u246 ( .B0(wbd_adr_o[4]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n178), .Y(
        oc8051_memory_interface1_n563) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u245 ( .A0(dptr_lo[5]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[5]), .Y(oc8051_memory_interface1_n177) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u244 ( .B0(wbd_adr_o[5]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n177), .Y(
        oc8051_memory_interface1_n564) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u243 ( .A0(dptr_lo[6]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[6]), .Y(oc8051_memory_interface1_n176) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u242 ( .B0(wbd_adr_o[6]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n176), .Y(
        oc8051_memory_interface1_n565) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u241 ( .A0(dptr_lo[7]), .A1(
        oc8051_memory_interface1_n173), .B0(oc8051_memory_interface1_n175), 
        .B1(ri[7]), .Y(oc8051_memory_interface1_n174) );
  AO1B2_X0P5M_A12TS oc8051_memory_interface1_u240 ( .B0(wbd_adr_o[7]), .B1(
        wbd_ack_i), .A0N(oc8051_memory_interface1_n174), .Y(
        oc8051_memory_interface1_n566) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u239 ( .A0(wbd_adr_o[8]), .A1(
        wbd_ack_i), .B0(dptr_hi[0]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n567) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u238 ( .A0(wbd_adr_o[9]), .A1(
        wbd_ack_i), .B0(dptr_hi[1]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n568) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u237 ( .A0(wbd_adr_o[10]), .A1(
        wbd_ack_i), .B0(dptr_hi[2]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n569) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u236 ( .A0(wbd_adr_o[11]), .A1(
        wbd_ack_i), .B0(dptr_hi[3]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n570) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u235 ( .A0(wbd_adr_o[12]), .A1(
        wbd_ack_i), .B0(dptr_hi[4]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n571) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u234 ( .A0(wbd_adr_o[13]), .A1(
        wbd_ack_i), .B0(dptr_hi[5]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n572) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u233 ( .A0(wbd_adr_o[14]), .A1(
        wbd_ack_i), .B0(dptr_hi[6]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n573) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u232 ( .A0(wbd_adr_o[15]), .A1(
        wbd_ack_i), .B0(dptr_hi[7]), .B1(oc8051_memory_interface1_n173), .Y(
        oc8051_memory_interface1_n574) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u231 ( .A0(wbd_dat_o[0]), .A1(
        wbd_ack_i), .B0(acc[0]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n575) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u230 ( .A0(wbd_dat_o[1]), .A1(
        wbd_ack_i), .B0(acc[1]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n576) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u229 ( .A0(wbd_dat_o[2]), .A1(
        wbd_ack_i), .B0(acc[2]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n577) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u228 ( .A0(wbd_dat_o[3]), .A1(
        wbd_ack_i), .B0(acc[3]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n578) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u227 ( .A0(wbd_dat_o[4]), .A1(
        wbd_ack_i), .B0(acc[4]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n579) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u226 ( .A0(wbd_dat_o[5]), .A1(
        wbd_ack_i), .B0(acc[5]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n580) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u225 ( .A0(wbd_dat_o[6]), .A1(
        wbd_ack_i), .B0(acc[6]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n581) );
  AO22_X0P5M_A12TS oc8051_memory_interface1_u224 ( .A0(wbd_dat_o[7]), .A1(
        wbd_ack_i), .B0(acc[7]), .B1(oc8051_memory_interface1_n1310), .Y(
        oc8051_memory_interface1_n582) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u223 ( .A(
        oc8051_memory_interface1_imem_wait), .Y(oc8051_memory_interface1_n170)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u222 ( .A0(
        oc8051_memory_interface1_n172), .A1(oc8051_memory_interface1_n170), 
        .B0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n583)
         );
  OAI21_X0P5M_A12TS oc8051_memory_interface1_u221 ( .A0(
        oc8051_memory_interface1_n169), .A1(oc8051_memory_interface1_n170), 
        .B0(oc8051_memory_interface1_n171), .Y(oc8051_memory_interface1_n584)
         );
  INV_X0P5B_A12TS oc8051_memory_interface1_u220 ( .A(wbd_ack_i), .Y(
        oc8051_memory_interface1_n813) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u219 ( .A(n2), .Y(
        oc8051_memory_interface1_n131) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u218 ( .A(
        oc8051_memory_interface1_istb_t), .B(oc8051_memory_interface1_n168), 
        .Y(oc8051_memory_interface1_n157) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u217 ( .A(wbi_dat_i[7]), .Y(
        oc8051_memory_interface1_n133) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u216 ( .A(
        oc8051_memory_interface1_istb_t), .B(oc8051_memory_interface1_n167), 
        .Y(oc8051_memory_interface1_n158) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u215 ( .A(
        oc8051_memory_interface1_cdata_7_), .Y(oc8051_memory_interface1_n166)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u214 ( .A0(
        oc8051_memory_interface1_n131), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n133), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n166), .Y(oc8051_memory_interface1_n804) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u213 ( .A(n2), .Y(
        oc8051_memory_interface1_n136) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u212 ( .A(wbi_dat_i[6]), .Y(
        oc8051_memory_interface1_n137) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u211 ( .A(
        oc8051_memory_interface1_cdata_6_), .Y(oc8051_memory_interface1_n165)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u210 ( .A0(
        oc8051_memory_interface1_n136), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n137), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n165), .Y(oc8051_memory_interface1_n803) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u209 ( .A(n2), .Y(
        oc8051_memory_interface1_n139) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u208 ( .A(wbi_dat_i[5]), .Y(
        oc8051_memory_interface1_n140) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u207 ( .A(
        oc8051_memory_interface1_cdata_5_), .Y(oc8051_memory_interface1_n164)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u206 ( .A0(
        oc8051_memory_interface1_n139), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n140), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n164), .Y(oc8051_memory_interface1_n802) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u205 ( .A(n2), .Y(
        oc8051_memory_interface1_n142) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u204 ( .A(wbi_dat_i[4]), .Y(
        oc8051_memory_interface1_n143) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u203 ( .A(
        oc8051_memory_interface1_cdata_4_), .Y(oc8051_memory_interface1_n163)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u202 ( .A0(
        oc8051_memory_interface1_n142), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n143), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n163), .Y(oc8051_memory_interface1_n801) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u201 ( .A(n2), .Y(
        oc8051_memory_interface1_n145) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u200 ( .A(wbi_dat_i[3]), .Y(
        oc8051_memory_interface1_n146) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u199 ( .A(
        oc8051_memory_interface1_cdata_3_), .Y(oc8051_memory_interface1_n162)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u198 ( .A0(
        oc8051_memory_interface1_n145), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n146), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n162), .Y(oc8051_memory_interface1_n800) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u197 ( .A(n2), .Y(
        oc8051_memory_interface1_n148) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u196 ( .A(wbi_dat_i[2]), .Y(
        oc8051_memory_interface1_n149) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u195 ( .A(
        oc8051_memory_interface1_cdata_2_), .Y(oc8051_memory_interface1_n161)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u194 ( .A0(
        oc8051_memory_interface1_n148), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n149), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n161), .Y(oc8051_memory_interface1_n799) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u193 ( .A(n2), .Y(
        oc8051_memory_interface1_n151) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u192 ( .A(wbi_dat_i[1]), .Y(
        oc8051_memory_interface1_n152) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u191 ( .A(
        oc8051_memory_interface1_cdata_1_), .Y(oc8051_memory_interface1_n160)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u190 ( .A0(
        oc8051_memory_interface1_n151), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n152), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n160), .Y(oc8051_memory_interface1_n798) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u189 ( .A(n2), .Y(
        oc8051_memory_interface1_n154) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u188 ( .A(wbi_dat_i[0]), .Y(
        oc8051_memory_interface1_n155) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u187 ( .A(
        oc8051_memory_interface1_cdata_0_), .Y(oc8051_memory_interface1_n159)
         );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u186 ( .A0(
        oc8051_memory_interface1_n154), .A1(oc8051_memory_interface1_n157), 
        .B0(oc8051_memory_interface1_n155), .B1(oc8051_memory_interface1_n158), 
        .C0(oc8051_memory_interface1_istb_t), .C1(
        oc8051_memory_interface1_n159), .Y(oc8051_memory_interface1_n797) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u185 ( .A(
        oc8051_memory_interface1_idat_cur_0_), .Y(
        oc8051_memory_interface1_n156) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u184 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n154), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n155), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n156), 
        .Y(oc8051_memory_interface1_n796) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u183 ( .A(
        oc8051_memory_interface1_idat_cur_1_), .Y(
        oc8051_memory_interface1_n153) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u182 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n151), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n152), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n153), 
        .Y(oc8051_memory_interface1_n795) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u181 ( .A(
        oc8051_memory_interface1_idat_cur_2_), .Y(
        oc8051_memory_interface1_n150) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u180 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n148), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n149), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n150), 
        .Y(oc8051_memory_interface1_n794) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u179 ( .A(
        oc8051_memory_interface1_idat_cur_3_), .Y(
        oc8051_memory_interface1_n147) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u178 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n145), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n146), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n147), 
        .Y(oc8051_memory_interface1_n793) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u177 ( .A(
        oc8051_memory_interface1_idat_cur_4_), .Y(
        oc8051_memory_interface1_n144) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u176 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n142), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n143), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n144), 
        .Y(oc8051_memory_interface1_n792) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u175 ( .A(
        oc8051_memory_interface1_idat_cur_5_), .Y(
        oc8051_memory_interface1_n141) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u174 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n139), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n140), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n141), 
        .Y(oc8051_memory_interface1_n791) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u173 ( .A(
        oc8051_memory_interface1_idat_cur_6_), .Y(
        oc8051_memory_interface1_n138) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u172 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n136), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n137), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n138), 
        .Y(oc8051_memory_interface1_n790) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u171 ( .A(
        oc8051_memory_interface1_idat_cur_7_), .Y(
        oc8051_memory_interface1_n135) );
  OAI222_X0P5M_A12TS oc8051_memory_interface1_u170 ( .A0(
        oc8051_memory_interface1_n130), .A1(oc8051_memory_interface1_n131), 
        .B0(oc8051_memory_interface1_n132), .B1(oc8051_memory_interface1_n133), 
        .C0(oc8051_memory_interface1_n134), .C1(oc8051_memory_interface1_n135), 
        .Y(oc8051_memory_interface1_n789) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u169 ( .A(ram_rd_sel[2]), .Y(
        oc8051_memory_interface1_n99) );
  NAND3_X0P5A_A12TS oc8051_memory_interface1_u168 ( .A(
        oc8051_memory_interface1_n113), .B(oc8051_memory_interface1_n99), .C(
        ram_rd_sel[1]), .Y(oc8051_memory_interface1_n104) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u167 ( .A(ram_rd_sel[1]), .Y(
        oc8051_memory_interface1_n105) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u166 ( .AN(
        oc8051_memory_interface1_n830), .B(oc8051_memory_interface1_n105), .Y(
        oc8051_memory_interface1_n101) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u165 ( .A(sp[0]), .B(
        oc8051_memory_interface1_n101), .Y(oc8051_memory_interface1_n128) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u164 ( .A(
        oc8051_memory_interface1_n830), .B(oc8051_memory_interface1_n105), .Y(
        oc8051_memory_interface1_n97) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u163 ( .A(
        oc8051_memory_interface1_n97), .Y(oc8051_memory_interface1_n107) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u162 ( .A(ram_rd_sel[1]), .B(
        ram_rd_sel[2]), .C(ram_rd_sel[0]), .Y(oc8051_memory_interface1_n117)
         );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u161 ( .A0(ri[0]), .A1(
        oc8051_memory_interface1_n107), .B0(op1_cur[0]), .B1(
        oc8051_memory_interface1_n117), .Y(oc8051_memory_interface1_n129) );
  AOI32_X0P5M_A12TS oc8051_memory_interface1_u160 ( .A0(ram_rd_sel[0]), .A1(
        oc8051_memory_interface1_n105), .A2(ram_rd_sel[2]), .B0(ri[1]), .B1(
        oc8051_memory_interface1_n107), .Y(oc8051_memory_interface1_n124) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u159 ( .A(op1_cur[1]), .B(
        oc8051_memory_interface1_n117), .Y(oc8051_memory_interface1_n125) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u158 ( .A(
        oc8051_memory_interface1_n104), .Y(oc8051_memory_interface1_n102) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u157 ( .A0(sp[1]), .A1(
        oc8051_memory_interface1_n101), .B0(oc8051_memory_interface1_n102), 
        .B1(op2_n[1]), .Y(oc8051_memory_interface1_n126) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u156 ( .A(sp[2]), .B(
        oc8051_memory_interface1_n101), .Y(oc8051_memory_interface1_n122) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u155 ( .A0(ri[2]), .A1(
        oc8051_memory_interface1_n107), .B0(op1_cur[2]), .B1(
        oc8051_memory_interface1_n117), .Y(oc8051_memory_interface1_n123) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u154 ( .A(sp[3]), .B(
        oc8051_memory_interface1_n101), .Y(oc8051_memory_interface1_n119) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u153 ( .A0(ri[3]), .A1(
        oc8051_memory_interface1_n107), .B0(bank_sel[0]), .B1(
        oc8051_memory_interface1_n117), .Y(oc8051_memory_interface1_n120) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u152 ( .A0(
        oc8051_memory_interface1_n118), .A1(oc8051_memory_interface1_n104), 
        .B0(oc8051_memory_interface1_n119), .C0(oc8051_memory_interface1_n120), 
        .Y(rd_addr[3]) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u151 ( .A(sp[4]), .B(
        oc8051_memory_interface1_n101), .Y(oc8051_memory_interface1_n115) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u150 ( .A(
        oc8051_memory_interface1_n99), .B(ram_rd_sel[0]), .Y(
        oc8051_memory_interface1_n108) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u149 ( .A0(bank_sel[1]), .A1(
        oc8051_memory_interface1_n117), .B0(ri[4]), .B1(
        oc8051_memory_interface1_n107), .C0(oc8051_memory_interface1_n108), 
        .Y(oc8051_memory_interface1_n116) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u148 ( .A0(
        oc8051_memory_interface1_n114), .A1(oc8051_memory_interface1_n104), 
        .B0(oc8051_memory_interface1_n115), .C0(oc8051_memory_interface1_n116), 
        .Y(rd_addr[4]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u147 ( .A(
        oc8051_memory_interface1_n113), .B(oc8051_memory_interface1_n99), .Y(
        oc8051_memory_interface1_n112) );
  MXIT2_X0P5M_A12TS oc8051_memory_interface1_u146 ( .A(
        oc8051_memory_interface1_n108), .B(oc8051_memory_interface1_n112), 
        .S0(ram_rd_sel[1]), .Y(oc8051_memory_interface1_n110) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u145 ( .A0(ri[5]), .A1(
        oc8051_memory_interface1_n107), .B0(sp[5]), .B1(
        oc8051_memory_interface1_n101), .Y(oc8051_memory_interface1_n111) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u144 ( .A0(
        oc8051_memory_interface1_n109), .A1(oc8051_memory_interface1_n104), 
        .B0(oc8051_memory_interface1_n110), .C0(oc8051_memory_interface1_n111), 
        .Y(rd_addr[5]) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u143 ( .A0(sp[6]), .A1(
        oc8051_memory_interface1_n101), .B0(ri[6]), .B1(
        oc8051_memory_interface1_n107), .C0(oc8051_memory_interface1_n108), 
        .Y(oc8051_memory_interface1_n106) );
  OAI221_X0P5M_A12TS oc8051_memory_interface1_u142 ( .A0(
        oc8051_memory_interface1_n103), .A1(oc8051_memory_interface1_n104), 
        .B0(oc8051_memory_interface1_n105), .B1(oc8051_memory_interface1_n99), 
        .C0(oc8051_memory_interface1_n106), .Y(rd_addr[6]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u141 ( .A(ri[7]), .Y(
        oc8051_memory_interface1_n98) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u140 ( .A0(sp[7]), .A1(
        oc8051_memory_interface1_n101), .B0(oc8051_memory_interface1_n102), 
        .B1(op2_n[7]), .Y(oc8051_memory_interface1_n100) );
  OAI211_X0P5M_A12TS oc8051_memory_interface1_u139 ( .A0(
        oc8051_memory_interface1_n97), .A1(oc8051_memory_interface1_n98), .B0(
        oc8051_memory_interface1_n99), .C0(oc8051_memory_interface1_n100), .Y(
        rd_addr[7]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u138 ( .A(
        oc8051_memory_interface1_n397), .Y(pc[9]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u137 ( .A(
        oc8051_memory_interface1_n395), .Y(pc[11]) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u136 ( .A(
        oc8051_memory_interface1_n393), .Y(pc[13]) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u135 ( .A(
        oc8051_memory_interface1_n86), .B(ram_wr_sel[0]), .Y(
        oc8051_memory_interface1_n79) );
  NOR2_X0P5A_A12TS oc8051_memory_interface1_u134 ( .A(ram_wr_sel[0]), .B(
        ram_wr_sel[1]), .Y(oc8051_memory_interface1_n87) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u133 ( .A0(
        oc8051_memory_interface1_ri_r[0]), .A1(oc8051_memory_interface1_n79), 
        .B0(oc8051_memory_interface1_rn_r[0]), .B1(
        oc8051_memory_interface1_n87), .Y(oc8051_memory_interface1_n94) );
  INV_X0P5B_A12TS oc8051_memory_interface1_u132 ( .A(ram_wr_sel[0]), .Y(
        oc8051_memory_interface1_n96) );
  NOR3_X0P5A_A12TS oc8051_memory_interface1_u131 ( .A(ram_wr_sel[1]), .B(
        ram_wr_sel[2]), .C(oc8051_memory_interface1_n96), .Y(
        oc8051_memory_interface1_n78) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u130 ( .AN(ram_wr_sel[2]), .B(
        ram_wr_sel[1]), .Y(oc8051_memory_interface1_n76) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u129 ( .AN(wr_ind), .B(
        oc8051_memory_interface1_n96), .Y(oc8051_memory_interface1_n75) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u128 ( .A0(
        oc8051_memory_interface1_imm_r[0]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_imm2_r[0]), .B1(
        oc8051_memory_interface1_n76), .C0(sp_w[0]), .C1(
        oc8051_memory_interface1_n75), .Y(oc8051_memory_interface1_n95) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u127 ( .A0(
        oc8051_memory_interface1_ri_r[1]), .A1(oc8051_memory_interface1_n79), 
        .B0(oc8051_memory_interface1_rn_r[1]), .B1(
        oc8051_memory_interface1_n87), .Y(oc8051_memory_interface1_n92) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u126 ( .A0(
        oc8051_memory_interface1_imm_r[1]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_imm2_r[1]), .B1(
        oc8051_memory_interface1_n76), .C0(sp_w[1]), .C1(
        oc8051_memory_interface1_n75), .Y(oc8051_memory_interface1_n93) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u125 ( .A0(
        oc8051_memory_interface1_ri_r[2]), .A1(oc8051_memory_interface1_n79), 
        .B0(oc8051_memory_interface1_rn_r[2]), .B1(
        oc8051_memory_interface1_n87), .Y(oc8051_memory_interface1_n90) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u124 ( .A0(
        oc8051_memory_interface1_imm_r[2]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_imm2_r[2]), .B1(
        oc8051_memory_interface1_n76), .C0(sp_w[2]), .C1(
        oc8051_memory_interface1_n75), .Y(oc8051_memory_interface1_n91) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u123 ( .A0(
        oc8051_memory_interface1_ri_r[3]), .A1(oc8051_memory_interface1_n79), 
        .B0(oc8051_memory_interface1_rn_r[3]), .B1(
        oc8051_memory_interface1_n87), .Y(oc8051_memory_interface1_n88) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u122 ( .A0(
        oc8051_memory_interface1_imm_r[3]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_imm2_r[3]), .B1(
        oc8051_memory_interface1_n76), .C0(sp_w[3]), .C1(
        oc8051_memory_interface1_n75), .Y(oc8051_memory_interface1_n89) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u121 ( .A(
        oc8051_memory_interface1_n88), .B(oc8051_memory_interface1_n89), .Y(
        wr_addr[3]) );
  AOI222_X0P5M_A12TS oc8051_memory_interface1_u120 ( .A0(
        oc8051_memory_interface1_rn_r[4]), .A1(oc8051_memory_interface1_n87), 
        .B0(oc8051_memory_interface1_imm_r[4]), .B1(
        oc8051_memory_interface1_n78), .C0(oc8051_memory_interface1_ri_r[4]), 
        .C1(oc8051_memory_interface1_n79), .Y(oc8051_memory_interface1_n84) );
  NOR2B_X0P5M_A12TS oc8051_memory_interface1_u119 ( .AN(ram_wr_sel[2]), .B(
        oc8051_memory_interface1_n86), .Y(oc8051_memory_interface1_n77) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u118 ( .A0(sp_w[4]), .A1(
        oc8051_memory_interface1_n75), .B0(oc8051_memory_interface1_imm2_r[4]), 
        .B1(oc8051_memory_interface1_n76), .C0(oc8051_memory_interface1_n77), 
        .Y(oc8051_memory_interface1_n85) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u117 ( .A(
        oc8051_memory_interface1_n84), .B(oc8051_memory_interface1_n85), .Y(
        wr_addr[4]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u116 ( .A0(
        oc8051_memory_interface1_imm_r[5]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_ri_r[5]), .B1(
        oc8051_memory_interface1_n79), .Y(oc8051_memory_interface1_n82) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u115 ( .A0(sp_w[5]), .A1(
        oc8051_memory_interface1_n75), .B0(oc8051_memory_interface1_imm2_r[5]), 
        .B1(oc8051_memory_interface1_n76), .C0(oc8051_memory_interface1_n77), 
        .Y(oc8051_memory_interface1_n83) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u114 ( .A(
        oc8051_memory_interface1_n82), .B(oc8051_memory_interface1_n83), .Y(
        wr_addr[5]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u113 ( .A0(
        oc8051_memory_interface1_imm_r[6]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_ri_r[6]), .B1(
        oc8051_memory_interface1_n79), .Y(oc8051_memory_interface1_n80) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u112 ( .A0(sp_w[6]), .A1(
        oc8051_memory_interface1_n75), .B0(oc8051_memory_interface1_imm2_r[6]), 
        .B1(oc8051_memory_interface1_n76), .C0(oc8051_memory_interface1_n77), 
        .Y(oc8051_memory_interface1_n81) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u111 ( .A(
        oc8051_memory_interface1_n80), .B(oc8051_memory_interface1_n81), .Y(
        wr_addr[6]) );
  AOI22_X0P5M_A12TS oc8051_memory_interface1_u110 ( .A0(
        oc8051_memory_interface1_imm_r[7]), .A1(oc8051_memory_interface1_n78), 
        .B0(oc8051_memory_interface1_ri_r[7]), .B1(
        oc8051_memory_interface1_n79), .Y(oc8051_memory_interface1_n73) );
  AOI221_X0P5M_A12TS oc8051_memory_interface1_u109 ( .A0(sp_w[7]), .A1(
        oc8051_memory_interface1_n75), .B0(oc8051_memory_interface1_imm2_r[7]), 
        .B1(oc8051_memory_interface1_n76), .C0(oc8051_memory_interface1_n77), 
        .Y(oc8051_memory_interface1_n74) );
  NAND2_X0P5A_A12TS oc8051_memory_interface1_u108 ( .A(
        oc8051_memory_interface1_n73), .B(oc8051_memory_interface1_n74), .Y(
        wr_addr[7]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u107 ( .A(
        oc8051_memory_interface1_idat_old_1_), .B(
        oc8051_memory_interface1_idat_old_9_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n50)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u106 ( .A(
        oc8051_memory_interface1_idat_cur_9_), .Y(oc8051_memory_interface1_n58) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u105 ( .A(
        oc8051_memory_interface1_n50), .B(oc8051_memory_interface1_n4), .C(
        oc8051_memory_interface1_n5), .D(oc8051_memory_interface1_n58), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_1_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u104 ( .A(
        oc8051_memory_interface1_idat_old_4_), .B(
        oc8051_memory_interface1_idat_old_12_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n53)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u103 ( .A(
        oc8051_memory_interface1_idat_cur_12_), .Y(
        oc8051_memory_interface1_n61) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u102 ( .A(
        oc8051_memory_interface1_n53), .B(oc8051_memory_interface1_n13), .C(
        oc8051_memory_interface1_n14), .D(oc8051_memory_interface1_n61), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_4_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u101 ( .A(
        oc8051_memory_interface1_idat_old_2_), .B(
        oc8051_memory_interface1_idat_old_10_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n51)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u100 ( .A(
        oc8051_memory_interface1_idat_cur_10_), .Y(
        oc8051_memory_interface1_n59) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u99 ( .A(
        oc8051_memory_interface1_n51), .B(oc8051_memory_interface1_n7), .C(
        oc8051_memory_interface1_n8), .D(oc8051_memory_interface1_n59), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_2_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u98 ( .A(
        oc8051_memory_interface1_idat_old_0_), .B(
        oc8051_memory_interface1_idat_old_8_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n49)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u97 ( .A(
        oc8051_memory_interface1_idat_cur_8_), .Y(oc8051_memory_interface1_n57) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u96 ( .A(
        oc8051_memory_interface1_n49), .B(oc8051_memory_interface1_n1), .C(
        oc8051_memory_interface1_n2), .D(oc8051_memory_interface1_n57), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_0_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u95 ( .A(
        oc8051_memory_interface1_idat_old_5_), .B(
        oc8051_memory_interface1_idat_old_13_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n54)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u94 ( .A(
        oc8051_memory_interface1_idat_cur_13_), .Y(
        oc8051_memory_interface1_n62) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u93 ( .A(
        oc8051_memory_interface1_n54), .B(oc8051_memory_interface1_n16), .C(
        oc8051_memory_interface1_n17), .D(oc8051_memory_interface1_n62), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_5_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u92 ( .A(
        oc8051_memory_interface1_idat_old_7_), .B(
        oc8051_memory_interface1_idat_old_15_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n56)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u91 ( .A(
        oc8051_memory_interface1_idat_cur_15_), .Y(
        oc8051_memory_interface1_n64) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u90 ( .A(
        oc8051_memory_interface1_n56), .B(oc8051_memory_interface1_n22), .C(
        oc8051_memory_interface1_n23), .D(oc8051_memory_interface1_n64), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_7_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u89 ( .A(
        oc8051_memory_interface1_idat_old_6_), .B(
        oc8051_memory_interface1_idat_old_14_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n55)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u88 ( .A(
        oc8051_memory_interface1_idat_cur_14_), .Y(
        oc8051_memory_interface1_n63) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u87 ( .A(
        oc8051_memory_interface1_n55), .B(oc8051_memory_interface1_n19), .C(
        oc8051_memory_interface1_n20), .D(oc8051_memory_interface1_n63), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_6_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u86 ( .A(
        oc8051_memory_interface1_idat_old_3_), .B(
        oc8051_memory_interface1_idat_old_11_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n52)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u85 ( .A(
        oc8051_memory_interface1_idat_cur_11_), .Y(
        oc8051_memory_interface1_n60) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u84 ( .A(
        oc8051_memory_interface1_n52), .B(oc8051_memory_interface1_n10), .C(
        oc8051_memory_interface1_n11), .D(oc8051_memory_interface1_n60), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op1_3_) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u83 ( .A(
        oc8051_memory_interface1_idat_cur_23_), .B(
        oc8051_memory_interface1_idat_cur_31_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n24)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u82 ( .A(
        oc8051_memory_interface1_idat_cur_22_), .B(
        oc8051_memory_interface1_idat_cur_30_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n21)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u81 ( .A(
        oc8051_memory_interface1_idat_cur_21_), .B(
        oc8051_memory_interface1_idat_cur_29_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n18)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u80 ( .A(
        oc8051_memory_interface1_idat_cur_20_), .B(
        oc8051_memory_interface1_idat_cur_28_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n15)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u79 ( .A(
        oc8051_memory_interface1_idat_cur_19_), .B(
        oc8051_memory_interface1_idat_cur_27_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n12)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u78 ( .A(
        oc8051_memory_interface1_idat_cur_18_), .B(
        oc8051_memory_interface1_idat_cur_26_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n9)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u77 ( .A(
        oc8051_memory_interface1_idat_cur_16_), .B(
        oc8051_memory_interface1_idat_cur_24_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n3)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u76 ( .A(
        oc8051_memory_interface1_idat_cur_7_), .B(
        oc8051_memory_interface1_idat_cur_15_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n23)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u75 ( .A(
        oc8051_memory_interface1_idat_cur_6_), .B(
        oc8051_memory_interface1_idat_cur_14_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n20)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u74 ( .A(
        oc8051_memory_interface1_idat_cur_5_), .B(
        oc8051_memory_interface1_idat_cur_13_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n17)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u73 ( .A(
        oc8051_memory_interface1_idat_cur_4_), .B(
        oc8051_memory_interface1_idat_cur_12_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n14)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u72 ( .A(
        oc8051_memory_interface1_idat_cur_3_), .B(
        oc8051_memory_interface1_idat_cur_11_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n11)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u71 ( .A(
        oc8051_memory_interface1_idat_cur_2_), .B(
        oc8051_memory_interface1_idat_cur_10_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n8)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u70 ( .A(
        oc8051_memory_interface1_idat_cur_0_), .B(
        oc8051_memory_interface1_idat_cur_8_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n2)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u69 ( .A(
        oc8051_memory_interface1_idat_cur_1_), .B(
        oc8051_memory_interface1_idat_cur_9_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n5)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u68 ( .A(
        oc8051_memory_interface1_idat_old_23_), .B(
        oc8051_memory_interface1_idat_old_31_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n22)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u67 ( .A(
        oc8051_memory_interface1_idat_old_22_), .B(
        oc8051_memory_interface1_idat_old_30_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n19)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u66 ( .A(
        oc8051_memory_interface1_idat_old_21_), .B(
        oc8051_memory_interface1_idat_old_29_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n16)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u65 ( .A(
        oc8051_memory_interface1_idat_old_20_), .B(
        oc8051_memory_interface1_idat_old_28_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n13)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u64 ( .A(
        oc8051_memory_interface1_idat_old_19_), .B(
        oc8051_memory_interface1_idat_old_27_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n10)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u63 ( .A(
        oc8051_memory_interface1_idat_old_18_), .B(
        oc8051_memory_interface1_idat_old_26_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n7)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u62 ( .A(
        oc8051_memory_interface1_idat_old_16_), .B(
        oc8051_memory_interface1_idat_old_24_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n1)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u61 ( .A(
        oc8051_memory_interface1_idat_old_17_), .B(
        oc8051_memory_interface1_idat_old_25_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n4)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u60 ( .A(
        oc8051_memory_interface1_idat_cur_31_), .Y(
        oc8051_memory_interface1_n72) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u59 ( .A(
        oc8051_memory_interface1_n22), .B(oc8051_memory_interface1_n23), .C(
        oc8051_memory_interface1_n24), .D(oc8051_memory_interface1_n72), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[7]) );
  MXT2_X1M_A12TS oc8051_memory_interface1_u58 ( .A(
        oc8051_memory_interface1_idat_old_31_), .B(
        oc8051_memory_interface1_idat_cur_7_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n46)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u57 ( .A(
        oc8051_memory_interface1_idat_old_26_), .B(
        oc8051_memory_interface1_idat_cur_2_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n31)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u56 ( .A(
        oc8051_memory_interface1_idat_old_24_), .B(
        oc8051_memory_interface1_idat_cur_0_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n25)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u55 ( .A(
        oc8051_memory_interface1_idat_old_25_), .B(
        oc8051_memory_interface1_idat_cur_1_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n28)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u54 ( .A(
        oc8051_memory_interface1_idat_old_28_), .B(
        oc8051_memory_interface1_idat_cur_4_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n37)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u53 ( .A(
        oc8051_memory_interface1_idat_old_30_), .B(
        oc8051_memory_interface1_idat_cur_6_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n43)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u52 ( .A(
        oc8051_memory_interface1_idat_old_27_), .B(
        oc8051_memory_interface1_idat_cur_3_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n34)
         );
  MXT2_X1M_A12TS oc8051_memory_interface1_u51 ( .A(
        oc8051_memory_interface1_idat_old_29_), .B(
        oc8051_memory_interface1_idat_cur_5_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n40)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u50 ( .A(
        oc8051_memory_interface1_idat_cur_30_), .Y(
        oc8051_memory_interface1_n71) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u49 ( .A(
        oc8051_memory_interface1_n19), .B(oc8051_memory_interface1_n20), .C(
        oc8051_memory_interface1_n21), .D(oc8051_memory_interface1_n71), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[6]) );
  INV_X1M_A12TS oc8051_memory_interface1_u48 ( .A(
        oc8051_memory_interface1_idat_cur_28_), .Y(
        oc8051_memory_interface1_n69) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u47 ( .A(
        oc8051_memory_interface1_n13), .B(oc8051_memory_interface1_n14), .C(
        oc8051_memory_interface1_n15), .D(oc8051_memory_interface1_n69), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[4]) );
  INV_X1M_A12TS oc8051_memory_interface1_u46 ( .A(
        oc8051_memory_interface1_idat_cur_27_), .Y(
        oc8051_memory_interface1_n68) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u45 ( .A(
        oc8051_memory_interface1_n10), .B(oc8051_memory_interface1_n11), .C(
        oc8051_memory_interface1_n12), .D(oc8051_memory_interface1_n68), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[3]) );
  INV_X1M_A12TS oc8051_memory_interface1_u44 ( .A(
        oc8051_memory_interface1_idat_cur_26_), .Y(
        oc8051_memory_interface1_n67) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u43 ( .A(
        oc8051_memory_interface1_n7), .B(oc8051_memory_interface1_n8), .C(
        oc8051_memory_interface1_n9), .D(oc8051_memory_interface1_n67), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[2]) );
  INV_X1M_A12TS oc8051_memory_interface1_u42 ( .A(
        oc8051_memory_interface1_idat_cur_29_), .Y(
        oc8051_memory_interface1_n70) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u41 ( .A(
        oc8051_memory_interface1_n16), .B(oc8051_memory_interface1_n17), .C(
        oc8051_memory_interface1_n18), .D(oc8051_memory_interface1_n70), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[5]) );
  INV_X1M_A12TS oc8051_memory_interface1_u40 ( .A(
        oc8051_memory_interface1_idat_cur_24_), .Y(
        oc8051_memory_interface1_n65) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u39 ( .A(
        oc8051_memory_interface1_n1), .B(oc8051_memory_interface1_n2), .C(
        oc8051_memory_interface1_n3), .D(oc8051_memory_interface1_n65), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[0]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u38 ( .A(
        oc8051_memory_interface1_n46), .B(
        oc8051_memory_interface1_idat_cur_23_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n48)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u37 ( .A(
        oc8051_memory_interface1_idat_old_15_), .B(
        oc8051_memory_interface1_idat_cur_15_), .C(
        oc8051_memory_interface1_idat_old_23_), .D(
        oc8051_memory_interface1_idat_cur_23_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n47)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u36 ( .A(
        oc8051_memory_interface1_n47), .B(oc8051_memory_interface1_n48), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[7]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u35 ( .A(
        oc8051_memory_interface1_n31), .B(
        oc8051_memory_interface1_idat_cur_18_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n33)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u34 ( .A(
        oc8051_memory_interface1_idat_old_10_), .B(
        oc8051_memory_interface1_idat_cur_10_), .C(
        oc8051_memory_interface1_idat_old_18_), .D(
        oc8051_memory_interface1_idat_cur_18_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n32)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u33 ( .A(
        oc8051_memory_interface1_n32), .B(oc8051_memory_interface1_n33), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[2]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u32 ( .A(
        oc8051_memory_interface1_n25), .B(
        oc8051_memory_interface1_idat_cur_16_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n27)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u31 ( .A(
        oc8051_memory_interface1_idat_old_8_), .B(
        oc8051_memory_interface1_idat_cur_8_), .C(
        oc8051_memory_interface1_idat_old_16_), .D(
        oc8051_memory_interface1_idat_cur_16_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n26)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u30 ( .A(
        oc8051_memory_interface1_n26), .B(oc8051_memory_interface1_n27), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[0]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u29 ( .A(
        oc8051_memory_interface1_n37), .B(
        oc8051_memory_interface1_idat_cur_20_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n39)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u28 ( .A(
        oc8051_memory_interface1_idat_old_12_), .B(
        oc8051_memory_interface1_idat_cur_12_), .C(
        oc8051_memory_interface1_idat_old_20_), .D(
        oc8051_memory_interface1_idat_cur_20_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n38)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u27 ( .A(
        oc8051_memory_interface1_n38), .B(oc8051_memory_interface1_n39), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[4]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u26 ( .A(
        oc8051_memory_interface1_n34), .B(
        oc8051_memory_interface1_idat_cur_19_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n36)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u25 ( .A(
        oc8051_memory_interface1_idat_old_11_), .B(
        oc8051_memory_interface1_idat_cur_11_), .C(
        oc8051_memory_interface1_idat_old_19_), .D(
        oc8051_memory_interface1_idat_cur_19_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n35)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u24 ( .A(
        oc8051_memory_interface1_n35), .B(oc8051_memory_interface1_n36), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[3]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u23 ( .A(
        oc8051_memory_interface1_n40), .B(
        oc8051_memory_interface1_idat_cur_21_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n42)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u22 ( .A(
        oc8051_memory_interface1_idat_old_13_), .B(
        oc8051_memory_interface1_idat_cur_13_), .C(
        oc8051_memory_interface1_idat_old_21_), .D(
        oc8051_memory_interface1_idat_cur_21_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n41)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u21 ( .A(
        oc8051_memory_interface1_n41), .B(oc8051_memory_interface1_n42), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[5]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u20 ( .A(
        oc8051_memory_interface1_n43), .B(
        oc8051_memory_interface1_idat_cur_22_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n45)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u19 ( .A(
        oc8051_memory_interface1_idat_old_14_), .B(
        oc8051_memory_interface1_idat_cur_14_), .C(
        oc8051_memory_interface1_idat_old_22_), .D(
        oc8051_memory_interface1_idat_cur_22_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n44)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u18 ( .A(
        oc8051_memory_interface1_n44), .B(oc8051_memory_interface1_n45), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[6]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u17 ( .A(
        oc8051_memory_interface1_n28), .B(
        oc8051_memory_interface1_idat_cur_17_), .S0(
        oc8051_memory_interface1_op_pos_2_), .Y(oc8051_memory_interface1_n30)
         );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u16 ( .A(
        oc8051_memory_interface1_idat_old_9_), .B(
        oc8051_memory_interface1_idat_cur_9_), .C(
        oc8051_memory_interface1_idat_old_17_), .D(
        oc8051_memory_interface1_idat_cur_17_), .S0(
        oc8051_memory_interface1_op_pos_2_), .S1(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n29)
         );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u15 ( .A(
        oc8051_memory_interface1_n29), .B(oc8051_memory_interface1_n30), .S0(
        oc8051_memory_interface1_op_pos_1_), .Y(
        oc8051_memory_interface1_op2[1]) );
  MXIT2_X0P7M_A12TS oc8051_memory_interface1_u14 ( .A(
        oc8051_memory_interface1_idat_cur_17_), .B(
        oc8051_memory_interface1_idat_cur_25_), .S0(
        oc8051_memory_interface1_op_pos_0_), .Y(oc8051_memory_interface1_n6)
         );
  INV_X1M_A12TS oc8051_memory_interface1_u13 ( .A(
        oc8051_memory_interface1_idat_cur_25_), .Y(
        oc8051_memory_interface1_n66) );
  MXIT4_X1M_A12TS oc8051_memory_interface1_u12 ( .A(
        oc8051_memory_interface1_n4), .B(oc8051_memory_interface1_n5), .C(
        oc8051_memory_interface1_n6), .D(oc8051_memory_interface1_n66), .S0(
        oc8051_memory_interface1_op_pos_1_), .S1(
        oc8051_memory_interface1_op_pos_2_), .Y(
        oc8051_memory_interface1_op3[1]) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u11 ( .A(
        oc8051_memory_interface1_n90), .B(oc8051_memory_interface1_n91), .Y(
        wr_addr[2]) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u10 ( .A(
        oc8051_memory_interface1_n92), .B(oc8051_memory_interface1_n93), .Y(
        wr_addr[1]) );
  NAND2_X1M_A12TS oc8051_memory_interface1_u9 ( .A(
        oc8051_memory_interface1_n94), .B(oc8051_memory_interface1_n95), .Y(
        wr_addr[0]) );
  NAND2_X0P5M_A12TS oc8051_memory_interface1_u8 ( .A(
        oc8051_memory_interface1_n134), .B(oc8051_memory_interface1_n167), .Y(
        oc8051_memory_interface1_n132) );
  OAI211_X1M_A12TS oc8051_memory_interface1_u7 ( .A0(
        oc8051_memory_interface1_n121), .A1(oc8051_memory_interface1_n104), 
        .B0(oc8051_memory_interface1_n122), .C0(oc8051_memory_interface1_n123), 
        .Y(rd_addr[2]) );
  NAND3_X2M_A12TS oc8051_memory_interface1_u6 ( .A(
        oc8051_memory_interface1_n124), .B(oc8051_memory_interface1_n125), .C(
        oc8051_memory_interface1_n126), .Y(rd_addr[1]) );
  OAI211_X2M_A12TS oc8051_memory_interface1_u5 ( .A0(
        oc8051_memory_interface1_n127), .A1(oc8051_memory_interface1_n104), 
        .B0(oc8051_memory_interface1_n128), .C0(oc8051_memory_interface1_n129), 
        .Y(rd_addr[0]) );
  INV_X1M_A12TS oc8051_memory_interface1_u4 ( .A(oc8051_memory_interface1_n194), .Y(oc8051_memory_interface1_n200) );
  NOR2_X2M_A12TS oc8051_memory_interface1_u3 ( .A(
        oc8051_memory_interface1_n200), .B(oc8051_memory_interface1_n187), .Y(
        oc8051_memory_interface1_n134) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_wr_r_reg ( .D(
        oc8051_memory_interface1_n5530), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_wr_r) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op_pos_reg_0_ ( .D(
        oc8051_memory_interface1_n492), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_op_pos_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op_pos_reg_2_ ( .D(
        oc8051_memory_interface1_n557), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_op_pos_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dstb_o_reg ( .D(
        oc8051_memory_interface1_n813), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_cyc_o) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dwe_o_reg ( .D(
        oc8051_memory_interface1_n1310), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_we_o) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op_pos_reg_1_ ( .D(
        oc8051_memory_interface1_n491), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_op_pos_1_) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_14_ ( .D(
        oc8051_memory_interface1_n476), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n392) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_9_ ( .D(
        oc8051_memory_interface1_n481), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n397) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_13_ ( .D(
        oc8051_memory_interface1_n477), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n393) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_11_ ( .D(
        oc8051_memory_interface1_n479), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n395) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_istb_t_reg ( .D(
        oc8051_memory_interface1_n583), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_istb_t) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_8_ ( .D(
        oc8051_memory_interface1_n482), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n398) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_15_ ( .D(
        oc8051_memory_interface1_n475), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n399) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_12_ ( .D(
        oc8051_memory_interface1_n478), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n394) );
  DFFRPQN_X1M_A12TS oc8051_memory_interface1_pc_reg_10_ ( .D(
        oc8051_memory_interface1_n480), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_memory_interface1_n396) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_16_ ( .D(
        oc8051_memory_interface1_n524), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_16_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_17_ ( .D(
        oc8051_memory_interface1_n522), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_17_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_18_ ( .D(
        oc8051_memory_interface1_n520), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_18_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_19_ ( .D(
        oc8051_memory_interface1_n518), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_19_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_20_ ( .D(
        oc8051_memory_interface1_n516), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_20_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_21_ ( .D(
        oc8051_memory_interface1_n514), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_21_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_22_ ( .D(
        oc8051_memory_interface1_n512), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_22_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_23_ ( .D(
        oc8051_memory_interface1_n510), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_23_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_8_ ( .D(
        oc8051_memory_interface1_n540), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_9_ ( .D(
        oc8051_memory_interface1_n538), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_10_ ( .D(
        oc8051_memory_interface1_n536), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_11_ ( .D(
        oc8051_memory_interface1_n534), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_12_ ( .D(
        oc8051_memory_interface1_n532), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_13_ ( .D(
        oc8051_memory_interface1_n530), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_14_ ( .D(
        oc8051_memory_interface1_n528), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_15_ ( .D(
        oc8051_memory_interface1_n526), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dack_ir_reg ( .D(wbd_ack_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_dack_ir) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_0_ ( .D(
        oc8051_memory_interface1_n796), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_1_ ( .D(
        oc8051_memory_interface1_n795), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_2_ ( .D(
        oc8051_memory_interface1_n794), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_3_ ( .D(
        oc8051_memory_interface1_n793), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_4_ ( .D(
        oc8051_memory_interface1_n792), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_5_ ( .D(
        oc8051_memory_interface1_n791), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_6_ ( .D(
        oc8051_memory_interface1_n790), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_7_ ( .D(
        oc8051_memory_interface1_n789), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_24_ ( .D(
        oc8051_memory_interface1_n508), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_24_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_25_ ( .D(
        oc8051_memory_interface1_n506), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_25_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_26_ ( .D(
        oc8051_memory_interface1_n504), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_26_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_27_ ( .D(
        oc8051_memory_interface1_n502), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_27_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_28_ ( .D(
        oc8051_memory_interface1_n500), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_28_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_29_ ( .D(
        oc8051_memory_interface1_n498), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_29_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_30_ ( .D(
        oc8051_memory_interface1_n496), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_30_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_cur_reg_31_ ( .D(
        oc8051_memory_interface1_n494), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_cur_31_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_24_ ( .D(
        oc8051_memory_interface1_n507), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_24_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_25_ ( .D(
        oc8051_memory_interface1_n505), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_25_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_26_ ( .D(
        oc8051_memory_interface1_n503), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_26_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_27_ ( .D(
        oc8051_memory_interface1_n501), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_27_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_28_ ( .D(
        oc8051_memory_interface1_n499), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_28_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_29_ ( .D(
        oc8051_memory_interface1_n497), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_29_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_30_ ( .D(
        oc8051_memory_interface1_n495), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_30_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_31_ ( .D(
        oc8051_memory_interface1_n493), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_31_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_11_ ( .D(
        oc8051_memory_interface1_n463), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_8_ ( .D(
        oc8051_memory_interface1_n539), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_9_ ( .D(
        oc8051_memory_interface1_n537), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_10_ ( .D(
        oc8051_memory_interface1_n535), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_11_ ( .D(
        oc8051_memory_interface1_n533), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_12_ ( .D(
        oc8051_memory_interface1_n531), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_13_ ( .D(
        oc8051_memory_interface1_n529), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_14_ ( .D(
        oc8051_memory_interface1_n527), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_15_ ( .D(
        oc8051_memory_interface1_n525), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_16_ ( .D(
        oc8051_memory_interface1_n523), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_16_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_17_ ( .D(
        oc8051_memory_interface1_n521), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_17_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_18_ ( .D(
        oc8051_memory_interface1_n519), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_18_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_19_ ( .D(
        oc8051_memory_interface1_n517), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_19_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_20_ ( .D(
        oc8051_memory_interface1_n515), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_20_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_21_ ( .D(
        oc8051_memory_interface1_n513), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_21_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_22_ ( .D(
        oc8051_memory_interface1_n511), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_22_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_23_ ( .D(
        oc8051_memory_interface1_n509), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_23_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_8_ ( .D(
        oc8051_memory_interface1_n466), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_4_ ( .D(
        oc8051_memory_interface1_n470), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_7_ ( .D(
        oc8051_memory_interface1_n467), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_3_ ( .D(
        oc8051_memory_interface1_n471), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_0_ ( .D(
        oc8051_memory_interface1_n555), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_1_ ( .D(
        oc8051_memory_interface1_n553), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_2_ ( .D(
        oc8051_memory_interface1_n551), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_3_ ( .D(
        oc8051_memory_interface1_n549), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_4_ ( .D(
        oc8051_memory_interface1_n547), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_5_ ( .D(
        oc8051_memory_interface1_n545), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_6_ ( .D(
        oc8051_memory_interface1_n543), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_idat_old_reg_7_ ( .D(
        oc8051_memory_interface1_n541), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_idat_old_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_1_ ( .D(
        oc8051_memory_interface1_n473), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_2_ ( .D(
        oc8051_memory_interface1_n472), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_12_ ( .D(
        oc8051_memory_interface1_n462), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_14_ ( .D(
        oc8051_memory_interface1_n460), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_6_ ( .D(
        oc8051_memory_interface1_n468), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_5_ ( .D(
        oc8051_memory_interface1_n469), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_1_ ( .D(
        oc8051_memory_interface1_n489), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[1])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_7_ ( .D(
        oc8051_memory_interface1_n483), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[7])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_15_ ( .D(
        oc8051_memory_interface1_n459), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_wr_r2_reg ( .D(
        oc8051_memory_interface1_pc_wr_r), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_wr_r2) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_5_ ( .D(
        oc8051_memory_interface1_n485), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[5])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_10_ ( .D(
        oc8051_memory_interface1_n464), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_ack_t_reg ( .D(
        oc8051_memory_interface1_n558), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_ack_t) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_0_ ( .D(
        oc8051_memory_interface1_n490), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[0])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_9_ ( .D(
        oc8051_memory_interface1_n465), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_4_ ( .D(
        oc8051_memory_interface1_n486), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[4])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_3_ ( .D(
        oc8051_memory_interface1_n487), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[3])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_2_ ( .D(
        oc8051_memory_interface1_n488), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[2])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imem_wait_reg ( .D(
        oc8051_memory_interface1_n584), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_imem_wait) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_0_ ( .D(
        oc8051_memory_interface1_n474), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_0_ ( .D(
        oc8051_memory_interface1_n797), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_2_ ( .D(
        oc8051_memory_interface1_n799), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_3_ ( .D(
        oc8051_memory_interface1_n800), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_5_ ( .D(
        oc8051_memory_interface1_n802), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_6_ ( .D(
        oc8051_memory_interface1_n803), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_7_ ( .D(
        oc8051_memory_interface1_n804), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_buf_reg_13_ ( .D(
        oc8051_memory_interface1_n461), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_pc_buf_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_pc_reg_6_ ( .D(
        oc8051_memory_interface1_n484), .CK(wb_clk_i), .R(wb_rst_i), .Q(pc[6])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_7_ ( .D(
        oc8051_memory_interface1_n447), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_12_ ( .D(
        oc8051_memory_interface1_n452), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_12_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_3_ ( .D(
        oc8051_memory_interface1_n443), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_4_ ( .D(
        oc8051_memory_interface1_n444), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_5_ ( .D(
        oc8051_memory_interface1_n445), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_6_ ( .D(
        oc8051_memory_interface1_n446), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_8_ ( .D(
        oc8051_memory_interface1_n448), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_8_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_9_ ( .D(
        oc8051_memory_interface1_n449), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_9_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_10_ ( .D(
        oc8051_memory_interface1_n450), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_10_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_11_ ( .D(
        oc8051_memory_interface1_n451), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_11_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_13_ ( .D(
        oc8051_memory_interface1_n453), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_13_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_14_ ( .D(
        oc8051_memory_interface1_n454), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_14_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_15_ ( .D(
        oc8051_memory_interface1_n455), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_15_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdone_reg ( .D(
        oc8051_memory_interface1_istb_t), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdone) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_0_ ( .D(
        oc8051_memory_interface1_n416), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_2_ ( .D(
        oc8051_memory_interface1_n418), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_3_ ( .D(
        oc8051_memory_interface1_n419), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_5_ ( .D(
        oc8051_memory_interface1_n421), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_6_ ( .D(
        oc8051_memory_interface1_n422), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_7_ ( .D(
        oc8051_memory_interface1_n423), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_1_ ( .D(
        oc8051_memory_interface1_n798), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_cdata_reg_4_ ( .D(
        oc8051_memory_interface1_n801), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_cdata_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_0_ ( .D(
        oc8051_memory_interface1_n424), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_1_ ( .D(
        oc8051_memory_interface1_n425), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_2_ ( .D(
        oc8051_memory_interface1_n426), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_3_ ( .D(
        oc8051_memory_interface1_n427), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_3_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_4_ ( .D(
        oc8051_memory_interface1_n428), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_5_ ( .D(
        oc8051_memory_interface1_n429), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_5_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_6_ ( .D(
        oc8051_memory_interface1_n430), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_6_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_vec_buff_reg_7_ ( .D(
        oc8051_memory_interface1_n431), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_vec_buff_7_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_1_ ( .D(
        oc8051_memory_interface1_n417), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_ir_reg_4_ ( .D(
        oc8051_memory_interface1_n420), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_ddat_ir_4_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dmem_wait_reg ( .D(
        oc8051_memory_interface1_n813), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_dmem_wait) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_reti_reg ( .D(
        oc8051_memory_interface1_n2000), .CK(wb_clk_i), .R(wb_rst_i), .Q(reti)
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_ack_reg ( .D(
        oc8051_memory_interface1_n3720), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        int_ack) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_0_ ( .D(
        oc8051_memory_interface1_n440), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_0_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_1_ ( .D(
        oc8051_memory_interface1_n441), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_1_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_iadr_t_reg_2_ ( .D(
        oc8051_memory_interface1_n442), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_iadr_t_2_) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_7_ ( .D(op3_n[7]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[7])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_0_ ( .D(op3_n[0]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[0])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_1_ ( .D(op3_n[1]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[1])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_2_ ( .D(op3_n[2]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[2])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_3_ ( .D(op3_n[3]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[3])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_4_ ( .D(op3_n[4]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[4])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_5_ ( .D(op3_n[5]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[5])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op3_buff_reg_6_ ( .D(op3_n[6]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op3_buff[6])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rd_ind_reg ( .D(
        oc8051_memory_interface1_n830), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_rd_ind) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_4_ ( .D(op3_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_5_ ( .D(op3_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_6_ ( .D(op3_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_7_ ( .D(op3_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_5_ ( .D(op2_n[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_6_ ( .D(op2_n[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_7_ ( .D(op2_n[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_0_ ( .D(ri[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_1_ ( .D(ri[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_2_ ( .D(ri[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_3_ ( .D(ri[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_0_ ( .D(op2_n[0]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[0])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_1_ ( .D(op2_n[1]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[1])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_2_ ( .D(op2_n[2]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[2])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_3_ ( .D(op2_n[3]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[3])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_4_ ( .D(op2_n[4]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[4])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_5_ ( .D(op2_n[5]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[5])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_6_ ( .D(op2_n[6]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[6])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_5_ ( .D(ri[5]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_6_ ( .D(ri[6]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_7_ ( .D(ri[7]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_0_ ( .D(op1_cur[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_1_ ( .D(op1_cur[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_2_ ( .D(op1_cur[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_3_ ( .D(bank_sel[0]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ri_r_reg_4_ ( .D(ri[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_ri_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_0_ ( .D(op2_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_1_ ( .D(op2_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_2_ ( .D(op2_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_3_ ( .D(op2_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rn_r_reg_4_ ( .D(bank_sel[1]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rn_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_0_ ( .D(op3_n[0]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_1_ ( .D(op3_n[1]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_2_ ( .D(op3_n[2]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm2_r_reg_3_ ( .D(op3_n[3]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm2_r[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_imm_r_reg_4_ ( .D(op2_n[4]), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_imm_r[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_rd_addr_r_reg ( .D(rd_addr[7]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_rd_addr_r) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_int_ack_buff_reg ( .D(
        oc8051_memory_interface1_int_ack_t), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_memory_interface1_int_ack_buff) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_op2_buff_reg_7_ ( .D(op2_n[7]), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_memory_interface1_op2_buff[7])
         );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_8_ ( .D(
        oc8051_memory_interface1_n567), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[8]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_9_ ( .D(
        oc8051_memory_interface1_n568), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[9]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_10_ ( .D(
        oc8051_memory_interface1_n569), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[10]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_11_ ( .D(
        oc8051_memory_interface1_n570), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[11]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_12_ ( .D(
        oc8051_memory_interface1_n571), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[12]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_13_ ( .D(
        oc8051_memory_interface1_n572), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[13]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_14_ ( .D(
        oc8051_memory_interface1_n573), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[14]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_15_ ( .D(
        oc8051_memory_interface1_n574), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[15]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_0_ ( .D(
        oc8051_memory_interface1_n575), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_1_ ( .D(
        oc8051_memory_interface1_n576), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_2_ ( .D(
        oc8051_memory_interface1_n577), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_3_ ( .D(
        oc8051_memory_interface1_n578), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_4_ ( .D(
        oc8051_memory_interface1_n579), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_5_ ( .D(
        oc8051_memory_interface1_n580), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_6_ ( .D(
        oc8051_memory_interface1_n581), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_ddat_o_reg_7_ ( .D(
        oc8051_memory_interface1_n582), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_dat_o[7]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_0_ ( .D(
        oc8051_memory_interface1_n559), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[0]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_1_ ( .D(
        oc8051_memory_interface1_n560), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[1]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_2_ ( .D(
        oc8051_memory_interface1_n561), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[2]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_3_ ( .D(
        oc8051_memory_interface1_n562), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[3]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_4_ ( .D(
        oc8051_memory_interface1_n563), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[4]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_5_ ( .D(
        oc8051_memory_interface1_n564), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[5]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_6_ ( .D(
        oc8051_memory_interface1_n565), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[6]) );
  DFFRPQ_X1M_A12TS oc8051_memory_interface1_dadr_ot_reg_7_ ( .D(
        oc8051_memory_interface1_n566), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        wbd_adr_o[7]) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u279 ( .A(rd_addr[3]), .B(rd_addr[6]), .Y(
        oc8051_sfr1_n219) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u278 ( .A(rd_addr[2]), .B(rd_addr[5]), .C(
        rd_addr[4]), .Y(oc8051_sfr1_n257) );
  AND4_X0P5M_A12TS oc8051_sfr1_u277 ( .A(wr_sfr[1]), .B(wr_sfr[0]), .C(
        oc8051_sfr1_n231), .D(oc8051_sfr1_n174), .Y(oc8051_sfr1_n35) );
  INV_X0P5B_A12TS oc8051_sfr1_u276 ( .A(rd_addr[2]), .Y(oc8051_sfr1_n172) );
  INV_X0P5B_A12TS oc8051_sfr1_u275 ( .A(rd_addr[3]), .Y(oc8051_sfr1_n183) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u274 ( .A(oc8051_sfr1_n174), .B(
        oc8051_sfr1_n185), .C(oc8051_sfr1_n172), .D(oc8051_sfr1_n183), .Y(
        oc8051_sfr1_n227) );
  INV_X0P5B_A12TS oc8051_sfr1_u273 ( .A(rd_addr[4]), .Y(oc8051_sfr1_n182) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u272 ( .A(oc8051_sfr1_n182), .B(rd_addr[5]), 
        .Y(oc8051_sfr1_n181) );
  INV_X0P5B_A12TS oc8051_sfr1_u271 ( .A(rd_addr[6]), .Y(oc8051_sfr1_n168) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u270 ( .AN(oc8051_sfr1_n181), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n42) );
  OAI211_X0P5M_A12TS oc8051_sfr1_u269 ( .A0(psw_set[1]), .A1(psw_set[0]), .B0(
        rd_addr[7]), .C0(oc8051_sfr1_n42), .Y(oc8051_sfr1_n228) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u268 ( .A(oc8051_sfr1_n174), .B(
        oc8051_sfr1_n172), .Y(oc8051_sfr1_n170) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u267 ( .A(wr_addr[3]), .B(oc8051_sfr1_n183), 
        .Y(oc8051_sfr1_n251) );
  INV_X0P5B_A12TS oc8051_sfr1_u266 ( .A(wr_addr[6]), .Y(oc8051_sfr1_n203) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u265 ( .A(oc8051_sfr1_n203), .B(rd_addr[6]), 
        .Y(oc8051_sfr1_n252) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u264 ( .A(wr_addr[4]), .B(rd_addr[4]), .Y(
        oc8051_sfr1_n255) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u263 ( .A(wr_addr[5]), .B(rd_addr[5]), .Y(
        oc8051_sfr1_n256) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u262 ( .A(oc8051_sfr1_n255), .B(
        oc8051_sfr1_n256), .Y(oc8051_sfr1_n253) );
  INV_X0P5B_A12TS oc8051_sfr1_u261 ( .A(wr_addr[7]), .Y(oc8051_sfr1_n250) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u260 ( .A(rd_addr[7]), .B(oc8051_sfr1_n250), 
        .Y(oc8051_sfr1_n254) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u259 ( .A(oc8051_sfr1_n251), .B(
        oc8051_sfr1_n252), .C(oc8051_sfr1_n253), .D(oc8051_sfr1_n254), .Y(
        oc8051_sfr1_n249) );
  AOI211_X0P5M_A12TS oc8051_sfr1_u258 ( .A0(oc8051_sfr1_n170), .A1(rd_addr[1]), 
        .B0(oc8051_sfr1_n249), .C0(oc8051_sfr1_n250), .Y(oc8051_sfr1_n236) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u257 ( .A(wr_addr[0]), .B(oc8051_sfr1_n174), 
        .Y(oc8051_sfr1_n246) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u256 ( .A(wr_addr[2]), .B(oc8051_sfr1_n172), 
        .Y(oc8051_sfr1_n247) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u255 ( .A(wr_addr[1]), .B(oc8051_sfr1_n185), 
        .Y(oc8051_sfr1_n248) );
  INV_X0P5B_A12TS oc8051_sfr1_u254 ( .A(oc8051_sfr1_n249), .Y(oc8051_sfr1_n210) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u253 ( .A(oc8051_sfr1_n246), .B(
        oc8051_sfr1_n247), .C(oc8051_sfr1_n248), .D(oc8051_sfr1_n210), .Y(
        oc8051_sfr1_n214) );
  INV_X0P5B_A12TS oc8051_sfr1_u252 ( .A(oc8051_sfr1_n214), .Y(oc8051_sfr1_n245) );
  INV_X0P5B_A12TS oc8051_sfr1_u251 ( .A(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_n200) );
  AND4_X0P5M_A12TS oc8051_sfr1_u250 ( .A(oc8051_sfr1_n245), .B(n_5_net_), .C(
        wr_addr[7]), .D(oc8051_sfr1_n200), .Y(oc8051_sfr1_n187) );
  AOI31_X0P5M_A12TS oc8051_sfr1_u249 ( .A0(oc8051_sfr1_wr_bit_r), .A1(n_5_net_), .A2(oc8051_sfr1_n236), .B0(oc8051_sfr1_n187), .Y(oc8051_sfr1_n229) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u248 ( .AN(wr_sfr[1]), .B(wr_sfr[0]), .Y(
        oc8051_sfr1_n198) );
  INV_X0P5B_A12TS oc8051_sfr1_u247 ( .A(rd_addr[5]), .Y(oc8051_sfr1_n186) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u246 ( .A(oc8051_sfr1_n186), .B(rd_addr[4]), 
        .C(oc8051_sfr1_n168), .Y(oc8051_sfr1_n40) );
  AND3_X0P5M_A12TS oc8051_sfr1_u245 ( .A(rd_addr[7]), .B(oc8051_sfr1_n183), 
        .C(oc8051_sfr1_n40), .Y(oc8051_sfr1_n235) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u244 ( .AN(wr_sfr[0]), .B(wr_sfr[1]), .Y(
        oc8051_sfr1_n197) );
  AND2_X0P5M_A12TS oc8051_sfr1_u243 ( .A(oc8051_sfr1_n197), .B(
        oc8051_sfr1_n235), .Y(oc8051_sfr1_n209) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_u242 ( .A0(oc8051_sfr1_n198), .A1(
        oc8051_sfr1_n235), .B0(oc8051_sfr1_n209), .C0(oc8051_sfr1_n174), .Y(
        oc8051_sfr1_n234) );
  INV_X0P5B_A12TS oc8051_sfr1_u241 ( .A(oc8051_sfr1_n234), .Y(oc8051_sfr1_n232) );
  AOI32_X0P5M_A12TS oc8051_sfr1_u240 ( .A0(wr_sfr[0]), .A1(oc8051_sfr1_n231), 
        .A2(wr_sfr[1]), .B0(oc8051_sfr1_n232), .B1(oc8051_sfr1_n233), .Y(
        oc8051_sfr1_n230) );
  OA211_X0P5M_A12TS oc8051_sfr1_u239 ( .A0(oc8051_sfr1_n227), .A1(
        oc8051_sfr1_n228), .B0(oc8051_sfr1_n229), .C0(oc8051_sfr1_n230), .Y(
        oc8051_sfr1_n226) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u238 ( .A(wait_data), .B(oc8051_sfr1_n35), .C(
        oc8051_sfr1_n226), .Y(oc8051_sfr1_n1020) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u237 ( .A(rd_addr[3]), .B(rd_addr[5]), .Y(
        oc8051_sfr1_n175) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u236 ( .A(oc8051_sfr1_n1350), .B(
        oc8051_sfr1_n1340), .S0(rd_addr[4]), .Y(oc8051_sfr1_n223) );
  NAND3_X0P5A_A12TS oc8051_sfr1_u235 ( .A(rd_addr[3]), .B(rd_addr[6]), .C(
        oc8051_sfr1_n1380), .Y(oc8051_sfr1_n224) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u234 ( .A(oc8051_sfr1_n186), .B(
        oc8051_sfr1_n182), .Y(oc8051_sfr1_n184) );
  NAND3_X0P5A_A12TS oc8051_sfr1_u233 ( .A(oc8051_sfr1_n184), .B(
        oc8051_sfr1_n219), .C(oc8051_sfr1_n1320), .Y(oc8051_sfr1_n225) );
  OAI211_X0P5M_A12TS oc8051_sfr1_u232 ( .A0(oc8051_sfr1_n175), .A1(
        oc8051_sfr1_n223), .B0(oc8051_sfr1_n224), .C0(oc8051_sfr1_n225), .Y(
        oc8051_sfr1_n215) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u231 ( .A(oc8051_sfr1_n183), .B(rd_addr[6]), 
        .Y(oc8051_sfr1_n173) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u230 ( .A0(oc8051_sfr1_n1360), .A1(
        oc8051_sfr1_n173), .B0(oc8051_sfr1_n1290), .B1(oc8051_sfr1_n183), .Y(
        oc8051_sfr1_n221) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u229 ( .A(oc8051_sfr1_n1370), .B(rd_addr[3]), 
        .Y(oc8051_sfr1_n222) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u228 ( .A(oc8051_sfr1_n221), .B(
        oc8051_sfr1_n222), .S0(rd_addr[4]), .Y(oc8051_sfr1_n220) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u227 ( .AN(oc8051_sfr1_n184), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n55) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u226 ( .A0(oc8051_sfr1_n220), .A1(
        oc8051_sfr1_n186), .B0(oc8051_sfr1_n1330), .B1(oc8051_sfr1_n55), .Y(
        oc8051_sfr1_n216) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u225 ( .A0(oc8051_sfr1_n1280), .A1(
        oc8051_sfr1_n42), .B0(oc8051_sfr1_n1270), .B1(oc8051_sfr1_n40), .Y(
        oc8051_sfr1_n217) );
  AND2_X0P5M_A12TS oc8051_sfr1_u224 ( .A(oc8051_sfr1_n181), .B(
        oc8051_sfr1_n219), .Y(oc8051_sfr1_n53) );
  AND3_X0P5M_A12TS oc8051_sfr1_u223 ( .A(oc8051_sfr1_n219), .B(
        oc8051_sfr1_n182), .C(rd_addr[5]), .Y(oc8051_sfr1_n41) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u222 ( .A0(oc8051_sfr1_n1300), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_n1310), .B1(oc8051_sfr1_n41), .Y(
        oc8051_sfr1_n218) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u221 ( .AN(oc8051_sfr1_n215), .B(
        oc8051_sfr1_n216), .C(oc8051_sfr1_n217), .D(oc8051_sfr1_n218), .Y(
        oc8051_sfr1_n212) );
  INV_X0P5B_A12TS oc8051_sfr1_u220 ( .A(n_5_net_), .Y(oc8051_sfr1_n204) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u219 ( .A(oc8051_sfr1_n200), .B(
        oc8051_sfr1_n214), .C(oc8051_sfr1_n204), .Y(oc8051_sfr1_n213) );
  AOI31_X0P5M_A12TS oc8051_sfr1_u218 ( .A0(wr_addr[2]), .A1(wr_addr[1]), .A2(
        wr_addr[0]), .B0(oc8051_sfr1_wr_bit_r), .Y(oc8051_sfr1_n211) );
  AND3_X0P5M_A12TS oc8051_sfr1_u217 ( .A(n_5_net_), .B(oc8051_sfr1_n210), .C(
        oc8051_sfr1_n211), .Y(oc8051_sfr1_n191) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u216 ( .A(oc8051_sfr1_n209), .B(
        oc8051_sfr1_n191), .Y(oc8051_sfr1_n208) );
  XOR2_X0P5M_A12TS oc8051_sfr1_u215 ( .A(oc8051_sfr1_prescaler_1_), .B(
        oc8051_sfr1_prescaler_0_), .Y(oc8051_sfr1_n1500) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u214 ( .A(oc8051_sfr1_prescaler_1_), .B(
        oc8051_sfr1_prescaler_0_), .Y(oc8051_sfr1_n31) );
  INV_X0P5B_A12TS oc8051_sfr1_u213 ( .A(oc8051_sfr1_n31), .Y(oc8051_sfr1_n205)
         );
  INV_X0P5B_A12TS oc8051_sfr1_u212 ( .A(oc8051_sfr1_prescaler_3_), .Y(
        oc8051_sfr1_n30) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u211 ( .A(oc8051_sfr1_n205), .B(
        oc8051_sfr1_n30), .Y(oc8051_sfr1_n206) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u210 ( .A(oc8051_sfr1_n206), .B(
        oc8051_sfr1_n205), .S0(oc8051_sfr1_prescaler_2_), .Y(oc8051_sfr1_n1510) );
  INV_X0P5B_A12TS oc8051_sfr1_u209 ( .A(oc8051_sfr1_prescaler_2_), .Y(
        oc8051_sfr1_n207) );
  OAI22_X0P5M_A12TS oc8051_sfr1_u208 ( .A0(oc8051_sfr1_n205), .A1(
        oc8051_sfr1_n30), .B0(oc8051_sfr1_n206), .B1(oc8051_sfr1_n207), .Y(
        oc8051_sfr1_n1520) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u207 ( .A(comp_sel[1]), .B(wr_addr[5]), .S0(
        wr_addr[4]), .Y(oc8051_sfr1_n202) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u206 ( .A(oc8051_sfr1_n202), .B(
        oc8051_sfr1_n203), .C(oc8051_sfr1_n204), .Y(oc8051_sfr1_n192) );
  OR3_X0P5M_A12TS oc8051_sfr1_u205 ( .A(wr_addr[1]), .B(wr_addr[2]), .C(
        wr_addr[0]), .Y(oc8051_sfr1_n199) );
  OAI21_X0P5M_A12TS oc8051_sfr1_u204 ( .A0(comp_sel[1]), .A1(wr_addr[5]), .B0(
        wr_addr[7]), .Y(oc8051_sfr1_n201) );
  AOI211_X0P5M_A12TS oc8051_sfr1_u203 ( .A0(oc8051_sfr1_n199), .A1(
        oc8051_sfr1_n200), .B0(oc8051_sfr1_n201), .C0(wr_addr[3]), .Y(
        oc8051_sfr1_n193) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u202 ( .A(oc8051_sfr1_n197), .B(
        oc8051_sfr1_n198), .Y(oc8051_sfr1_n195) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u201 ( .A(psw_set[1]), .B(psw_set[0]), .Y(
        oc8051_sfr1_n196) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u200 ( .A(oc8051_sfr1_n195), .B(
        oc8051_sfr1_n196), .S0(comp_sel[1]), .Y(oc8051_sfr1_n194) );
  AOI21_X0P5M_A12TS oc8051_sfr1_u199 ( .A0(oc8051_sfr1_n192), .A1(
        oc8051_sfr1_n193), .B0(oc8051_sfr1_n194), .Y(oc8051_sfr1_n189) );
  NAND2_X0P5A_A12TS oc8051_sfr1_u198 ( .A(comp_sel[1]), .B(oc8051_sfr1_n191), 
        .Y(oc8051_sfr1_n190) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u197 ( .A(oc8051_sfr1_n189), .B(
        oc8051_sfr1_n190), .S0(comp_sel[0]), .Y(oc8051_sfr1_n188) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u196 ( .A(oc8051_sfr1_n187), .B(
        oc8051_sfr1_n188), .Y(comp_wait) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u195 ( .A(oc8051_sfr1_n35), .B(
        oc8051_sfr1_n1020), .Y(oc8051_sfr1_n33) );
  NOR2_X0P5A_A12TS oc8051_sfr1_u194 ( .A(oc8051_sfr1_n172), .B(
        oc8051_sfr1_n186), .Y(oc8051_sfr1_n71) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u193 ( .A(rd_addr[0]), .B(rd_addr[6]), .C(
        oc8051_sfr1_n172), .Y(oc8051_sfr1_n72) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u192 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(
        oc8051_sfr1_n183), .Y(oc8051_sfr1_n169) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u191 ( .A0(oc8051_sfr1_ip_7_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[7]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[7]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n176) );
  AND2_X0P5M_A12TS oc8051_sfr1_u190 ( .A(oc8051_sfr1_n173), .B(
        oc8051_sfr1_n167), .Y(oc8051_sfr1_n68) );
  AND4_X0P5M_A12TS oc8051_sfr1_u189 ( .A(oc8051_sfr1_n174), .B(
        oc8051_sfr1_n185), .C(oc8051_sfr1_n182), .D(oc8051_sfr1_n186), .Y(
        oc8051_sfr1_n171) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u188 ( .AN(oc8051_sfr1_n171), .B(rd_addr[3]), 
        .Y(oc8051_sfr1_n69) );
  AND2_X0P5M_A12TS oc8051_sfr1_u187 ( .A(oc8051_sfr1_n173), .B(
        oc8051_sfr1_n170), .Y(oc8051_sfr1_n70) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u186 ( .A0(oc8051_sfr1_tl0[7]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_7_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[7]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n177) );
  AND3_X0P5M_A12TS oc8051_sfr1_u185 ( .A(oc8051_sfr1_n172), .B(
        oc8051_sfr1_n168), .C(oc8051_sfr1_n184), .Y(oc8051_sfr1_n65) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u184 ( .A(rd_addr[1]), .B(rd_addr[3]), .C(
        oc8051_sfr1_n174), .Y(oc8051_sfr1_n66) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u183 ( .A0(oc8051_sfr1_p3_data_7_), .A1(
        oc8051_sfr1_n65), .B0(sp[7]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[7]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n178) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u182 ( .AN(oc8051_sfr1_n167), .B(rd_addr[3]), 
        .Y(oc8051_sfr1_n60) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u181 ( .A(oc8051_sfr1_n182), .B(rd_addr[0]), 
        .C(oc8051_sfr1_n183), .Y(oc8051_sfr1_n61) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u180 ( .AN(oc8051_sfr1_n181), .B(
        oc8051_sfr1_n174), .Y(oc8051_sfr1_n63) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u179 ( .A(rd_addr[3]), .B(rd_addr[5]), .C(
        oc8051_sfr1_n172), .Y(oc8051_sfr1_n64) );
  AO22_X0P5M_A12TS oc8051_sfr1_u178 ( .A0(oc8051_sfr1_sbuf[7]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[7]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n180) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u177 ( .A0(dptr_lo[7]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_7_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n180), 
        .Y(oc8051_sfr1_n179) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u176 ( .A(oc8051_sfr1_n176), .B(
        oc8051_sfr1_n177), .C(oc8051_sfr1_n178), .D(oc8051_sfr1_n179), .Y(
        oc8051_sfr1_n160) );
  INV_X0P5B_A12TS oc8051_sfr1_u175 ( .A(oc8051_sfr1_n175), .Y(oc8051_sfr1_n54)
         );
  AOI222_X0P5M_A12TS oc8051_sfr1_u174 ( .A0(oc8051_sfr1_p1_data_7_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_7_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_7_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n161) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u173 ( .A(oc8051_sfr1_n168), .B(rd_addr[2]), 
        .C(oc8051_sfr1_n174), .Y(oc8051_sfr1_n51) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u172 ( .A(oc8051_sfr1_n168), .B(rd_addr[0]), 
        .C(oc8051_sfr1_n172), .Y(oc8051_sfr1_n52) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u171 ( .A0(oc8051_sfr1_rcap2h[7]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[7]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n164) );
  AND3_X0P5M_A12TS oc8051_sfr1_u170 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(
        oc8051_sfr1_n173), .Y(oc8051_sfr1_n49) );
  AND3_X0P5M_A12TS oc8051_sfr1_u169 ( .A(oc8051_sfr1_n171), .B(
        oc8051_sfr1_n172), .C(oc8051_sfr1_n173), .Y(oc8051_sfr1_n50) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u168 ( .A0(oc8051_sfr1_tl1[7]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_7_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n165) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u167 ( .AN(oc8051_sfr1_n170), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n46) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u166 ( .AN(oc8051_sfr1_n169), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n47) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_u165 ( .AN(oc8051_sfr1_n167), .B(
        oc8051_sfr1_n168), .Y(oc8051_sfr1_n48) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u164 ( .A0(oc8051_sfr1_th2[7]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_7_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[7]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n166)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u163 ( .A(oc8051_sfr1_n164), .B(
        oc8051_sfr1_n165), .C(oc8051_sfr1_n166), .Y(oc8051_sfr1_n162) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u162 ( .A0(acc[7]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_7_), .B1(oc8051_sfr1_n41), .C0(cy), .C1(
        oc8051_sfr1_n42), .Y(oc8051_sfr1_n163) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u161 ( .AN(oc8051_sfr1_n160), .B(
        oc8051_sfr1_n161), .C(oc8051_sfr1_n162), .D(oc8051_sfr1_n163), .Y(
        oc8051_sfr1_n159) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u160 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n159), .B0(des_acc[7]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n158) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u159 ( .B0(sfr_out[7]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n158), .Y(oc8051_sfr1_n237) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u158 ( .A0(oc8051_sfr1_ip_6_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[6]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[6]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n153) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u157 ( .A0(oc8051_sfr1_tl0[6]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_6_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[6]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n154) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u156 ( .A0(oc8051_sfr1_p3_data_6_), .A1(
        oc8051_sfr1_n65), .B0(sp[6]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[6]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n155) );
  AO22_X0P5M_A12TS oc8051_sfr1_u155 ( .A0(oc8051_sfr1_sbuf[6]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[6]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n157) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u154 ( .A0(dptr_lo[6]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_6_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n157), 
        .Y(oc8051_sfr1_n156) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u153 ( .A(oc8051_sfr1_n153), .B(
        oc8051_sfr1_n154), .C(oc8051_sfr1_n155), .D(oc8051_sfr1_n156), .Y(
        oc8051_sfr1_n146) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u152 ( .A0(oc8051_sfr1_p1_data_6_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_6_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_6_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n147) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u151 ( .A0(oc8051_sfr1_rcap2h[6]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[6]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n150) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u150 ( .A0(oc8051_sfr1_tl1[6]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tr1), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n151) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u149 ( .A0(oc8051_sfr1_th2[6]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_6_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[6]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n152)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u148 ( .A(oc8051_sfr1_n150), .B(
        oc8051_sfr1_n151), .C(oc8051_sfr1_n152), .Y(oc8051_sfr1_n148) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u147 ( .A0(acc[6]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_6_), .B1(oc8051_sfr1_n41), .C0(srcac), .C1(
        oc8051_sfr1_n42), .Y(oc8051_sfr1_n149) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u146 ( .AN(oc8051_sfr1_n146), .B(
        oc8051_sfr1_n147), .C(oc8051_sfr1_n148), .D(oc8051_sfr1_n149), .Y(
        oc8051_sfr1_n145) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u145 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n145), .B0(des_acc[6]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n144) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u144 ( .B0(sfr_out[6]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n144), .Y(oc8051_sfr1_n238) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u143 ( .A0(oc8051_sfr1_ip_5_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[5]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[5]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n139) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u142 ( .A0(oc8051_sfr1_tl0[5]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_5_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[5]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n140) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u141 ( .A0(oc8051_sfr1_p3_data_5_), .A1(
        oc8051_sfr1_n65), .B0(sp[5]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[5]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n141) );
  AO22_X0P5M_A12TS oc8051_sfr1_u140 ( .A0(oc8051_sfr1_sbuf[5]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[5]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n143) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u139 ( .A0(dptr_lo[5]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_5_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n143), 
        .Y(oc8051_sfr1_n142) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u138 ( .A(oc8051_sfr1_n139), .B(
        oc8051_sfr1_n140), .C(oc8051_sfr1_n141), .D(oc8051_sfr1_n142), .Y(
        oc8051_sfr1_n132) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u137 ( .A0(oc8051_sfr1_p1_data_5_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_5_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_5_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n133) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u136 ( .A0(oc8051_sfr1_rcap2h[5]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[5]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n136) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u135 ( .A0(oc8051_sfr1_tl1[5]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_5_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n137) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u134 ( .A0(oc8051_sfr1_th2[5]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_rclk), .B1(oc8051_sfr1_n47), .C0(
        oc8051_sfr1_rcap2l[5]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n138) );
  AND3_X0P5M_A12TS oc8051_sfr1_u133 ( .A(oc8051_sfr1_n136), .B(
        oc8051_sfr1_n137), .C(oc8051_sfr1_n138), .Y(oc8051_sfr1_n134) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u132 ( .A0(acc[5]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_5_), .B1(oc8051_sfr1_n41), .C0(
        oc8051_sfr1_psw_5_), .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n135) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u131 ( .AN(oc8051_sfr1_n132), .B(
        oc8051_sfr1_n133), .C(oc8051_sfr1_n134), .D(oc8051_sfr1_n135), .Y(
        oc8051_sfr1_n131) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u130 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n131), .B0(des_acc[5]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n130) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u129 ( .B0(sfr_out[5]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n130), .Y(oc8051_sfr1_n239) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u128 ( .A0(oc8051_sfr1_ip_4_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[4]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[4]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n125) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u127 ( .A0(oc8051_sfr1_tl0[4]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_4_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[4]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n126) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u126 ( .A0(oc8051_sfr1_p3_data_4_), .A1(
        oc8051_sfr1_n65), .B0(sp[4]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[4]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n127) );
  AO22_X0P5M_A12TS oc8051_sfr1_u125 ( .A0(oc8051_sfr1_sbuf[4]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[4]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n129) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u124 ( .A0(dptr_lo[4]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_4_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n129), 
        .Y(oc8051_sfr1_n128) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u123 ( .A(oc8051_sfr1_n125), .B(
        oc8051_sfr1_n126), .C(oc8051_sfr1_n127), .D(oc8051_sfr1_n128), .Y(
        oc8051_sfr1_n118) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u122 ( .A0(oc8051_sfr1_p1_data_4_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_4_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_4_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n119) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u121 ( .A0(oc8051_sfr1_rcap2h[4]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[4]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n122) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u120 ( .A0(oc8051_sfr1_tl1[4]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tr0), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n123) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u119 ( .A0(oc8051_sfr1_th2[4]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_tclk), .B1(oc8051_sfr1_n47), .C0(
        oc8051_sfr1_rcap2l[4]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n124) );
  AND3_X0P5M_A12TS oc8051_sfr1_u118 ( .A(oc8051_sfr1_n122), .B(
        oc8051_sfr1_n123), .C(oc8051_sfr1_n124), .Y(oc8051_sfr1_n120) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u117 ( .A0(acc[4]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_4_), .B1(oc8051_sfr1_n41), .C0(
        oc8051_sfr1_psw_4_), .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n121) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u116 ( .AN(oc8051_sfr1_n118), .B(
        oc8051_sfr1_n119), .C(oc8051_sfr1_n120), .D(oc8051_sfr1_n121), .Y(
        oc8051_sfr1_n117) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u115 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n117), .B0(des_acc[4]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n116) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u114 ( .B0(sfr_out[4]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n116), .Y(oc8051_sfr1_n240) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u113 ( .A0(oc8051_sfr1_ip_3_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[3]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[3]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n111) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u112 ( .A0(oc8051_sfr1_tl0[3]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_3_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[3]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n112) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u111 ( .A0(oc8051_sfr1_p3_data_3_), .A1(
        oc8051_sfr1_n65), .B0(sp[3]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[3]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n113) );
  AO22_X0P5M_A12TS oc8051_sfr1_u110 ( .A0(oc8051_sfr1_sbuf[3]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[3]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n115) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u109 ( .A0(dptr_lo[3]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_3_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n115), 
        .Y(oc8051_sfr1_n114) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u108 ( .A(oc8051_sfr1_n111), .B(
        oc8051_sfr1_n112), .C(oc8051_sfr1_n113), .D(oc8051_sfr1_n114), .Y(
        oc8051_sfr1_n104) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u107 ( .A0(oc8051_sfr1_p1_data_3_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_3_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_3_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n105) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u106 ( .A0(oc8051_sfr1_rcap2h[3]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[3]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n108) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u105 ( .A0(oc8051_sfr1_tl1[3]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_3_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n109) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u104 ( .A0(oc8051_sfr1_th2[3]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_3_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[3]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n110)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u103 ( .A(oc8051_sfr1_n108), .B(
        oc8051_sfr1_n109), .C(oc8051_sfr1_n110), .Y(oc8051_sfr1_n106) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u102 ( .A0(acc[3]), .A1(oc8051_sfr1_n40), 
        .B0(oc8051_sfr1_p2_data_3_), .B1(oc8051_sfr1_n41), .C0(
        oc8051_sfr1_psw_3_), .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n107) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u101 ( .AN(oc8051_sfr1_n104), .B(
        oc8051_sfr1_n105), .C(oc8051_sfr1_n106), .D(oc8051_sfr1_n107), .Y(
        oc8051_sfr1_n103) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u100 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n103), .B0(des_acc[3]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n102) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u99 ( .B0(sfr_out[3]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n102), .Y(oc8051_sfr1_n241) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u98 ( .A0(oc8051_sfr1_ip_2_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[2]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[2]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n97) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u97 ( .A0(oc8051_sfr1_tl0[2]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_2_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[2]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n98) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u96 ( .A0(oc8051_sfr1_p3_data_2_), .A1(
        oc8051_sfr1_n65), .B0(sp[2]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[2]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n99) );
  AO22_X0P5M_A12TS oc8051_sfr1_u95 ( .A0(oc8051_sfr1_sbuf[2]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[2]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n101) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u94 ( .A0(dptr_lo[2]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_2_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n101), 
        .Y(oc8051_sfr1_n100) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u93 ( .A(oc8051_sfr1_n97), .B(oc8051_sfr1_n98), 
        .C(oc8051_sfr1_n99), .D(oc8051_sfr1_n100), .Y(oc8051_sfr1_n90) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u92 ( .A0(oc8051_sfr1_p1_data_2_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_2_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_2_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n91) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u91 ( .A0(oc8051_sfr1_rcap2h[2]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[2]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n94) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u90 ( .A0(oc8051_sfr1_tl1[2]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_2_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n95) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u89 ( .A0(oc8051_sfr1_th2[2]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_2_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[2]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n96)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u88 ( .A(oc8051_sfr1_n94), .B(oc8051_sfr1_n95), 
        .C(oc8051_sfr1_n96), .Y(oc8051_sfr1_n92) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u87 ( .A0(acc[2]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_2_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_2_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n93) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u86 ( .AN(oc8051_sfr1_n90), .B(
        oc8051_sfr1_n91), .C(oc8051_sfr1_n92), .D(oc8051_sfr1_n93), .Y(
        oc8051_sfr1_n89) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u85 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n89), .B0(des_acc[2]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n88) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u84 ( .B0(sfr_out[2]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n88), .Y(oc8051_sfr1_n242) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u83 ( .A0(oc8051_sfr1_ip_1_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[1]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[1]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n83) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u82 ( .A0(oc8051_sfr1_tl0[1]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_1_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[1]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n84) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u81 ( .A0(oc8051_sfr1_p3_data_1_), .A1(
        oc8051_sfr1_n65), .B0(sp[1]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[1]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n85) );
  AO22_X0P5M_A12TS oc8051_sfr1_u80 ( .A0(oc8051_sfr1_sbuf[1]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[1]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n87) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u79 ( .A0(dptr_lo[1]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_1_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n87), 
        .Y(oc8051_sfr1_n86) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u78 ( .A(oc8051_sfr1_n83), .B(oc8051_sfr1_n84), 
        .C(oc8051_sfr1_n85), .D(oc8051_sfr1_n86), .Y(oc8051_sfr1_n76) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u77 ( .A0(oc8051_sfr1_p1_data_1_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_1_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_1_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n77) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u76 ( .A0(oc8051_sfr1_rcap2h[1]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[1]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n80) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u75 ( .A0(oc8051_sfr1_tl1[1]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_1_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n81) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u74 ( .A0(oc8051_sfr1_th2[1]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_1_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[1]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n82)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u73 ( .A(oc8051_sfr1_n80), .B(oc8051_sfr1_n81), 
        .C(oc8051_sfr1_n82), .Y(oc8051_sfr1_n78) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u72 ( .A0(acc[1]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_1_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_1_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n79) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u71 ( .AN(oc8051_sfr1_n76), .B(
        oc8051_sfr1_n77), .C(oc8051_sfr1_n78), .D(oc8051_sfr1_n79), .Y(
        oc8051_sfr1_n75) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u70 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n75), .B0(des_acc[1]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n74) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u69 ( .B0(sfr_out[1]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n74), .Y(oc8051_sfr1_n243) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u68 ( .A0(oc8051_sfr1_ip_0_), .A1(
        oc8051_sfr1_n71), .B0(oc8051_sfr1_th0[0]), .B1(oc8051_sfr1_n72), .C0(
        oc8051_sfr1_tmod[0]), .C1(oc8051_sfr1_n73), .Y(oc8051_sfr1_n56) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u67 ( .A0(oc8051_sfr1_tl0[0]), .A1(
        oc8051_sfr1_n68), .B0(oc8051_sfr1_p0_data_0_), .B1(oc8051_sfr1_n69), 
        .C0(oc8051_sfr1_th1[0]), .C1(oc8051_sfr1_n70), .Y(oc8051_sfr1_n57) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u66 ( .A0(oc8051_sfr1_p3_data_0_), .A1(
        oc8051_sfr1_n65), .B0(sp[0]), .B1(oc8051_sfr1_n66), .C0(dptr_hi[0]), 
        .C1(oc8051_sfr1_n67), .Y(oc8051_sfr1_n58) );
  AO22_X0P5M_A12TS oc8051_sfr1_u65 ( .A0(oc8051_sfr1_sbuf[0]), .A1(
        oc8051_sfr1_n63), .B0(oc8051_sfr1_pcon[0]), .B1(oc8051_sfr1_n64), .Y(
        oc8051_sfr1_n62) );
  AOI221_X0P5M_A12TS oc8051_sfr1_u64 ( .A0(dptr_lo[0]), .A1(oc8051_sfr1_n60), 
        .B0(oc8051_sfr1_scon_0_), .B1(oc8051_sfr1_n61), .C0(oc8051_sfr1_n62), 
        .Y(oc8051_sfr1_n59) );
  NAND4_X0P5A_A12TS oc8051_sfr1_u63 ( .A(oc8051_sfr1_n56), .B(oc8051_sfr1_n57), 
        .C(oc8051_sfr1_n58), .D(oc8051_sfr1_n59), .Y(oc8051_sfr1_n36) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u62 ( .A0(oc8051_sfr1_p1_data_0_), .A1(
        oc8051_sfr1_n53), .B0(oc8051_sfr1_ie_0_), .B1(oc8051_sfr1_n54), .C0(
        oc8051_sfr1_b_reg_0_), .C1(oc8051_sfr1_n55), .Y(oc8051_sfr1_n37) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u61 ( .A0(oc8051_sfr1_rcap2h[0]), .A1(
        oc8051_sfr1_n51), .B0(oc8051_sfr1_tl2[0]), .B1(oc8051_sfr1_n52), .Y(
        oc8051_sfr1_n43) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u60 ( .A0(oc8051_sfr1_tl1[0]), .A1(
        oc8051_sfr1_n49), .B0(oc8051_sfr1_tcon_0_), .B1(oc8051_sfr1_n50), .Y(
        oc8051_sfr1_n44) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u59 ( .A0(oc8051_sfr1_th2[0]), .A1(
        oc8051_sfr1_n46), .B0(oc8051_sfr1_t2con_0_), .B1(oc8051_sfr1_n47), 
        .C0(oc8051_sfr1_rcap2l[0]), .C1(oc8051_sfr1_n48), .Y(oc8051_sfr1_n45)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_u58 ( .A(oc8051_sfr1_n43), .B(oc8051_sfr1_n44), 
        .C(oc8051_sfr1_n45), .Y(oc8051_sfr1_n38) );
  AOI222_X0P5M_A12TS oc8051_sfr1_u57 ( .A0(acc[0]), .A1(oc8051_sfr1_n40), .B0(
        oc8051_sfr1_p2_data_0_), .B1(oc8051_sfr1_n41), .C0(oc8051_sfr1_psw_0_), 
        .C1(oc8051_sfr1_n42), .Y(oc8051_sfr1_n39) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_u56 ( .AN(oc8051_sfr1_n36), .B(
        oc8051_sfr1_n37), .C(oc8051_sfr1_n38), .D(oc8051_sfr1_n39), .Y(
        oc8051_sfr1_n34) );
  AOI22_X0P5M_A12TS oc8051_sfr1_u55 ( .A0(oc8051_sfr1_n33), .A1(
        oc8051_sfr1_n34), .B0(des_acc[0]), .B1(oc8051_sfr1_n35), .Y(
        oc8051_sfr1_n32) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_u54 ( .B0(sfr_out[0]), .B1(oc8051_sfr1_n1020), 
        .A0N(oc8051_sfr1_n32), .Y(oc8051_sfr1_n244) );
  NOR3_X0P5A_A12TS oc8051_sfr1_u53 ( .A(oc8051_sfr1_n30), .B(
        oc8051_sfr1_prescaler_2_), .C(oc8051_sfr1_n31), .Y(oc8051_sfr1_n259)
         );
  INV_X0P5B_A12TS oc8051_sfr1_u52 ( .A(oc8051_sfr1_prescaler_0_), .Y(
        oc8051_sfr1_n258) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u51 ( .A(oc8051_sfr1_ip_0_), .B(
        oc8051_sfr1_ip_2_), .C(oc8051_sfr1_ip_1_), .D(oc8051_sfr1_ip_3_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n22) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u50 ( .A(oc8051_sfr1_scon_0_), .B(
        oc8051_sfr1_scon_2_), .C(oc8051_sfr1_scon_1_), .D(oc8051_sfr1_scon_3_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n18) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u49 ( .A(oc8051_sfr1_ie_4_), .B(
        oc8051_sfr1_ie_6_), .C(oc8051_sfr1_ie_5_), .D(oc8051_sfr1_ie_7_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n21) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u48 ( .A(oc8051_sfr1_ip_4_), .B(
        oc8051_sfr1_ip_6_), .C(oc8051_sfr1_ip_5_), .D(oc8051_sfr1_ip_7_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n23) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u47 ( .A(oc8051_sfr1_scon_4_), .B(
        oc8051_sfr1_scon_6_), .C(oc8051_sfr1_scon_5_), .D(oc8051_sfr1_scon_7_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n19) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u46 ( .A(oc8051_sfr1_ie_0_), .B(
        oc8051_sfr1_ie_2_), .C(oc8051_sfr1_ie_1_), .D(oc8051_sfr1_ie_3_), .S0(
        rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n20) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u45 ( .A(oc8051_sfr1_n22), .B(oc8051_sfr1_n23), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1340) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u44 ( .A(oc8051_sfr1_n20), .B(oc8051_sfr1_n21), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1350) );
  MXIT2_X0P7M_A12TS oc8051_sfr1_u43 ( .A(oc8051_sfr1_n212), .B(descy), .S0(
        oc8051_sfr1_n213), .Y(oc8051_sfr1_n7) );
  MXIT2_X0P7M_A12TS oc8051_sfr1_u42 ( .A(oc8051_sfr1_n6), .B(oc8051_sfr1_n7), 
        .S0(oc8051_sfr1_n208), .Y(oc8051_sfr1_n1400) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u41 ( .A(oc8051_sfr1_n18), .B(oc8051_sfr1_n19), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1370) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u40 ( .A(oc8051_sfr1_p1_data_0_), .B(
        oc8051_sfr1_p1_data_2_), .C(oc8051_sfr1_p1_data_1_), .D(
        oc8051_sfr1_p1_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n26) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u39 ( .A(oc8051_sfr1_p2_data_4_), .B(
        oc8051_sfr1_p2_data_6_), .C(oc8051_sfr1_p2_data_5_), .D(
        oc8051_sfr1_p2_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n25) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u38 ( .A(oc8051_sfr1_p1_data_4_), .B(
        oc8051_sfr1_p1_data_6_), .C(oc8051_sfr1_p1_data_5_), .D(
        oc8051_sfr1_p1_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n27) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u37 ( .A(oc8051_sfr1_p2_data_0_), .B(
        oc8051_sfr1_p2_data_2_), .C(oc8051_sfr1_p2_data_1_), .D(
        oc8051_sfr1_p2_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n24) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u36 ( .A(oc8051_sfr1_n26), .B(oc8051_sfr1_n27), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1300) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_u35 ( .A(oc8051_sfr1_n24), .B(oc8051_sfr1_n25), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1310) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u34 ( .A(wr_dat[0]), .B(wr_dat[2]), .C(
        wr_dat[1]), .D(wr_dat[3]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n28) );
  MXIT4_X0P5M_A12TS oc8051_sfr1_u33 ( .A(wr_dat[4]), .B(wr_dat[6]), .C(
        wr_dat[5]), .D(wr_dat[7]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n29) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u32 ( .A(oc8051_sfr1_b_reg_4_), .B(
        oc8051_sfr1_b_reg_6_), .C(oc8051_sfr1_b_reg_5_), .D(
        oc8051_sfr1_b_reg_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n15) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u31 ( .A(oc8051_sfr1_b_reg_0_), .B(
        oc8051_sfr1_b_reg_2_), .C(oc8051_sfr1_b_reg_1_), .D(
        oc8051_sfr1_b_reg_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n14) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u30 ( .A(oc8051_sfr1_n14), .B(oc8051_sfr1_n15), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1330) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u29 ( .A(acc[4]), .B(acc[6]), .C(acc[5]), .D(
        acc[7]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n13) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u28 ( .A(acc[0]), .B(acc[2]), .C(acc[1]), .D(
        acc[3]), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n12) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u27 ( .A(oc8051_sfr1_n12), .B(oc8051_sfr1_n13), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1270) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u26 ( .A(oc8051_sfr1_tr0), .B(oc8051_sfr1_tr1), 
        .C(oc8051_sfr1_tcon_5_), .D(oc8051_sfr1_tcon_7_), .S0(rd_addr[1]), 
        .S1(rd_addr[0]), .Y(oc8051_sfr1_n9) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u25 ( .A(oc8051_sfr1_tcon_0_), .B(
        oc8051_sfr1_tcon_2_), .C(oc8051_sfr1_tcon_1_), .D(oc8051_sfr1_tcon_3_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n8) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u24 ( .A(oc8051_sfr1_n8), .B(oc8051_sfr1_n9), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1360) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u23 ( .A(oc8051_sfr1_psw_4_), .B(srcac), .C(
        oc8051_sfr1_psw_5_), .D(cy), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n11) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u22 ( .A(oc8051_sfr1_psw_0_), .B(
        oc8051_sfr1_psw_2_), .C(oc8051_sfr1_psw_1_), .D(oc8051_sfr1_psw_3_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n10) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u21 ( .A(oc8051_sfr1_n10), .B(oc8051_sfr1_n11), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1280) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u20 ( .A(oc8051_sfr1_t2con_0_), .B(
        oc8051_sfr1_t2con_2_), .C(oc8051_sfr1_t2con_1_), .D(
        oc8051_sfr1_t2con_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n16) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u19 ( .A(oc8051_sfr1_n16), .B(oc8051_sfr1_n17), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1380) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u18 ( .A(oc8051_sfr1_tclk), .B(
        oc8051_sfr1_t2con_6_), .C(oc8051_sfr1_rclk), .D(oc8051_sfr1_t2con_7_), 
        .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(oc8051_sfr1_n17) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u17 ( .A(oc8051_sfr1_n28), .B(oc8051_sfr1_n29), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n6) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u16 ( .A(oc8051_sfr1_p0_data_4_), .B(
        oc8051_sfr1_p0_data_6_), .C(oc8051_sfr1_p0_data_5_), .D(
        oc8051_sfr1_p0_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n3) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u15 ( .A(oc8051_sfr1_p0_data_0_), .B(
        oc8051_sfr1_p0_data_2_), .C(oc8051_sfr1_p0_data_1_), .D(
        oc8051_sfr1_p0_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n2) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u14 ( .A(oc8051_sfr1_n2), .B(oc8051_sfr1_n3), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1290) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u13 ( .A(oc8051_sfr1_p3_data_0_), .B(
        oc8051_sfr1_p3_data_2_), .C(oc8051_sfr1_p3_data_1_), .D(
        oc8051_sfr1_p3_data_3_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n4) );
  MXT2_X0P5M_A12TS oc8051_sfr1_u12 ( .A(oc8051_sfr1_n4), .B(oc8051_sfr1_n5), 
        .S0(rd_addr[2]), .Y(oc8051_sfr1_n1320) );
  MXT4_X0P5M_A12TS oc8051_sfr1_u11 ( .A(oc8051_sfr1_p3_data_4_), .B(
        oc8051_sfr1_p3_data_6_), .C(oc8051_sfr1_p3_data_5_), .D(
        oc8051_sfr1_p3_data_7_), .S0(rd_addr[1]), .S1(rd_addr[0]), .Y(
        oc8051_sfr1_n5) );
  NOR2_X0P5M_A12TS oc8051_sfr1_u10 ( .A(rd_addr[2]), .B(rd_addr[1]), .Y(
        oc8051_sfr1_n233) );
  AND4_X0P7M_A12TS oc8051_sfr1_u9 ( .A(rd_addr[1]), .B(oc8051_sfr1_n219), .C(
        rd_addr[7]), .D(oc8051_sfr1_n257), .Y(oc8051_sfr1_n231) );
  AND3_X0P7M_A12TS oc8051_sfr1_u8 ( .A(rd_addr[0]), .B(oc8051_sfr1_n182), .C(
        oc8051_sfr1_n169), .Y(oc8051_sfr1_n73) );
  AND4_X0P7M_A12TS oc8051_sfr1_u7 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(
        oc8051_sfr1_n172), .D(oc8051_sfr1_n183), .Y(oc8051_sfr1_n67) );
  NOR2_X0P5M_A12TS oc8051_sfr1_u6 ( .A(oc8051_sfr1_n185), .B(rd_addr[0]), .Y(
        oc8051_sfr1_n167) );
  INV_X0P5M_A12TS oc8051_sfr1_u5 ( .A(rd_addr[1]), .Y(oc8051_sfr1_n185) );
  INV_X0P5M_A12TS oc8051_sfr1_u4 ( .A(rd_addr[0]), .Y(oc8051_sfr1_n174) );
  TIELO_X1M_A12TS oc8051_sfr1_u3 ( .Y(oc8051_sfr1_int_src_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_wr_bit_r_reg ( .D(bit_addr_o), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_wr_bit_r) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_wait_data_reg ( .D(oc8051_sfr1_n1020), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(wait_data) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_pres_ow_reg ( .D(oc8051_sfr1_n259), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_pres_ow) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_2_ ( .D(oc8051_sfr1_n1510), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_0_ ( .D(oc8051_sfr1_n258), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_1_ ( .D(oc8051_sfr1_n1500), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_7_ ( .D(oc8051_sfr1_n237), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_6_ ( .D(oc8051_sfr1_n238), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_5_ ( .D(oc8051_sfr1_n239), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_4_ ( .D(oc8051_sfr1_n240), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_3_ ( .D(oc8051_sfr1_n241), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_2_ ( .D(oc8051_sfr1_n242), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_1_ ( .D(oc8051_sfr1_n243), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_dat0_reg_0_ ( .D(oc8051_sfr1_n244), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_out[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_prescaler_reg_3_ ( .D(oc8051_sfr1_n1520), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_prescaler_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_bit_out_reg ( .D(oc8051_sfr1_n1400), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(sfr_bit) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u77 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_acc1_n61) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u76 ( .A(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_acc1_n60) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u75 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_acc1_n11) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u74 ( .A(
        oc8051_sfr1_oc8051_acc1_n61), .B(oc8051_sfr1_oc8051_acc1_n60), .C(
        oc8051_sfr1_oc8051_acc1_n11), .Y(oc8051_sfr1_oc8051_acc1_n62) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u73 ( .A(n_5_net_), .Y(
        oc8051_sfr1_oc8051_acc1_n66) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u72 ( .A(
        oc8051_sfr1_oc8051_acc1_n66), .B(wr_addr[4]), .C(wr_addr[3]), .Y(
        oc8051_sfr1_oc8051_acc1_n65) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u71 ( .A(wr_addr[6]), .B(
        wr_addr[5]), .C(wr_addr[7]), .D(oc8051_sfr1_oc8051_acc1_n65), .Y(
        oc8051_sfr1_oc8051_acc1_n63) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u70 ( .AN(wr_sfr[1]), .B(
        wr_sfr[0]), .Y(oc8051_sfr1_oc8051_acc1_n64) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u69 ( .A0(
        oc8051_sfr1_oc8051_acc1_n62), .A1(oc8051_sfr1_wr_bit_r), .A2(
        oc8051_sfr1_oc8051_acc1_n63), .B0(oc8051_sfr1_oc8051_acc1_n64), .Y(
        oc8051_sfr1_oc8051_acc1_n57) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u68 ( .AN(wr_sfr[1]), .B(wr_sfr[0]), .Y(oc8051_sfr1_oc8051_acc1_n9) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u67 ( .AN(
        oc8051_sfr1_oc8051_acc1_n63), .B(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_acc1_n59) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u66 ( .A(
        oc8051_sfr1_oc8051_acc1_n57), .B(oc8051_sfr1_oc8051_acc1_n9), .C(
        oc8051_sfr1_oc8051_acc1_n59), .Y(oc8051_sfr1_oc8051_acc1_n33) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u65 ( .A(descy), .B(
        oc8051_sfr1_oc8051_acc1_n33), .Y(oc8051_sfr1_oc8051_acc1_n19) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u64 ( .A(oc8051_sfr1_oc8051_acc1_n19), .Y(oc8051_sfr1_oc8051_acc1_n32) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u63 ( .A(oc8051_sfr1_oc8051_acc1_n62), .Y(oc8051_sfr1_oc8051_acc1_n53) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u62 ( .A0(
        oc8051_sfr1_oc8051_acc1_n32), .A1(oc8051_sfr1_oc8051_acc1_n53), .B0(
        des2[0]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n54) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u61 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_acc1_n60), .C(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_acc1_n49) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u60 ( .A(
        oc8051_sfr1_oc8051_acc1_n11), .B(oc8051_sfr1_oc8051_acc1_n60), .C(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_acc1_n45) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u59 ( .A(
        oc8051_sfr1_oc8051_acc1_n61), .B(oc8051_sfr1_oc8051_acc1_n60), .C(
        wr_addr[0]), .Y(oc8051_sfr1_oc8051_acc1_n47) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u58 ( .A(
        oc8051_sfr1_oc8051_acc1_n49), .B(oc8051_sfr1_oc8051_acc1_n45), .C(
        oc8051_sfr1_oc8051_acc1_n47), .Y(oc8051_sfr1_oc8051_acc1_n34) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u57 ( .A(
        oc8051_sfr1_oc8051_acc1_n11), .B(oc8051_sfr1_oc8051_acc1_n61), .C(
        wr_addr[2]), .Y(oc8051_sfr1_oc8051_acc1_n46) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u56 ( .A(oc8051_sfr1_oc8051_acc1_n46), .Y(oc8051_sfr1_oc8051_acc1_n31) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u55 ( .A(
        oc8051_sfr1_oc8051_acc1_n34), .B(oc8051_sfr1_oc8051_acc1_n31), .Y(
        oc8051_sfr1_oc8051_acc1_n24) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u54 ( .A(oc8051_sfr1_oc8051_acc1_n33), .Y(oc8051_sfr1_oc8051_acc1_n25) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u53 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_acc1_n33), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_acc1_n23) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u52 ( .A(
        oc8051_sfr1_oc8051_acc1_n60), .B(wr_addr[1]), .C(
        oc8051_sfr1_oc8051_acc1_n11), .Y(oc8051_sfr1_oc8051_acc1_n27) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u51 ( .A(oc8051_sfr1_oc8051_acc1_n59), .Y(oc8051_sfr1_oc8051_acc1_n58) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u50 ( .A(
        oc8051_sfr1_oc8051_acc1_n58), .B(oc8051_sfr1_oc8051_acc1_n9), .C(
        oc8051_sfr1_oc8051_acc1_n57), .Y(oc8051_sfr1_oc8051_acc1_n22) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u49 ( .A0(
        oc8051_sfr1_oc8051_acc1_n33), .A1(oc8051_sfr1_oc8051_acc1_n27), .B0(
        oc8051_sfr1_oc8051_acc1_n22), .Y(oc8051_sfr1_oc8051_acc1_n17) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u48 ( .A0(
        oc8051_sfr1_oc8051_acc1_n24), .A1(oc8051_sfr1_oc8051_acc1_n25), .B0(
        oc8051_sfr1_oc8051_acc1_n23), .C0(oc8051_sfr1_oc8051_acc1_n17), .Y(
        oc8051_sfr1_oc8051_acc1_n56) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u47 ( .AN(
        oc8051_sfr1_oc8051_acc1_n57), .B(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n8) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u46 ( .A0(acc[0]), .A1(
        oc8051_sfr1_oc8051_acc1_n56), .B0(des_acc[0]), .B1(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n55) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u45 ( .A(
        oc8051_sfr1_oc8051_acc1_n54), .B(oc8051_sfr1_oc8051_acc1_n55), .Y(
        oc8051_sfr1_oc8051_acc1_acc_0_) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u44 ( .A(
        oc8051_sfr1_oc8051_acc1_n49), .B(oc8051_sfr1_oc8051_acc1_n45), .C(
        oc8051_sfr1_oc8051_acc1_n46), .Y(oc8051_sfr1_oc8051_acc1_n52) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u43 ( .A(
        oc8051_sfr1_oc8051_acc1_n33), .B(oc8051_sfr1_oc8051_acc1_n53), .Y(
        oc8051_sfr1_oc8051_acc1_n26) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u42 ( .A(
        oc8051_sfr1_oc8051_acc1_n26), .B(oc8051_sfr1_oc8051_acc1_n23), .C(
        oc8051_sfr1_oc8051_acc1_n17), .Y(oc8051_sfr1_oc8051_acc1_n35) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u41 ( .A0(
        oc8051_sfr1_oc8051_acc1_n33), .A1(oc8051_sfr1_oc8051_acc1_n52), .B0(
        oc8051_sfr1_oc8051_acc1_n35), .C0(acc[1]), .Y(
        oc8051_sfr1_oc8051_acc1_n50) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u40 ( .A0(des_acc[1]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[1]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n51) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u39 ( .A0(
        oc8051_sfr1_oc8051_acc1_n19), .A1(oc8051_sfr1_oc8051_acc1_n47), .B0(
        oc8051_sfr1_oc8051_acc1_n50), .C0(oc8051_sfr1_oc8051_acc1_n51), .Y(
        oc8051_sfr1_oc8051_acc1_acc_1_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u38 ( .A(des_acc[2]), .B(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n42) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u37 ( .A(oc8051_sfr1_oc8051_acc1_n49), .Y(oc8051_sfr1_oc8051_acc1_n39) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u36 ( .A(oc8051_sfr1_oc8051_acc1_n35), .Y(oc8051_sfr1_oc8051_acc1_n48) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u35 ( .A0(
        oc8051_sfr1_oc8051_acc1_n46), .A1(oc8051_sfr1_oc8051_acc1_n47), .B0(
        oc8051_sfr1_oc8051_acc1_n25), .C0(oc8051_sfr1_oc8051_acc1_n48), .Y(
        oc8051_sfr1_oc8051_acc1_n41) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u34 ( .A0(
        oc8051_sfr1_oc8051_acc1_n39), .A1(oc8051_sfr1_oc8051_acc1_n33), .B0(
        oc8051_sfr1_oc8051_acc1_n41), .C0(acc[2]), .Y(
        oc8051_sfr1_oc8051_acc1_n43) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u33 ( .A(oc8051_sfr1_oc8051_acc1_n45), .Y(oc8051_sfr1_oc8051_acc1_n40) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u32 ( .A0(
        oc8051_sfr1_oc8051_acc1_n32), .A1(oc8051_sfr1_oc8051_acc1_n40), .B0(
        des2[2]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n44) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u31 ( .A(
        oc8051_sfr1_oc8051_acc1_n42), .B(oc8051_sfr1_oc8051_acc1_n43), .C(
        oc8051_sfr1_oc8051_acc1_n44), .Y(oc8051_sfr1_oc8051_acc1_acc_2_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u30 ( .A(des_acc[3]), .B(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n36) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u29 ( .A0(
        oc8051_sfr1_oc8051_acc1_n40), .A1(oc8051_sfr1_oc8051_acc1_n33), .B0(
        oc8051_sfr1_oc8051_acc1_n41), .C0(acc[3]), .Y(
        oc8051_sfr1_oc8051_acc1_n37) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u28 ( .A0(
        oc8051_sfr1_oc8051_acc1_n39), .A1(oc8051_sfr1_oc8051_acc1_n32), .B0(
        des2[3]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n38) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u27 ( .A(
        oc8051_sfr1_oc8051_acc1_n36), .B(oc8051_sfr1_oc8051_acc1_n37), .C(
        oc8051_sfr1_oc8051_acc1_n38), .Y(oc8051_sfr1_oc8051_acc1_acc_3_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u26 ( .A(des_acc[4]), .B(
        oc8051_sfr1_oc8051_acc1_n8), .Y(oc8051_sfr1_oc8051_acc1_n28) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u25 ( .A0(
        oc8051_sfr1_oc8051_acc1_n33), .A1(oc8051_sfr1_oc8051_acc1_n34), .B0(
        oc8051_sfr1_oc8051_acc1_n35), .C0(acc[4]), .Y(
        oc8051_sfr1_oc8051_acc1_n29) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u24 ( .A0(
        oc8051_sfr1_oc8051_acc1_n31), .A1(oc8051_sfr1_oc8051_acc1_n32), .B0(
        des2[4]), .B1(oc8051_sfr1_oc8051_acc1_n9), .Y(
        oc8051_sfr1_oc8051_acc1_n30) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u23 ( .A(
        oc8051_sfr1_oc8051_acc1_n28), .B(oc8051_sfr1_oc8051_acc1_n29), .C(
        oc8051_sfr1_oc8051_acc1_n30), .Y(oc8051_sfr1_oc8051_acc1_acc_4_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u22 ( .A(oc8051_sfr1_oc8051_acc1_n27), .Y(oc8051_sfr1_oc8051_acc1_n18) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u21 ( .A0(
        oc8051_sfr1_oc8051_acc1_n24), .A1(oc8051_sfr1_oc8051_acc1_n25), .B0(
        oc8051_sfr1_oc8051_acc1_n26), .Y(oc8051_sfr1_oc8051_acc1_n16) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_acc1_u20 ( .A(oc8051_sfr1_oc8051_acc1_n23), .Y(oc8051_sfr1_oc8051_acc1_n10) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u19 ( .A0(
        oc8051_sfr1_oc8051_acc1_n16), .A1(oc8051_sfr1_oc8051_acc1_n10), .A2(
        oc8051_sfr1_oc8051_acc1_n22), .B0(acc[5]), .Y(
        oc8051_sfr1_oc8051_acc1_n20) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u18 ( .A0(des_acc[5]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[5]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n21) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u17 ( .A0(
        oc8051_sfr1_oc8051_acc1_n18), .A1(oc8051_sfr1_oc8051_acc1_n19), .B0(
        oc8051_sfr1_oc8051_acc1_n20), .C0(oc8051_sfr1_oc8051_acc1_n21), .Y(
        oc8051_sfr1_oc8051_acc1_acc_5_) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u16 ( .AN(
        oc8051_sfr1_oc8051_acc1_n16), .B(oc8051_sfr1_oc8051_acc1_n17), .Y(
        oc8051_sfr1_oc8051_acc1_n12) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u15 ( .A0(
        oc8051_sfr1_oc8051_acc1_n10), .A1(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_acc1_n12), .C0(acc[6]), .Y(
        oc8051_sfr1_oc8051_acc1_n13) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u14 ( .A(descy), .B(
        oc8051_sfr1_oc8051_acc1_n11), .C(oc8051_sfr1_oc8051_acc1_n10), .Y(
        oc8051_sfr1_oc8051_acc1_n14) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u13 ( .A0(des_acc[6]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[6]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n15) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u12 ( .A(
        oc8051_sfr1_oc8051_acc1_n13), .B(oc8051_sfr1_oc8051_acc1_n14), .C(
        oc8051_sfr1_oc8051_acc1_n15), .Y(oc8051_sfr1_oc8051_acc1_acc_6_) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u11 ( .A0(
        oc8051_sfr1_oc8051_acc1_n10), .A1(oc8051_sfr1_oc8051_acc1_n11), .B0(
        oc8051_sfr1_oc8051_acc1_n12), .C0(acc[7]), .Y(
        oc8051_sfr1_oc8051_acc1_n5) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u10 ( .A0(des_acc[7]), .A1(
        oc8051_sfr1_oc8051_acc1_n8), .B0(des2[7]), .B1(
        oc8051_sfr1_oc8051_acc1_n9), .Y(oc8051_sfr1_oc8051_acc1_n7) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_acc1_u9 ( .A(oc8051_sfr1_oc8051_acc1_n5), .B(oc8051_sfr1_oc8051_acc1_n6), .C(oc8051_sfr1_oc8051_acc1_n7), .Y(
        oc8051_sfr1_oc8051_acc1_acc_7_) );
  XNOR2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u8 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_1_), .B(oc8051_sfr1_oc8051_acc1_acc_0_), 
        .Y(oc8051_sfr1_oc8051_acc1_n4) );
  XNOR3_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u7 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_2_), .B(oc8051_sfr1_oc8051_acc1_acc_3_), 
        .C(oc8051_sfr1_oc8051_acc1_n4), .Y(oc8051_sfr1_oc8051_acc1_n1) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u6 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_5_), .B(oc8051_sfr1_oc8051_acc1_acc_4_), 
        .Y(oc8051_sfr1_oc8051_acc1_n3) );
  XOR3_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u5 ( .A(
        oc8051_sfr1_oc8051_acc1_acc_7_), .B(oc8051_sfr1_oc8051_acc1_n3), .C(
        oc8051_sfr1_oc8051_acc1_acc_6_), .Y(oc8051_sfr1_oc8051_acc1_n2) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u4 ( .A(oc8051_sfr1_oc8051_acc1_n1), 
        .B(oc8051_sfr1_oc8051_acc1_n2), .Y(oc8051_sfr1_psw_0_) );
  NAND3_X0P5M_A12TS oc8051_sfr1_oc8051_acc1_u3 ( .A(descy), .B(wr_addr[0]), 
        .C(oc8051_sfr1_oc8051_acc1_n10), .Y(oc8051_sfr1_oc8051_acc1_n6) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_0_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_2_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_6_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_1_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_4_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_3_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_7_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_acc1_data_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_acc1_acc_5_), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        acc[5]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_b_register_u37 ( .A(oc8051_sfr1_wr_bit_r), 
        .Y(oc8051_sfr1_oc8051_b_register_n5) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u36 ( .AN(wr_addr[4]), .B(
        wr_addr[3]), .Y(oc8051_sfr1_oc8051_b_register_n28) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u35 ( .A(wr_addr[7]), .B(
        wr_addr[6]), .C(oc8051_sfr1_oc8051_b_register_n28), .D(wr_addr[5]), 
        .Y(oc8051_sfr1_oc8051_b_register_n25) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u34 ( .A(
        oc8051_sfr1_oc8051_b_register_n25), .B(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_b_register_n27) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_b_register_u33 ( .A(descy), .B(
        oc8051_sfr1_oc8051_b_register_n27), .Y(
        oc8051_sfr1_oc8051_b_register_n6) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u32 ( .B0(des_acc[0]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n23) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_b_register_u31 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_b_register_n9) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_b_register_u30 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_b_register_n12) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u29 ( .A(n_5_net_), .B(
        oc8051_sfr1_oc8051_b_register_n27), .Y(
        oc8051_sfr1_oc8051_b_register_n15) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u28 ( .AN(
        oc8051_sfr1_oc8051_b_register_n15), .B(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_b_register_n18) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_b_register_u27 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_wr_bit_r), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_b_register_n26) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u26 ( .A(
        oc8051_sfr1_oc8051_b_register_n25), .B(
        oc8051_sfr1_oc8051_b_register_n9), .C(n_5_net_), .D(
        oc8051_sfr1_oc8051_b_register_n26), .Y(
        oc8051_sfr1_oc8051_b_register_n4) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u25 ( .A0(
        oc8051_sfr1_oc8051_b_register_n9), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(
        oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n24) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u24 ( .A(
        oc8051_sfr1_oc8051_b_register_n23), .B(oc8051_sfr1_b_reg_0_), .S0(
        oc8051_sfr1_oc8051_b_register_n24), .Y(
        oc8051_sfr1_oc8051_b_register_n32) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u23 ( .B0(des_acc[1]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n21) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u22 ( .A0(wr_addr[0]), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(
        oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n22) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u21 ( .A(
        oc8051_sfr1_oc8051_b_register_n21), .B(oc8051_sfr1_b_reg_1_), .S0(
        oc8051_sfr1_oc8051_b_register_n22), .Y(
        oc8051_sfr1_oc8051_b_register_n33) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u20 ( .B0(des_acc[2]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n19) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u19 ( .A0(wr_addr[1]), .A1(
        oc8051_sfr1_oc8051_b_register_n9), .A2(
        oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n20) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u18 ( .A(
        oc8051_sfr1_oc8051_b_register_n19), .B(oc8051_sfr1_b_reg_2_), .S0(
        oc8051_sfr1_oc8051_b_register_n20), .Y(
        oc8051_sfr1_oc8051_b_register_n34) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u17 ( .B0(des_acc[3]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n16) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u16 ( .A0(wr_addr[1]), .A1(
        wr_addr[0]), .A2(oc8051_sfr1_oc8051_b_register_n18), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n17) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u15 ( .A(
        oc8051_sfr1_oc8051_b_register_n16), .B(oc8051_sfr1_b_reg_3_), .S0(
        oc8051_sfr1_oc8051_b_register_n17), .Y(
        oc8051_sfr1_oc8051_b_register_n35) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u14 ( .B0(des_acc[4]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n13) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u13 ( .A(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_b_register_n15), .Y(
        oc8051_sfr1_oc8051_b_register_n3) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u12 ( .A0(
        oc8051_sfr1_oc8051_b_register_n9), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(
        oc8051_sfr1_oc8051_b_register_n3), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n14) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u11 ( .A(
        oc8051_sfr1_oc8051_b_register_n13), .B(oc8051_sfr1_b_reg_4_), .S0(
        oc8051_sfr1_oc8051_b_register_n14), .Y(
        oc8051_sfr1_oc8051_b_register_n36) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u10 ( .B0(des_acc[5]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(
        oc8051_sfr1_oc8051_b_register_n10) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u9 ( .A0(
        oc8051_sfr1_oc8051_b_register_n3), .A1(
        oc8051_sfr1_oc8051_b_register_n12), .A2(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(
        oc8051_sfr1_oc8051_b_register_n11) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u8 ( .A(
        oc8051_sfr1_oc8051_b_register_n10), .B(oc8051_sfr1_b_reg_5_), .S0(
        oc8051_sfr1_oc8051_b_register_n11), .Y(
        oc8051_sfr1_oc8051_b_register_n37) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u7 ( .B0(des_acc[6]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(oc8051_sfr1_oc8051_b_register_n7) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u6 ( .A0(
        oc8051_sfr1_oc8051_b_register_n3), .A1(
        oc8051_sfr1_oc8051_b_register_n9), .A2(wr_addr[1]), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(oc8051_sfr1_oc8051_b_register_n8) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u5 ( .A(
        oc8051_sfr1_oc8051_b_register_n7), .B(oc8051_sfr1_b_reg_6_), .S0(
        oc8051_sfr1_oc8051_b_register_n8), .Y(
        oc8051_sfr1_oc8051_b_register_n38) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u4 ( .B0(des_acc[7]), .B1(
        oc8051_sfr1_oc8051_b_register_n5), .A0N(
        oc8051_sfr1_oc8051_b_register_n6), .Y(oc8051_sfr1_oc8051_b_register_n1) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u3 ( .A0(wr_addr[0]), .A1(
        oc8051_sfr1_oc8051_b_register_n3), .A2(wr_addr[1]), .B0(
        oc8051_sfr1_oc8051_b_register_n4), .Y(oc8051_sfr1_oc8051_b_register_n2) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_b_register_u2 ( .A(
        oc8051_sfr1_oc8051_b_register_n1), .B(oc8051_sfr1_b_reg_7_), .S0(
        oc8051_sfr1_oc8051_b_register_n2), .Y(
        oc8051_sfr1_oc8051_b_register_n39) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_b_register_n34), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_b_register_n38), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_b_register_n32), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_b_register_n36), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_b_register_n33), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_b_register_n37), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_b_register_n35), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_b_register_data_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_b_register_n39), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_b_reg_7_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u55 ( .A(ram_rd_sel[2]), .Y(
        oc8051_sfr1_oc8051_sp1_n36) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u54 ( .A(oc8051_sfr1_oc8051_sp1_n36), 
        .B(ram_rd_sel[0]), .C(ram_rd_sel[1]), .Y(oc8051_sfr1_oc8051_sp1_n22)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u53 ( .A(wb_rst_i), .Y(
        oc8051_sfr1_oc8051_sp1_n37) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_sp1_u52 ( .A(wr_addr[7]), .B(wr_addr[0]), .C(oc8051_sfr1_oc8051_sp1_n35), .D(n_5_net_), .Y(oc8051_sfr1_oc8051_sp1_n34)
         );
  OR6_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u51 ( .A(oc8051_sfr1_wr_bit_r), .B(
        wr_addr[6]), .C(wr_addr[5]), .D(wr_addr[4]), .E(wr_addr[3]), .F(
        oc8051_sfr1_oc8051_sp1_n34), .Y(oc8051_sfr1_oc8051_sp1_n33) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u50 ( .A(oc8051_sfr1_oc8051_sp1_n33), 
        .Y(oc8051_sfr1_oc8051_sp1_n2) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u49 ( .AN(ram_wr_sel[2]), .B(
        ram_wr_sel[0]), .C(ram_wr_sel[1]), .Y(oc8051_sfr1_oc8051_sp1_n8) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u48 ( .A(oc8051_sfr1_oc8051_sp1_n8), 
        .Y(oc8051_sfr1_oc8051_sp1_n1) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_sp1_u47 ( .A(oc8051_sfr1_oc8051_sp1_n2), 
        .B(oc8051_sfr1_oc8051_sp1_n1), .Y(oc8051_sfr1_oc8051_sp1_n5) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_sp1_u46 ( .A(oc8051_sfr1_oc8051_sp1_n8), 
        .B(oc8051_sfr1_oc8051_sp1_n2), .Y(oc8051_sfr1_oc8051_sp1_n4) );
  AO21_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u45 ( .A0(oc8051_sfr1_oc8051_sp1_pop), .A1(oc8051_sfr1_oc8051_sp1_n5), .B0(oc8051_sfr1_oc8051_sp1_n4), .Y(
        oc8051_sfr1_oc8051_sp1_n31) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u44 ( .AN(oc8051_sfr1_oc8051_sp1_n5), .B(oc8051_sfr1_oc8051_sp1_pop), .Y(oc8051_sfr1_oc8051_sp1_n32) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u43 ( .A(oc8051_sfr1_oc8051_sp1_n31), .B(oc8051_sfr1_oc8051_sp1_n32), .S0(oc8051_sfr1_oc8051_sp1_sp_0_), .Y(
        oc8051_sfr1_oc8051_sp1_n30) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u42 ( .B0(wr_dat[0]), .B1(
        oc8051_sfr1_oc8051_sp1_n2), .A0N(oc8051_sfr1_oc8051_sp1_n30), .Y(sp[0]) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u41 ( .A1N(
        oc8051_sfr1_oc8051_sp1_pop), .A0(oc8051_sfr1_oc8051_sp1_n8), .B0(
        oc8051_sfr1_oc8051_sp1_sp_0_), .Y(oc8051_sfr1_oc8051_sp1_n26) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u40 ( .A(oc8051_sfr1_oc8051_sp1_n4), 
        .B(oc8051_sfr1_oc8051_sp1_n5), .C(oc8051_sfr1_oc8051_sp1_n5), .D(
        oc8051_sfr1_oc8051_sp1_n4), .S0(oc8051_sfr1_oc8051_sp1_n26), .S1(
        oc8051_sfr1_oc8051_sp1_sp_1_), .Y(oc8051_sfr1_oc8051_sp1_n29) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u39 ( .A(oc8051_sfr1_oc8051_sp1_sp_1_), .Y(oc8051_sfr1_oc8051_sp1_n27) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u38 ( .AN(
        oc8051_sfr1_oc8051_sp1_n26), .B(oc8051_sfr1_oc8051_sp1_sp_1_), .Y(
        oc8051_sfr1_oc8051_sp1_n28) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u37 ( .A0(
        oc8051_sfr1_oc8051_sp1_n26), .A1(oc8051_sfr1_oc8051_sp1_n27), .B0(
        oc8051_sfr1_oc8051_sp1_n1), .B1(oc8051_sfr1_oc8051_sp1_n28), .Y(
        oc8051_sfr1_oc8051_sp1_n23) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u36 ( .A(oc8051_sfr1_oc8051_sp1_n5), 
        .B(oc8051_sfr1_oc8051_sp1_n4), .C(oc8051_sfr1_oc8051_sp1_n4), .D(
        oc8051_sfr1_oc8051_sp1_n5), .S0(oc8051_sfr1_oc8051_sp1_sp_2_), .S1(
        oc8051_sfr1_oc8051_sp1_n23), .Y(oc8051_sfr1_oc8051_sp1_n25) );
  AO21_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u35 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n25), .Y(sp[2])
         );
  OR2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u34 ( .A(oc8051_sfr1_oc8051_sp1_sp_2_), .B(oc8051_sfr1_oc8051_sp1_n23), .Y(oc8051_sfr1_oc8051_sp1_n24) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u33 ( .A0(
        oc8051_sfr1_oc8051_sp1_n23), .A1(oc8051_sfr1_oc8051_sp1_sp_2_), .B0(
        oc8051_sfr1_oc8051_sp1_n8), .B1(oc8051_sfr1_oc8051_sp1_n24), .Y(
        oc8051_sfr1_oc8051_sp1_n18) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u32 ( .A(oc8051_sfr1_oc8051_sp1_n4), 
        .B(oc8051_sfr1_oc8051_sp1_n5), .C(oc8051_sfr1_oc8051_sp1_n5), .D(
        oc8051_sfr1_oc8051_sp1_n4), .S0(oc8051_sfr1_oc8051_sp1_sp_3_), .S1(
        oc8051_sfr1_oc8051_sp1_n18), .Y(oc8051_sfr1_oc8051_sp1_n21) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u31 ( .A(oc8051_sfr1_oc8051_sp1_sp_3_), .Y(oc8051_sfr1_oc8051_sp1_n19) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u30 ( .AN(
        oc8051_sfr1_oc8051_sp1_n18), .B(oc8051_sfr1_oc8051_sp1_sp_3_), .Y(
        oc8051_sfr1_oc8051_sp1_n20) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u29 ( .A0(
        oc8051_sfr1_oc8051_sp1_n18), .A1(oc8051_sfr1_oc8051_sp1_n19), .B0(
        oc8051_sfr1_oc8051_sp1_n1), .B1(oc8051_sfr1_oc8051_sp1_n20), .Y(
        oc8051_sfr1_oc8051_sp1_n15) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u28 ( .A(oc8051_sfr1_oc8051_sp1_n5), 
        .B(oc8051_sfr1_oc8051_sp1_n4), .C(oc8051_sfr1_oc8051_sp1_n4), .D(
        oc8051_sfr1_oc8051_sp1_n5), .S0(oc8051_sfr1_oc8051_sp1_sp_4_), .S1(
        oc8051_sfr1_oc8051_sp1_n15), .Y(oc8051_sfr1_oc8051_sp1_n17) );
  OR2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u27 ( .A(oc8051_sfr1_oc8051_sp1_sp_4_), .B(oc8051_sfr1_oc8051_sp1_n15), .Y(oc8051_sfr1_oc8051_sp1_n16) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u26 ( .A0(
        oc8051_sfr1_oc8051_sp1_n15), .A1(oc8051_sfr1_oc8051_sp1_sp_4_), .B0(
        oc8051_sfr1_oc8051_sp1_n8), .B1(oc8051_sfr1_oc8051_sp1_n16), .Y(
        oc8051_sfr1_oc8051_sp1_n11) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u25 ( .A(oc8051_sfr1_oc8051_sp1_n4), 
        .B(oc8051_sfr1_oc8051_sp1_n5), .C(oc8051_sfr1_oc8051_sp1_n5), .D(
        oc8051_sfr1_oc8051_sp1_n4), .S0(oc8051_sfr1_oc8051_sp1_sp_5_), .S1(
        oc8051_sfr1_oc8051_sp1_n11), .Y(oc8051_sfr1_oc8051_sp1_n14) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_sp1_u24 ( .A(oc8051_sfr1_oc8051_sp1_sp_5_), .Y(oc8051_sfr1_oc8051_sp1_n12) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u23 ( .AN(
        oc8051_sfr1_oc8051_sp1_n11), .B(oc8051_sfr1_oc8051_sp1_sp_5_), .Y(
        oc8051_sfr1_oc8051_sp1_n13) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u22 ( .A0(
        oc8051_sfr1_oc8051_sp1_n11), .A1(oc8051_sfr1_oc8051_sp1_n12), .B0(
        oc8051_sfr1_oc8051_sp1_n1), .B1(oc8051_sfr1_oc8051_sp1_n13), .Y(
        oc8051_sfr1_oc8051_sp1_n9) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u21 ( .A(oc8051_sfr1_oc8051_sp1_n5), 
        .B(oc8051_sfr1_oc8051_sp1_n4), .C(oc8051_sfr1_oc8051_sp1_n4), .D(
        oc8051_sfr1_oc8051_sp1_n5), .S0(oc8051_sfr1_oc8051_sp1_sp_6_), .S1(
        oc8051_sfr1_oc8051_sp1_n9), .Y(oc8051_sfr1_oc8051_sp1_n10) );
  OR2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u20 ( .A(oc8051_sfr1_oc8051_sp1_sp_6_), .B(oc8051_sfr1_oc8051_sp1_n9), .Y(oc8051_sfr1_oc8051_sp1_n7) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u19 ( .A0(oc8051_sfr1_oc8051_sp1_n7), .A1(oc8051_sfr1_oc8051_sp1_n8), .B0(oc8051_sfr1_oc8051_sp1_sp_6_), .B1(
        oc8051_sfr1_oc8051_sp1_n9), .Y(oc8051_sfr1_oc8051_sp1_n6) );
  MXT4_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u18 ( .A(oc8051_sfr1_oc8051_sp1_n4), 
        .B(oc8051_sfr1_oc8051_sp1_n5), .C(oc8051_sfr1_oc8051_sp1_n5), .D(
        oc8051_sfr1_oc8051_sp1_n4), .S0(oc8051_sfr1_oc8051_sp1_sp_7_), .S1(
        oc8051_sfr1_oc8051_sp1_n6), .Y(oc8051_sfr1_oc8051_sp1_n3) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u17 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_0_), .B(oc8051_sfr1_oc8051_sp1_n130), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[0]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u16 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_1_), .B(oc8051_sfr1_oc8051_sp1_n140), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[1]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u15 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_2_), .B(oc8051_sfr1_oc8051_sp1_n150), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[2]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u14 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_3_), .B(oc8051_sfr1_oc8051_sp1_n160), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[3]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u13 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_4_), .B(oc8051_sfr1_oc8051_sp1_n170), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[4]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u12 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_5_), .B(oc8051_sfr1_oc8051_sp1_n180), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[5]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u11 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_6_), .B(oc8051_sfr1_oc8051_sp1_n190), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[6]) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u10 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_7_), .B(oc8051_sfr1_oc8051_sp1_n200), .S0(
        oc8051_sfr1_oc8051_sp1_n1), .Y(sp_w[7]) );
  AO21_X0P7M_A12TS oc8051_sfr1_oc8051_sp1_u9 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n29), .Y(sp[1])
         );
  AO21_X0P7M_A12TS oc8051_sfr1_oc8051_sp1_u8 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n10), .Y(sp[6])
         );
  AO21_X0P7M_A12TS oc8051_sfr1_oc8051_sp1_u7 ( .A0(wr_dat[5]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n14), .Y(sp[5])
         );
  AO21_X0P7M_A12TS oc8051_sfr1_oc8051_sp1_u6 ( .A0(wr_dat[7]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n3), .Y(sp[7])
         );
  AO21_X0P7M_A12TS oc8051_sfr1_oc8051_sp1_u5 ( .A0(wr_dat[4]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n17), .Y(sp[4])
         );
  AO21_X0P7M_A12TS oc8051_sfr1_oc8051_sp1_u4 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_sp1_n2), .B0(oc8051_sfr1_oc8051_sp1_n21), .Y(sp[3])
         );
  NOR2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_u3 ( .A(wr_addr[2]), .B(wr_addr[1]), 
        .Y(oc8051_sfr1_oc8051_sp1_n35) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_5_ ( .D(sp[5]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_3_ ( .D(sp[3]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_4_ ( .D(sp[4]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_6_ ( .D(sp[6]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_6_) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_0_ ( .D(sp[0]), .CK(wb_clk_i), 
        .SN(oc8051_sfr1_oc8051_sp1_n37), .Q(oc8051_sfr1_oc8051_sp1_sp_0_) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_2_ ( .D(sp[2]), .CK(wb_clk_i), 
        .SN(oc8051_sfr1_oc8051_sp1_n37), .Q(oc8051_sfr1_oc8051_sp1_sp_2_) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_1_ ( .D(sp[1]), .CK(wb_clk_i), 
        .SN(oc8051_sfr1_oc8051_sp1_n37), .Q(oc8051_sfr1_oc8051_sp1_sp_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_sp_reg_7_ ( .D(sp[7]), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_sp1_sp_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_sp1_pop_reg ( .D(
        oc8051_sfr1_oc8051_sp1_n22), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_sp1_pop) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u2 ( .A(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[7]), .B(
        oc8051_sfr1_oc8051_sp1_sp_7_), .Y(oc8051_sfr1_oc8051_sp1_n200) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_0_), .Y(oc8051_sfr1_oc8051_sp1_n130) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_1 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_1_), .B(oc8051_sfr1_oc8051_sp1_sp_0_), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[2]), .S(
        oc8051_sfr1_oc8051_sp1_n140) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_5 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_5_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[5]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[6]), .S(
        oc8051_sfr1_oc8051_sp1_n180) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_3 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_3_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[3]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[4]), .S(
        oc8051_sfr1_oc8051_sp1_n160) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_4 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_4_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[4]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[5]), .S(
        oc8051_sfr1_oc8051_sp1_n170) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_2 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_2_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[2]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[3]), .S(
        oc8051_sfr1_oc8051_sp1_n150) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_sp1_add_102_s2_u1_1_6 ( .A(
        oc8051_sfr1_oc8051_sp1_sp_6_), .B(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[6]), .CO(
        oc8051_sfr1_oc8051_sp1_add_102_s2_carry[7]), .S(
        oc8051_sfr1_oc8051_sp1_n190) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u32 ( .A(wr_sfr[1]), .B(wr_sfr[0]), 
        .Y(oc8051_sfr1_oc8051_dptr1_n4) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u31 ( .AN(wr_addr[2]), .B(
        wr_addr[1]), .C(n_5_net_), .D(wr_addr[7]), .Y(
        oc8051_sfr1_oc8051_dptr1_n15) );
  OR6_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u30 ( .A(oc8051_sfr1_wr_bit_r), .B(
        wr_addr[6]), .C(wr_addr[5]), .D(wr_addr[4]), .E(wr_addr[3]), .F(
        oc8051_sfr1_oc8051_dptr1_n15), .Y(oc8051_sfr1_oc8051_dptr1_n2) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_dptr1_u29 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_dptr1_n3) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_dptr1_u28 ( .A(
        oc8051_sfr1_oc8051_dptr1_n2), .B(oc8051_sfr1_oc8051_dptr1_n4), .C(
        oc8051_sfr1_oc8051_dptr1_n3), .Y(oc8051_sfr1_oc8051_dptr1_n7) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_dptr1_u27 ( .A(
        oc8051_sfr1_oc8051_dptr1_n4), .B(oc8051_sfr1_oc8051_dptr1_n7), .Y(
        oc8051_sfr1_oc8051_dptr1_n6) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u26 ( .A0(dptr_hi[0]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[0]), .Y(oc8051_sfr1_oc8051_dptr1_n14) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u25 ( .B0(des2[0]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n14), .Y(
        oc8051_sfr1_oc8051_dptr1_n18) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u24 ( .A0(dptr_hi[1]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[1]), .Y(oc8051_sfr1_oc8051_dptr1_n13) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u23 ( .B0(des2[1]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n13), .Y(
        oc8051_sfr1_oc8051_dptr1_n19) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u22 ( .A0(dptr_hi[2]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[2]), .Y(oc8051_sfr1_oc8051_dptr1_n12) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u21 ( .B0(des2[2]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n12), .Y(
        oc8051_sfr1_oc8051_dptr1_n20) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u20 ( .A0(dptr_hi[3]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[3]), .Y(oc8051_sfr1_oc8051_dptr1_n11) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u19 ( .B0(des2[3]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n11), .Y(
        oc8051_sfr1_oc8051_dptr1_n21) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u18 ( .A0(dptr_hi[4]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[4]), .Y(oc8051_sfr1_oc8051_dptr1_n10) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u17 ( .B0(des2[4]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n10), .Y(
        oc8051_sfr1_oc8051_dptr1_n22) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u16 ( .A0(dptr_hi[5]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[5]), .Y(oc8051_sfr1_oc8051_dptr1_n9) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u15 ( .B0(des2[5]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n9), .Y(
        oc8051_sfr1_oc8051_dptr1_n23) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u14 ( .A0(dptr_hi[6]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[6]), .Y(oc8051_sfr1_oc8051_dptr1_n8) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u13 ( .B0(des2[6]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n8), .Y(
        oc8051_sfr1_oc8051_dptr1_n24) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u12 ( .A0(dptr_hi[7]), .A1(
        oc8051_sfr1_oc8051_dptr1_n6), .B0(oc8051_sfr1_oc8051_dptr1_n7), .B1(
        des_acc[7]), .Y(oc8051_sfr1_oc8051_dptr1_n5) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u11 ( .B0(des2[7]), .B1(
        oc8051_sfr1_oc8051_dptr1_n4), .A0N(oc8051_sfr1_oc8051_dptr1_n5), .Y(
        oc8051_sfr1_oc8051_dptr1_n25) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u10 ( .A1N(
        oc8051_sfr1_oc8051_dptr1_n2), .A0(oc8051_sfr1_oc8051_dptr1_n3), .B0(
        oc8051_sfr1_oc8051_dptr1_n4), .Y(oc8051_sfr1_oc8051_dptr1_n1) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u9 ( .A(des_acc[0]), .B(dptr_lo[0]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n26) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u8 ( .A(des_acc[1]), .B(dptr_lo[1]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n27) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u7 ( .A(des_acc[2]), .B(dptr_lo[2]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n28) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u6 ( .A(des_acc[3]), .B(dptr_lo[3]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n29) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u5 ( .A(des_acc[4]), .B(dptr_lo[4]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n30) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u4 ( .A(des_acc[5]), .B(dptr_lo[5]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n31) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u3 ( .A(des_acc[6]), .B(dptr_lo[6]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n32) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_dptr1_u2 ( .A(des_acc[7]), .B(dptr_lo[7]), .S0(oc8051_sfr1_oc8051_dptr1_n1), .Y(oc8051_sfr1_oc8051_dptr1_n33) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_0_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n18), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_1_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n19), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_2_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n20), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_3_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n21), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_4_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n22), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_5_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n23), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_6_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n24), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_hi_reg_7_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n25), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_hi[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_0_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n26), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_1_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n27), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_2_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n28), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_3_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n29), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_4_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n30), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_5_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n31), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_6_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n32), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_dptr1_data_lo_reg_7_ ( .D(
        oc8051_sfr1_oc8051_dptr1_n33), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        dptr_lo[7]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u51 ( .A(n_5_net_), .Y(
        oc8051_sfr1_oc8051_psw1_n40) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u50 ( .A(
        oc8051_sfr1_oc8051_psw1_n40), .B(wr_addr[5]), .C(wr_addr[3]), .Y(
        oc8051_sfr1_oc8051_psw1_n39) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u49 ( .A(wr_addr[6]), .B(wr_addr[4]), .C(wr_addr[7]), .D(oc8051_sfr1_oc8051_psw1_n39), .Y(
        oc8051_sfr1_oc8051_psw1_n37) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u48 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_psw1_n10) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u47 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_wr_bit_r), .C(wr_addr[2]), .Y(oc8051_sfr1_oc8051_psw1_n38)
         );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u46 ( .A(
        oc8051_sfr1_oc8051_psw1_n37), .B(oc8051_sfr1_oc8051_psw1_n10), .C(
        oc8051_sfr1_oc8051_psw1_n38), .Y(oc8051_sfr1_oc8051_psw1_n16) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u45 ( .A(wr_dat[3]), .B(
        oc8051_sfr1_psw_3_), .S0(oc8051_sfr1_oc8051_psw1_n16), .Y(bank_sel[0])
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u44 ( .A(wr_dat[4]), .B(
        oc8051_sfr1_psw_4_), .S0(oc8051_sfr1_oc8051_psw1_n16), .Y(bank_sel[1])
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u43 ( .A(oc8051_sfr1_oc8051_psw1_n16), .Y(oc8051_sfr1_oc8051_psw1_n7) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u42 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_psw1_n37), .Y(oc8051_sfr1_oc8051_psw1_n36) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u41 ( .A(oc8051_sfr1_oc8051_psw1_n36), .Y(oc8051_sfr1_oc8051_psw1_n24) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u40 ( .A(descy), .B(
        oc8051_sfr1_oc8051_psw1_n24), .Y(oc8051_sfr1_oc8051_psw1_n20) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u39 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_psw1_n8) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u38 ( .A(
        oc8051_sfr1_oc8051_psw1_n36), .B(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_psw1_n28) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u37 ( .A0(wr_addr[0]), .A1(
        oc8051_sfr1_oc8051_psw1_n8), .A2(oc8051_sfr1_oc8051_psw1_n28), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n35) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u36 ( .A(
        oc8051_sfr1_oc8051_psw1_n34), .B(oc8051_sfr1_psw_1_), .S0(
        oc8051_sfr1_oc8051_psw1_n35), .Y(oc8051_sfr1_oc8051_psw1_n43) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u35 ( .B0(wr_dat[2]), .B1(
        oc8051_sfr1_oc8051_psw1_n7), .A0N(oc8051_sfr1_oc8051_psw1_n20), .Y(
        oc8051_sfr1_oc8051_psw1_n31) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u34 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_psw1_n8), .Y(oc8051_sfr1_oc8051_psw1_n33) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u33 ( .A(oc8051_sfr1_oc8051_psw1_n7), .B(oc8051_sfr1_oc8051_psw1_n24), .Y(oc8051_sfr1_oc8051_psw1_n6) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u32 ( .A(oc8051_sfr1_oc8051_psw1_n6), .B(psw_set[1]), .Y(oc8051_sfr1_oc8051_psw1_n14) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u31 ( .A0(
        oc8051_sfr1_oc8051_psw1_n33), .A1(oc8051_sfr1_oc8051_psw1_n28), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .C0(oc8051_sfr1_oc8051_psw1_n14), .Y(
        oc8051_sfr1_oc8051_psw1_n32) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u30 ( .A(
        oc8051_sfr1_oc8051_psw1_n31), .B(oc8051_sfr1_psw_2_), .S0(
        oc8051_sfr1_oc8051_psw1_n32), .Y(oc8051_sfr1_oc8051_psw1_n29) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u29 ( .A(
        oc8051_sfr1_oc8051_psw1_n6), .B(psw_set[1]), .C(desov), .Y(
        oc8051_sfr1_oc8051_psw1_n30) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u28 ( .A(
        oc8051_sfr1_oc8051_psw1_n29), .B(oc8051_sfr1_oc8051_psw1_n30), .Y(
        oc8051_sfr1_oc8051_psw1_n44) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u27 ( .A(oc8051_sfr1_oc8051_psw1_n20), .Y(oc8051_sfr1_oc8051_psw1_n11) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u26 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_psw1_n7), .B0(oc8051_sfr1_oc8051_psw1_n11), .Y(
        oc8051_sfr1_oc8051_psw1_n25) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u25 ( .A(oc8051_sfr1_psw_3_), .Y(
        oc8051_sfr1_oc8051_psw1_n26) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u24 ( .A0(wr_addr[1]), .A1(
        wr_addr[0]), .A2(oc8051_sfr1_oc8051_psw1_n28), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n27) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u23 ( .A(
        oc8051_sfr1_oc8051_psw1_n25), .B(oc8051_sfr1_oc8051_psw1_n26), .S0(
        oc8051_sfr1_oc8051_psw1_n27), .Y(oc8051_sfr1_oc8051_psw1_n45) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u22 ( .A(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_psw1_n24), .Y(oc8051_sfr1_oc8051_psw1_n9) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u21 ( .A(oc8051_sfr1_oc8051_psw1_n9), .B(wr_addr[1]), .Y(oc8051_sfr1_oc8051_psw1_n19) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u20 ( .A(
        oc8051_sfr1_oc8051_psw1_n19), .B(oc8051_sfr1_oc8051_psw1_n10), .Y(
        oc8051_sfr1_oc8051_psw1_n21) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u19 ( .A(
        oc8051_sfr1_oc8051_psw1_n21), .B(oc8051_sfr1_psw_4_), .Y(
        oc8051_sfr1_oc8051_psw1_n23) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u18 ( .A(
        oc8051_sfr1_oc8051_psw1_n23), .B(wr_dat[4]), .S0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n22) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u17 ( .A0(
        oc8051_sfr1_oc8051_psw1_n21), .A1(oc8051_sfr1_oc8051_psw1_n20), .B0(
        oc8051_sfr1_oc8051_psw1_n22), .Y(oc8051_sfr1_oc8051_psw1_n46) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u16 ( .A0(
        oc8051_sfr1_oc8051_psw1_n19), .A1(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_psw1_n7), .Y(oc8051_sfr1_oc8051_psw1_n18) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u15 ( .A(
        oc8051_sfr1_oc8051_psw1_n17), .B(oc8051_sfr1_psw_5_), .S0(
        oc8051_sfr1_oc8051_psw1_n18), .Y(oc8051_sfr1_oc8051_psw1_n47) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u14 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_psw1_n7), .B0(desac), .B1(
        oc8051_sfr1_oc8051_psw1_n6), .C0(oc8051_sfr1_oc8051_psw1_n11), .Y(
        oc8051_sfr1_oc8051_psw1_n12) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u13 ( .A0(
        oc8051_sfr1_oc8051_psw1_n8), .A1(wr_addr[0]), .A2(
        oc8051_sfr1_oc8051_psw1_n9), .B0(oc8051_sfr1_oc8051_psw1_n16), .Y(
        oc8051_sfr1_oc8051_psw1_n15) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u12 ( .A0(psw_set[0]), .A1(
        oc8051_sfr1_oc8051_psw1_n14), .B0(oc8051_sfr1_oc8051_psw1_n15), .Y(
        oc8051_sfr1_oc8051_psw1_n13) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u11 ( .A(
        oc8051_sfr1_oc8051_psw1_n12), .B(oc8051_sfr1_oc8051_psw1_n1), .S0(
        oc8051_sfr1_oc8051_psw1_n13), .Y(oc8051_sfr1_oc8051_psw1_n48) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u10 ( .A0(
        oc8051_sfr1_oc8051_psw1_n6), .A1(descy), .B0(wr_dat[7]), .B1(
        oc8051_sfr1_oc8051_psw1_n7), .C0(oc8051_sfr1_oc8051_psw1_n11), .Y(
        oc8051_sfr1_oc8051_psw1_n2) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u9 ( .A(cy), .Y(
        oc8051_sfr1_oc8051_psw1_n3) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u8 ( .A(oc8051_sfr1_oc8051_psw1_n8), 
        .B(oc8051_sfr1_oc8051_psw1_n9), .C(oc8051_sfr1_oc8051_psw1_n10), .Y(
        oc8051_sfr1_oc8051_psw1_n5) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_psw1_u7 ( .A(oc8051_sfr1_oc8051_psw1_n5), 
        .B(oc8051_sfr1_oc8051_psw1_n6), .C(oc8051_sfr1_oc8051_psw1_n7), .Y(
        oc8051_sfr1_oc8051_psw1_n4) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u6 ( .A(oc8051_sfr1_oc8051_psw1_n2), .B(oc8051_sfr1_oc8051_psw1_n3), .S0(oc8051_sfr1_oc8051_psw1_n4), .Y(
        oc8051_sfr1_oc8051_psw1_n49) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_psw1_u5 ( .A(oc8051_sfr1_oc8051_psw1_n1), 
        .Y(srcac) );
  AO21B_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u4 ( .A0(wr_dat[5]), .A1(
        oc8051_sfr1_oc8051_psw1_n7), .B0N(oc8051_sfr1_oc8051_psw1_n20), .Y(
        oc8051_sfr1_oc8051_psw1_n17) );
  AO21B_X0P5M_A12TS oc8051_sfr1_oc8051_psw1_u3 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_psw1_n7), .B0N(oc8051_sfr1_oc8051_psw1_n20), .Y(
        oc8051_sfr1_oc8051_psw1_n34) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_6_ ( .D(
        oc8051_sfr1_oc8051_psw1_n48), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_psw1_n1) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_7_ ( .D(
        oc8051_sfr1_oc8051_psw1_n49), .CK(wb_clk_i), .R(wb_rst_i), .Q(cy) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_3_ ( .D(
        oc8051_sfr1_oc8051_psw1_n45), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_4_ ( .D(
        oc8051_sfr1_oc8051_psw1_n46), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_2_ ( .D(
        oc8051_sfr1_oc8051_psw1_n44), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_1_ ( .D(
        oc8051_sfr1_oc8051_psw1_n43), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_psw1_data_reg_5_ ( .D(
        oc8051_sfr1_oc8051_psw1_n47), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_psw_5_) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u171 ( .AN(oc8051_sfr1_wr_bit_r), .B(n_5_net_), .Y(oc8051_sfr1_oc8051_ports1_n48) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u170 ( .A(
        oc8051_sfr1_oc8051_ports1_n48), .Y(oc8051_sfr1_oc8051_ports1_n45) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u169 ( .A(wr_addr[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n81) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u168 ( .A(
        oc8051_sfr1_oc8051_ports1_n45), .B(oc8051_sfr1_oc8051_ports1_n81), .C(
        wr_addr[4]), .Y(oc8051_sfr1_oc8051_ports1_n82) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u167 ( .A(n_5_net_), .B(
        oc8051_sfr1_oc8051_ports1_n81), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u166 ( .A(
        oc8051_sfr1_oc8051_ports1_n85), .Y(oc8051_sfr1_oc8051_ports1_n88) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u165 ( .A(wr_addr[1]), .B(
        wr_addr[2]), .C(wr_addr[0]), .Y(oc8051_sfr1_oc8051_ports1_n43) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u164 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n43), .Y(
        oc8051_sfr1_oc8051_ports1_n103) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u163 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(descy), .Y(oc8051_sfr1_oc8051_ports1_n105) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u162 ( .A(
        oc8051_sfr1_oc8051_ports1_n105), .Y(oc8051_sfr1_oc8051_ports1_n86) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u161 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_ports1_n105), .Y(oc8051_sfr1_oc8051_ports1_n87)
         );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u160 ( .A0(wr_dat[0]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n40) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u159 ( .A(
        oc8051_sfr1_oc8051_ports1_n43), .Y(oc8051_sfr1_oc8051_ports1_n42) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u158 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n42), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n104) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u157 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n103), 
        .B0(oc8051_sfr1_oc8051_ports1_n40), .C0(oc8051_sfr1_oc8051_ports1_n104), .Y(oc8051_sfr1_oc8051_ports1_n132) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u156 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n91) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u155 ( .A(wr_addr[1]), .B(
        wr_addr[2]), .C(oc8051_sfr1_oc8051_ports1_n91), .Y(
        oc8051_sfr1_oc8051_ports1_n38) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u154 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n38), .Y(
        oc8051_sfr1_oc8051_ports1_n101) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u153 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n35) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u152 ( .A(
        oc8051_sfr1_oc8051_ports1_n38), .Y(oc8051_sfr1_oc8051_ports1_n37) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u151 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n37), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n102) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u150 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n101), 
        .B0(oc8051_sfr1_oc8051_ports1_n35), .C0(oc8051_sfr1_oc8051_ports1_n102), .Y(oc8051_sfr1_oc8051_ports1_n133) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u149 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n94) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u148 ( .A(wr_addr[0]), .B(
        wr_addr[2]), .C(oc8051_sfr1_oc8051_ports1_n94), .Y(
        oc8051_sfr1_oc8051_ports1_n33) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u147 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n33), .Y(
        oc8051_sfr1_oc8051_ports1_n99) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u146 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n30) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u145 ( .A(
        oc8051_sfr1_oc8051_ports1_n33), .Y(oc8051_sfr1_oc8051_ports1_n32) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u144 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n32), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n100) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u143 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n99), 
        .B0(oc8051_sfr1_oc8051_ports1_n30), .C0(oc8051_sfr1_oc8051_ports1_n100), .Y(oc8051_sfr1_oc8051_ports1_n134) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u142 ( .A(
        oc8051_sfr1_oc8051_ports1_n91), .B(wr_addr[2]), .C(
        oc8051_sfr1_oc8051_ports1_n94), .Y(oc8051_sfr1_oc8051_ports1_n28) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u141 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n28), .Y(
        oc8051_sfr1_oc8051_ports1_n97) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u140 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n25) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u139 ( .A(
        oc8051_sfr1_oc8051_ports1_n28), .Y(oc8051_sfr1_oc8051_ports1_n27) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u138 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n27), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n98) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u137 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n97), 
        .B0(oc8051_sfr1_oc8051_ports1_n25), .C0(oc8051_sfr1_oc8051_ports1_n98), 
        .Y(oc8051_sfr1_oc8051_ports1_n135) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u136 ( .A(
        oc8051_sfr1_oc8051_ports1_n91), .B(oc8051_sfr1_oc8051_ports1_n94), .C(
        wr_addr[2]), .Y(oc8051_sfr1_oc8051_ports1_n22) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u135 ( .A(
        oc8051_sfr1_oc8051_ports1_n22), .Y(oc8051_sfr1_oc8051_ports1_n23) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u134 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n23), .Y(
        oc8051_sfr1_oc8051_ports1_n95) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u133 ( .A0(wr_dat[4]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n20) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u132 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n22), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n96) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u131 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n95), 
        .B0(oc8051_sfr1_oc8051_ports1_n20), .C0(oc8051_sfr1_oc8051_ports1_n96), 
        .Y(oc8051_sfr1_oc8051_ports1_n136) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u130 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_ports1_n94), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u129 ( .A(
        oc8051_sfr1_oc8051_ports1_n17), .Y(oc8051_sfr1_oc8051_ports1_n18) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u128 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n18), .Y(
        oc8051_sfr1_oc8051_ports1_n92) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u127 ( .A0(wr_dat[5]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n15) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u126 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n17), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n93) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u125 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n92), 
        .B0(oc8051_sfr1_oc8051_ports1_n15), .C0(oc8051_sfr1_oc8051_ports1_n93), 
        .Y(oc8051_sfr1_oc8051_ports1_n137) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u124 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_ports1_n91), .C(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n12) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u123 ( .A(
        oc8051_sfr1_oc8051_ports1_n12), .Y(oc8051_sfr1_oc8051_ports1_n13) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u122 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n13), .Y(
        oc8051_sfr1_oc8051_ports1_n89) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u121 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n10) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u120 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n12), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n90) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u119 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n89), 
        .B0(oc8051_sfr1_oc8051_ports1_n10), .C0(oc8051_sfr1_oc8051_ports1_n90), 
        .Y(oc8051_sfr1_oc8051_ports1_n138) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u118 ( .A(wr_addr[1]), .B(
        wr_addr[0]), .C(wr_addr[2]), .Y(oc8051_sfr1_oc8051_ports1_n5) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u117 ( .A(
        oc8051_sfr1_oc8051_ports1_n5), .Y(oc8051_sfr1_oc8051_ports1_n8) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u116 ( .A(
        oc8051_sfr1_oc8051_ports1_n88), .B(oc8051_sfr1_oc8051_ports1_n8), .Y(
        oc8051_sfr1_oc8051_ports1_n83) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u115 ( .A0(wr_dat[7]), .A1(
        oc8051_sfr1_oc8051_ports1_n86), .B0(oc8051_sfr1_oc8051_ports1_n87), 
        .Y(oc8051_sfr1_oc8051_ports1_n3) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u114 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n5), .B0(
        oc8051_sfr1_oc8051_ports1_n85), .C0(p1_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n84) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u113 ( .A0(
        oc8051_sfr1_oc8051_ports1_n82), .A1(oc8051_sfr1_oc8051_ports1_n83), 
        .B0(oc8051_sfr1_oc8051_ports1_n3), .C0(oc8051_sfr1_oc8051_ports1_n84), 
        .Y(oc8051_sfr1_oc8051_ports1_n139) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u112 ( .A(p0_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n79) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u111 ( .A(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n44) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u110 ( .A(
        oc8051_sfr1_oc8051_ports1_n44), .B(oc8051_sfr1_oc8051_ports1_n81), .C(
        n_5_net_), .Y(oc8051_sfr1_oc8051_ports1_n66) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u109 ( .A0(
        oc8051_sfr1_oc8051_ports1_n42), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n80)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u108 ( .A(
        oc8051_sfr1_oc8051_ports1_n79), .B(oc8051_sfr1_oc8051_ports1_n40), 
        .S0(oc8051_sfr1_oc8051_ports1_n80), .Y(oc8051_sfr1_oc8051_ports1_n140)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u107 ( .A(p0_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n77) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u106 ( .A0(
        oc8051_sfr1_oc8051_ports1_n37), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n78)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u105 ( .A(
        oc8051_sfr1_oc8051_ports1_n77), .B(oc8051_sfr1_oc8051_ports1_n35), 
        .S0(oc8051_sfr1_oc8051_ports1_n78), .Y(oc8051_sfr1_oc8051_ports1_n141)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u104 ( .A(p0_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n75) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u103 ( .A0(
        oc8051_sfr1_oc8051_ports1_n32), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n76)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u102 ( .A(
        oc8051_sfr1_oc8051_ports1_n75), .B(oc8051_sfr1_oc8051_ports1_n30), 
        .S0(oc8051_sfr1_oc8051_ports1_n76), .Y(oc8051_sfr1_oc8051_ports1_n142)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u101 ( .A(p0_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n73) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u100 ( .A0(
        oc8051_sfr1_oc8051_ports1_n27), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n74)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u99 ( .A(
        oc8051_sfr1_oc8051_ports1_n73), .B(oc8051_sfr1_oc8051_ports1_n25), 
        .S0(oc8051_sfr1_oc8051_ports1_n74), .Y(oc8051_sfr1_oc8051_ports1_n143)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u98 ( .A(p0_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n71) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u97 ( .A0(
        oc8051_sfr1_oc8051_ports1_n22), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n72)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u96 ( .A(
        oc8051_sfr1_oc8051_ports1_n71), .B(oc8051_sfr1_oc8051_ports1_n20), 
        .S0(oc8051_sfr1_oc8051_ports1_n72), .Y(oc8051_sfr1_oc8051_ports1_n144)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u95 ( .A(p0_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n69) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u94 ( .A0(
        oc8051_sfr1_oc8051_ports1_n17), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n70)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u93 ( .A(
        oc8051_sfr1_oc8051_ports1_n69), .B(oc8051_sfr1_oc8051_ports1_n15), 
        .S0(oc8051_sfr1_oc8051_ports1_n70), .Y(oc8051_sfr1_oc8051_ports1_n145)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u92 ( .A(p0_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n67) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u91 ( .A0(
        oc8051_sfr1_oc8051_ports1_n12), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n68)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u90 ( .A(
        oc8051_sfr1_oc8051_ports1_n67), .B(oc8051_sfr1_oc8051_ports1_n10), 
        .S0(oc8051_sfr1_oc8051_ports1_n68), .Y(oc8051_sfr1_oc8051_ports1_n146)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u89 ( .A(p0_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n64) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u88 ( .A0(
        oc8051_sfr1_oc8051_ports1_n5), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n66), .Y(oc8051_sfr1_oc8051_ports1_n65)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u87 ( .A(
        oc8051_sfr1_oc8051_ports1_n64), .B(oc8051_sfr1_oc8051_ports1_n3), .S0(
        oc8051_sfr1_oc8051_ports1_n65), .Y(oc8051_sfr1_oc8051_ports1_n147) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u86 ( .A(p3_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n62) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u85 ( .A(wr_addr[5]), .B(
        n_5_net_), .C(wr_addr[4]), .Y(oc8051_sfr1_oc8051_ports1_n49) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u84 ( .A0(
        oc8051_sfr1_oc8051_ports1_n42), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n63)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u83 ( .A(
        oc8051_sfr1_oc8051_ports1_n62), .B(oc8051_sfr1_oc8051_ports1_n40), 
        .S0(oc8051_sfr1_oc8051_ports1_n63), .Y(oc8051_sfr1_oc8051_ports1_n148)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u82 ( .A(p3_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n60) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u81 ( .A0(
        oc8051_sfr1_oc8051_ports1_n37), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n61)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u80 ( .A(
        oc8051_sfr1_oc8051_ports1_n60), .B(oc8051_sfr1_oc8051_ports1_n35), 
        .S0(oc8051_sfr1_oc8051_ports1_n61), .Y(oc8051_sfr1_oc8051_ports1_n149)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u79 ( .A(p3_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n58) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u78 ( .A0(
        oc8051_sfr1_oc8051_ports1_n32), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n59)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u77 ( .A(
        oc8051_sfr1_oc8051_ports1_n58), .B(oc8051_sfr1_oc8051_ports1_n30), 
        .S0(oc8051_sfr1_oc8051_ports1_n59), .Y(oc8051_sfr1_oc8051_ports1_n150)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u76 ( .A(p3_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n56) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u75 ( .A0(
        oc8051_sfr1_oc8051_ports1_n27), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n57)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u74 ( .A(
        oc8051_sfr1_oc8051_ports1_n56), .B(oc8051_sfr1_oc8051_ports1_n25), 
        .S0(oc8051_sfr1_oc8051_ports1_n57), .Y(oc8051_sfr1_oc8051_ports1_n151)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u73 ( .A(p3_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n54) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u72 ( .A0(
        oc8051_sfr1_oc8051_ports1_n22), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n55)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u71 ( .A(
        oc8051_sfr1_oc8051_ports1_n54), .B(oc8051_sfr1_oc8051_ports1_n20), 
        .S0(oc8051_sfr1_oc8051_ports1_n55), .Y(oc8051_sfr1_oc8051_ports1_n152)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u70 ( .A(p3_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n52) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u69 ( .A0(
        oc8051_sfr1_oc8051_ports1_n17), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n53)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u68 ( .A(
        oc8051_sfr1_oc8051_ports1_n52), .B(oc8051_sfr1_oc8051_ports1_n15), 
        .S0(oc8051_sfr1_oc8051_ports1_n53), .Y(oc8051_sfr1_oc8051_ports1_n153)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u67 ( .A(p3_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n50) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u66 ( .A0(
        oc8051_sfr1_oc8051_ports1_n12), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n51)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u65 ( .A(
        oc8051_sfr1_oc8051_ports1_n50), .B(oc8051_sfr1_oc8051_ports1_n10), 
        .S0(oc8051_sfr1_oc8051_ports1_n51), .Y(oc8051_sfr1_oc8051_ports1_n154)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u64 ( .A(p3_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n46) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u63 ( .A0(
        oc8051_sfr1_oc8051_ports1_n5), .A1(oc8051_sfr1_oc8051_ports1_n48), 
        .B0(oc8051_sfr1_oc8051_ports1_n49), .Y(oc8051_sfr1_oc8051_ports1_n47)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u62 ( .A(
        oc8051_sfr1_oc8051_ports1_n46), .B(oc8051_sfr1_oc8051_ports1_n3), .S0(
        oc8051_sfr1_oc8051_ports1_n47), .Y(oc8051_sfr1_oc8051_ports1_n155) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u61 ( .A(wr_addr[5]), .B(
        oc8051_sfr1_oc8051_ports1_n44), .C(oc8051_sfr1_oc8051_ports1_n45), .Y(
        oc8051_sfr1_oc8051_ports1_n1) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u60 ( .A(n_5_net_), .B(
        oc8051_sfr1_oc8051_ports1_n44), .C(wr_addr[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n6) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_ports1_u59 ( .A(
        oc8051_sfr1_oc8051_ports1_n6), .Y(oc8051_sfr1_oc8051_ports1_n7) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u58 ( .A(
        oc8051_sfr1_oc8051_ports1_n43), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n39) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u57 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n42), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[0]), .Y(
        oc8051_sfr1_oc8051_ports1_n41) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u56 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n39), 
        .B0(oc8051_sfr1_oc8051_ports1_n40), .C0(oc8051_sfr1_oc8051_ports1_n41), 
        .Y(oc8051_sfr1_oc8051_ports1_n156) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u55 ( .A(
        oc8051_sfr1_oc8051_ports1_n38), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n34) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u54 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n37), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[1]), .Y(
        oc8051_sfr1_oc8051_ports1_n36) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u53 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n34), 
        .B0(oc8051_sfr1_oc8051_ports1_n35), .C0(oc8051_sfr1_oc8051_ports1_n36), 
        .Y(oc8051_sfr1_oc8051_ports1_n157) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u52 ( .A(
        oc8051_sfr1_oc8051_ports1_n33), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n29) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u51 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n32), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[2]), .Y(
        oc8051_sfr1_oc8051_ports1_n31) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u50 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n29), 
        .B0(oc8051_sfr1_oc8051_ports1_n30), .C0(oc8051_sfr1_oc8051_ports1_n31), 
        .Y(oc8051_sfr1_oc8051_ports1_n158) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u49 ( .A(
        oc8051_sfr1_oc8051_ports1_n28), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n24) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u48 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n27), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[3]), .Y(
        oc8051_sfr1_oc8051_ports1_n26) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u47 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n24), 
        .B0(oc8051_sfr1_oc8051_ports1_n25), .C0(oc8051_sfr1_oc8051_ports1_n26), 
        .Y(oc8051_sfr1_oc8051_ports1_n159) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u46 ( .A(
        oc8051_sfr1_oc8051_ports1_n23), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n19) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u45 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n22), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[4]), .Y(
        oc8051_sfr1_oc8051_ports1_n21) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u44 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n19), 
        .B0(oc8051_sfr1_oc8051_ports1_n20), .C0(oc8051_sfr1_oc8051_ports1_n21), 
        .Y(oc8051_sfr1_oc8051_ports1_n160) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u43 ( .A(
        oc8051_sfr1_oc8051_ports1_n18), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n14) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u42 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n17), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[5]), .Y(
        oc8051_sfr1_oc8051_ports1_n16) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u41 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n14), 
        .B0(oc8051_sfr1_oc8051_ports1_n15), .C0(oc8051_sfr1_oc8051_ports1_n16), 
        .Y(oc8051_sfr1_oc8051_ports1_n161) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u40 ( .A(
        oc8051_sfr1_oc8051_ports1_n13), .B(oc8051_sfr1_oc8051_ports1_n7), .Y(
        oc8051_sfr1_oc8051_ports1_n9) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u39 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n12), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[6]), .Y(
        oc8051_sfr1_oc8051_ports1_n11) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u38 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n9), .B0(
        oc8051_sfr1_oc8051_ports1_n10), .C0(oc8051_sfr1_oc8051_ports1_n11), 
        .Y(oc8051_sfr1_oc8051_ports1_n162) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_ports1_u37 ( .A(
        oc8051_sfr1_oc8051_ports1_n7), .B(oc8051_sfr1_oc8051_ports1_n8), .Y(
        oc8051_sfr1_oc8051_ports1_n2) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u36 ( .A0(
        oc8051_sfr1_wr_bit_r), .A1(oc8051_sfr1_oc8051_ports1_n5), .B0(
        oc8051_sfr1_oc8051_ports1_n6), .C0(p2_o[7]), .Y(
        oc8051_sfr1_oc8051_ports1_n4) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u35 ( .A0(
        oc8051_sfr1_oc8051_ports1_n1), .A1(oc8051_sfr1_oc8051_ports1_n2), .B0(
        oc8051_sfr1_oc8051_ports1_n3), .C0(oc8051_sfr1_oc8051_ports1_n4), .Y(
        oc8051_sfr1_oc8051_ports1_n163) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u34 ( .A(p0_i[0]), .B(p0_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u33 ( .A(p0_i[1]), .B(p0_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u32 ( .A(p0_i[2]), .B(p0_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u31 ( .A(p0_i[3]), .B(p0_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u30 ( .A(p0_i[4]), .B(p0_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u29 ( .A(p0_i[5]), .B(p0_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u28 ( .A(p0_i[6]), .B(p0_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u27 ( .A(p0_i[7]), .B(p0_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p0_data_7_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u26 ( .A(p1_i[0]), .B(p1_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u25 ( .A(p1_i[1]), .B(p1_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u24 ( .A(p1_i[2]), .B(p1_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u23 ( .A(p1_i[3]), .B(p1_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u22 ( .A(p1_i[4]), .B(p1_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u21 ( .A(p1_i[5]), .B(p1_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u20 ( .A(p1_i[6]), .B(p1_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u19 ( .A(p1_i[7]), .B(p1_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p1_data_7_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u18 ( .A(p2_i[0]), .B(p2_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u17 ( .A(p2_i[1]), .B(p2_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u16 ( .A(p2_i[2]), .B(p2_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u15 ( .A(p2_i[3]), .B(p2_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u14 ( .A(p2_i[4]), .B(p2_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u13 ( .A(p2_i[5]), .B(p2_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u12 ( .A(p2_i[6]), .B(p2_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u11 ( .A(p2_i[7]), .B(p2_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p2_data_7_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u10 ( .A(p3_i[0]), .B(p3_o[0]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_0_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u9 ( .A(p3_i[1]), .B(p3_o[1]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_1_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u8 ( .A(p3_i[2]), .B(p3_o[2]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_2_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u7 ( .A(p3_i[3]), .B(p3_o[3]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_3_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u6 ( .A(p3_i[4]), .B(p3_o[4]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_4_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u5 ( .A(p3_i[5]), .B(p3_o[5]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_5_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u4 ( .A(p3_i[6]), .B(p3_o[6]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_6_) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_u3 ( .A(p3_i[7]), .B(p3_o[7]), 
        .S0(rmw), .Y(oc8051_sfr1_p3_data_7_) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_ports1_u2 ( .A(wb_rst_i), .Y(
        oc8051_sfr1_oc8051_ports1_n106) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n140), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n141), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n142), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n143), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n144), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n145), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n146), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p0_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n147), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p0_o[7]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n148), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n149), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n150), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n151), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n152), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n153), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n154), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p3_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n155), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p3_o[7]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n132), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n133), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n134), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n135), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n136), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n137), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n138), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p1_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n139), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p1_o[7]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_0_ ( .D(
        oc8051_sfr1_oc8051_ports1_n156), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[0]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_1_ ( .D(
        oc8051_sfr1_oc8051_ports1_n157), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[1]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_2_ ( .D(
        oc8051_sfr1_oc8051_ports1_n158), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[2]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_3_ ( .D(
        oc8051_sfr1_oc8051_ports1_n159), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[3]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_4_ ( .D(
        oc8051_sfr1_oc8051_ports1_n160), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[4]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_5_ ( .D(
        oc8051_sfr1_oc8051_ports1_n161), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[5]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_6_ ( .D(
        oc8051_sfr1_oc8051_ports1_n162), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[6]) );
  DFFSQ_X0P5M_A12TS oc8051_sfr1_oc8051_ports1_p2_out_reg_7_ ( .D(
        oc8051_sfr1_oc8051_ports1_n163), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_ports1_n106), .Q(p2_o[7]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u241 ( .A(oc8051_sfr1_pcon[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n164) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u240 ( .A(oc8051_sfr1_scon_6_), .Y(
        oc8051_sfr1_oc8051_uatr1_n36) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u239 ( .A(
        oc8051_sfr1_oc8051_uatr1_n205), .Y(oc8051_sfr1_oc8051_uatr1_n168) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u238 ( .A(oc8051_sfr1_tf1), .Y(
        oc8051_sfr1_oc8051_uatr1_n169) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u237 ( .A(
        oc8051_sfr1_oc8051_uatr1_n168), .B(oc8051_sfr1_oc8051_uatr1_n169), .Y(
        oc8051_sfr1_oc8051_uatr1_n166) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u236 ( .A(
        oc8051_sfr1_oc8051_uatr1_n166), .B(oc8051_sfr1_brate2), .S0(
        oc8051_sfr1_tclk), .Y(oc8051_sfr1_oc8051_uatr1_n167) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u235 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n36), .A1(oc8051_sfr1_scon_7_), .B0(
        oc8051_sfr1_oc8051_uatr1_n167), .Y(oc8051_sfr1_oc8051_uatr1_n8) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u234 ( .A1N(
        oc8051_sfr1_oc8051_uatr1_smod_clk_tr), .A0(
        oc8051_sfr1_oc8051_uatr1_n164), .B0(oc8051_sfr1_oc8051_uatr1_n8), .Y(
        oc8051_sfr1_oc8051_uatr1_n174) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u233 ( .A(
        oc8051_sfr1_oc8051_uatr1_n166), .B(oc8051_sfr1_brate2), .S0(
        oc8051_sfr1_rclk), .Y(oc8051_sfr1_oc8051_uatr1_n165) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u232 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n36), .A1(oc8051_sfr1_scon_7_), .B0(
        oc8051_sfr1_oc8051_uatr1_n165), .Y(oc8051_sfr1_oc8051_uatr1_n94) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u231 ( .A1N(
        oc8051_sfr1_oc8051_uatr1_smod_clk_re), .A0(
        oc8051_sfr1_oc8051_uatr1_n164), .B0(oc8051_sfr1_oc8051_uatr1_n94), .Y(
        oc8051_sfr1_oc8051_uatr1_n269) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u230 ( .A(oc8051_sfr1_scon_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n120) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u229 ( .A(
        oc8051_sfr1_oc8051_uatr1_n180), .B(oc8051_sfr1_oc8051_uatr1_n120), .Y(
        oc8051_sfr1_uart_int) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u228 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_), .B(oc8051_sfr1_sbuf[7]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n181) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u227 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_), .B(oc8051_sfr1_sbuf[6]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n182) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u226 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_), .B(oc8051_sfr1_sbuf[5]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n183) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u225 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_), .B(oc8051_sfr1_sbuf[4]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n184) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u224 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_), .B(oc8051_sfr1_sbuf[3]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n185) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u223 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_), .B(oc8051_sfr1_sbuf[2]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n186) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u222 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_), .B(oc8051_sfr1_sbuf[1]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n187) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u221 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_), .B(oc8051_sfr1_sbuf[0]), 
        .S0(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n188) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u220 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_uatr1_n28) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u219 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_uatr1_n27) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u218 ( .A(
        oc8051_sfr1_oc8051_uatr1_n28), .B(oc8051_sfr1_oc8051_uatr1_n27), .Y(
        oc8051_sfr1_oc8051_uatr1_n22) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u217 ( .A(wr_addr[6]), .B(
        wr_addr[5]), .Y(oc8051_sfr1_oc8051_uatr1_n163) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u216 ( .A(wr_addr[7]), .B(n_5_net_), .C(oc8051_sfr1_oc8051_uatr1_n163), .Y(oc8051_sfr1_oc8051_uatr1_n132) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u215 ( .A(wr_addr[3]), .B(
        oc8051_sfr1_wr_bit_r), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_uatr1_n162) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u214 ( .A(oc8051_sfr1_pcon[0]), 
        .B(wr_dat[0]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n190) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u213 ( .A(oc8051_sfr1_pcon[1]), 
        .B(wr_dat[1]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n191) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u212 ( .A(oc8051_sfr1_pcon[2]), 
        .B(wr_dat[2]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n192) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u211 ( .A(oc8051_sfr1_pcon[3]), 
        .B(wr_dat[3]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n193) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u210 ( .A(oc8051_sfr1_pcon[4]), 
        .B(wr_dat[4]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n194) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u209 ( .A(oc8051_sfr1_pcon[5]), 
        .B(wr_dat[5]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n195) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u208 ( .A(oc8051_sfr1_pcon[6]), 
        .B(wr_dat[6]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n196) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u207 ( .A(oc8051_sfr1_pcon[7]), 
        .B(wr_dat[7]), .S0(oc8051_sfr1_oc8051_uatr1_n161), .Y(
        oc8051_sfr1_oc8051_uatr1_n197) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u206 ( .A(oc8051_sfr1_scon_7_), .Y(
        oc8051_sfr1_oc8051_uatr1_n40) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u205 ( .A(
        oc8051_sfr1_oc8051_uatr1_n36), .B(oc8051_sfr1_oc8051_uatr1_n40), .Y(
        oc8051_sfr1_oc8051_uatr1_n91) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u204 ( .A(
        oc8051_sfr1_oc8051_uatr1_receive), .B(oc8051_sfr1_oc8051_uatr1_n91), 
        .C(oc8051_sfr1_oc8051_uatr1_shift_re), .Y(
        oc8051_sfr1_oc8051_uatr1_n150) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u203 ( .A(
        oc8051_sfr1_oc8051_uatr1_n150), .Y(oc8051_sfr1_oc8051_uatr1_n143) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u202 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_done), .B(oc8051_sfr1_oc8051_uatr1_n143), 
        .Y(oc8051_sfr1_oc8051_uatr1_n98) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u201 ( .A(
        oc8051_sfr1_oc8051_uatr1_n98), .Y(oc8051_sfr1_oc8051_uatr1_n104) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u200 ( .A(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .B(
        oc8051_sfr1_oc8051_uatr1_n104), .C(
        oc8051_sfr1_oc8051_uatr1_re_count_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n111) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u199 ( .A(
        oc8051_sfr1_oc8051_uatr1_n91), .Y(oc8051_sfr1_oc8051_uatr1_n79) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u198 ( .A(oc8051_sfr1_pres_ow), 
        .B(oc8051_sfr1_oc8051_uatr1_n79), .C(oc8051_sfr1_oc8051_uatr1_receive), 
        .Y(oc8051_sfr1_oc8051_uatr1_n106) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u197 ( .A(
        oc8051_sfr1_oc8051_uatr1_n106), .Y(oc8051_sfr1_oc8051_uatr1_n109) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u196 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_done), .Y(oc8051_sfr1_oc8051_uatr1_n130)
         );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u195 ( .A(
        oc8051_sfr1_oc8051_uatr1_n109), .B(oc8051_sfr1_oc8051_uatr1_n143), .C(
        oc8051_sfr1_oc8051_uatr1_n130), .Y(oc8051_sfr1_oc8051_uatr1_n140) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u194 ( .A(
        oc8051_sfr1_oc8051_uatr1_n140), .B(oc8051_sfr1_oc8051_uatr1_shift_re), 
        .C(oc8051_sfr1_scon_4_), .D(oc8051_sfr1_oc8051_uatr1_n91), .Y(
        oc8051_sfr1_oc8051_uatr1_n151) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u193 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n140), .B(oc8051_sfr1_oc8051_uatr1_n91), .Y(
        oc8051_sfr1_oc8051_uatr1_n138) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u192 ( .A(oc8051_sfr1_scon_0_), 
        .B(oc8051_sfr1_oc8051_uatr1_receive), .Y(oc8051_sfr1_oc8051_uatr1_n136) );
  AOI32_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u191 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n138), .A1(oc8051_sfr1_scon_4_), .A2(
        oc8051_sfr1_oc8051_uatr1_n136), .B0(oc8051_sfr1_oc8051_uatr1_n109), 
        .B1(oc8051_sfr1_oc8051_uatr1_rx_done), .Y(
        oc8051_sfr1_oc8051_uatr1_n160) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u190 ( .A(
        oc8051_sfr1_oc8051_uatr1_n111), .B(oc8051_sfr1_oc8051_uatr1_n151), .C(
        oc8051_sfr1_oc8051_uatr1_n160), .Y(oc8051_sfr1_oc8051_uatr1_n103) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u189 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_), .Y(
        oc8051_sfr1_oc8051_uatr1_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u188 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_), .Y(
        oc8051_sfr1_oc8051_uatr1_n101) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u187 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n104), .A1(oc8051_sfr1_oc8051_uatr1_n109), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .Y(oc8051_sfr1_oc8051_uatr1_n107)
         );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u186 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n103), .A1(oc8051_sfr1_oc8051_uatr1_n159), 
        .B0(oc8051_sfr1_oc8051_uatr1_n101), .B1(oc8051_sfr1_oc8051_uatr1_n107), 
        .Y(oc8051_sfr1_oc8051_uatr1_n206) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u185 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_), .Y(
        oc8051_sfr1_oc8051_uatr1_n158) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u184 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_), .Y(
        oc8051_sfr1_oc8051_uatr1_n157) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u183 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n158), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .B1(oc8051_sfr1_oc8051_uatr1_n157), 
        .C0(oc8051_sfr1_oc8051_uatr1_n151), .Y(oc8051_sfr1_oc8051_uatr1_n207)
         );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u182 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n103), .A1(oc8051_sfr1_oc8051_uatr1_n158), 
        .B0(oc8051_sfr1_oc8051_uatr1_n107), .B1(oc8051_sfr1_oc8051_uatr1_n159), 
        .Y(oc8051_sfr1_oc8051_uatr1_n208) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u181 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_), .Y(
        oc8051_sfr1_oc8051_uatr1_n156) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u180 ( .A(
        oc8051_sfr1_oc8051_uatr1_n151), .Y(oc8051_sfr1_oc8051_uatr1_n137) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u179 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n138), .A1(oc8051_sfr1_oc8051_uatr1_n137), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .Y(oc8051_sfr1_oc8051_uatr1_n108)
         );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u178 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n157), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .B1(oc8051_sfr1_oc8051_uatr1_n156), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n209)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u177 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_), .Y(
        oc8051_sfr1_oc8051_uatr1_n155) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u176 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n156), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .B1(oc8051_sfr1_oc8051_uatr1_n155), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n210)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u175 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_), .Y(
        oc8051_sfr1_oc8051_uatr1_n154) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u174 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n155), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .B1(oc8051_sfr1_oc8051_uatr1_n154), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n211)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u173 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_), .Y(
        oc8051_sfr1_oc8051_uatr1_n153) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u172 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n154), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .B1(oc8051_sfr1_oc8051_uatr1_n153), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n212)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u171 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n152) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u170 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n153), 
        .B0(oc8051_sfr1_oc8051_uatr1_n103), .B1(oc8051_sfr1_oc8051_uatr1_n152), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n213)
         );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u169 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n107), .A1(oc8051_sfr1_oc8051_uatr1_n152), 
        .B0(oc8051_sfr1_oc8051_uatr1_n202), .B1(oc8051_sfr1_oc8051_uatr1_n103), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n214)
         );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u168 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n202), .A1(oc8051_sfr1_oc8051_uatr1_n107), 
        .B0(oc8051_sfr1_oc8051_uatr1_n203), .B1(oc8051_sfr1_oc8051_uatr1_n103), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n215)
         );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u167 ( .A(
        oc8051_sfr1_oc8051_uatr1_n151), .B(oc8051_sfr1_oc8051_uatr1_n98), .Y(
        oc8051_sfr1_oc8051_uatr1_n142) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u166 ( .A(
        oc8051_sfr1_oc8051_uatr1_n143), .B(oc8051_sfr1_oc8051_uatr1_n142), .C(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n144) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u165 ( .A(
        oc8051_sfr1_oc8051_uatr1_n144), .B(
        oc8051_sfr1_oc8051_uatr1_re_count_1_), .C(
        oc8051_sfr1_oc8051_uatr1_re_count_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n148) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u164 ( .A0(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .A1(
        oc8051_sfr1_oc8051_uatr1_n150), .B0(oc8051_sfr1_oc8051_uatr1_n142), 
        .Y(oc8051_sfr1_oc8051_uatr1_n145) );
  AOI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u163 ( .A1N(
        oc8051_sfr1_oc8051_uatr1_re_count_1_), .A0(
        oc8051_sfr1_oc8051_uatr1_n143), .B0(oc8051_sfr1_oc8051_uatr1_n145), 
        .Y(oc8051_sfr1_oc8051_uatr1_n147) );
  OA21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u162 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n150), .A1(
        oc8051_sfr1_oc8051_uatr1_re_count_2_), .B0(
        oc8051_sfr1_oc8051_uatr1_n147), .Y(oc8051_sfr1_oc8051_uatr1_n149) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u161 ( .A(
        oc8051_sfr1_oc8051_uatr1_n148), .B(oc8051_sfr1_oc8051_uatr1_n149), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n216) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u160 ( .A(
        oc8051_sfr1_oc8051_uatr1_n144), .B(
        oc8051_sfr1_oc8051_uatr1_re_count_1_), .Y(
        oc8051_sfr1_oc8051_uatr1_n146) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u159 ( .A(
        oc8051_sfr1_oc8051_uatr1_n146), .B(oc8051_sfr1_oc8051_uatr1_n147), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n217) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u158 ( .A(
        oc8051_sfr1_oc8051_uatr1_n144), .B(oc8051_sfr1_oc8051_uatr1_n145), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_1_), .Y(
        oc8051_sfr1_oc8051_uatr1_n218) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u157 ( .A(
        oc8051_sfr1_oc8051_uatr1_n143), .B(oc8051_sfr1_oc8051_uatr1_n142), .Y(
        oc8051_sfr1_oc8051_uatr1_n141) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u156 ( .A(
        oc8051_sfr1_oc8051_uatr1_n141), .B(oc8051_sfr1_oc8051_uatr1_n142), 
        .S0(oc8051_sfr1_oc8051_uatr1_re_count_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n219) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u155 ( .A(oc8051_sfr1_scon_4_), .Y(
        oc8051_sfr1_oc8051_uatr1_n26) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u154 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n91), .A1(oc8051_sfr1_oc8051_uatr1_n26), .A2(
        oc8051_sfr1_oc8051_uatr1_n140), .B0(oc8051_sfr1_oc8051_uatr1_n137), 
        .Y(oc8051_sfr1_oc8051_uatr1_n139) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u153 ( .A(rxd_i), .B(
        oc8051_sfr1_oc8051_uatr1_rxd_r), .S0(oc8051_sfr1_oc8051_uatr1_n139), 
        .Y(oc8051_sfr1_oc8051_uatr1_n220) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u152 ( .A(rxd_i), .Y(
        oc8051_sfr1_oc8051_uatr1_n96) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u151 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n137), .A1(oc8051_sfr1_oc8051_uatr1_n96), 
        .A2(oc8051_sfr1_oc8051_uatr1_rxd_r), .B0(oc8051_sfr1_oc8051_uatr1_n138), .Y(oc8051_sfr1_oc8051_uatr1_n133) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u150 ( .A(
        oc8051_sfr1_oc8051_uatr1_receive), .Y(oc8051_sfr1_oc8051_uatr1_n134)
         );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u149 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n136), .A1(oc8051_sfr1_scon_4_), .B0(
        oc8051_sfr1_oc8051_uatr1_n130), .C0(oc8051_sfr1_oc8051_uatr1_n137), 
        .Y(oc8051_sfr1_oc8051_uatr1_n135) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u148 ( .A(
        oc8051_sfr1_oc8051_uatr1_n133), .B(oc8051_sfr1_oc8051_uatr1_n134), 
        .S0(oc8051_sfr1_oc8051_uatr1_n135), .Y(oc8051_sfr1_oc8051_uatr1_n221)
         );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u147 ( .A(wr_addr[3]), .B(
        oc8051_sfr1_oc8051_uatr1_n132), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_uatr1_n131) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u146 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_uatr1_n131), .Y(oc8051_sfr1_oc8051_uatr1_n42) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u145 ( .A(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_uatr1_n41) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u144 ( .AN(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_uatr1_n131), .C(oc8051_sfr1_oc8051_uatr1_n28), 
        .D(oc8051_sfr1_oc8051_uatr1_n41), .Y(oc8051_sfr1_oc8051_uatr1_n92) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u143 ( .A(
        oc8051_sfr1_oc8051_uatr1_n92), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_uatr1_n20) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u142 ( .A(
        oc8051_sfr1_oc8051_uatr1_n20), .Y(oc8051_sfr1_oc8051_uatr1_n118) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u141 ( .A(
        oc8051_sfr1_oc8051_uatr1_n198), .B(oc8051_sfr1_oc8051_uatr1_n42), .C(
        oc8051_sfr1_oc8051_uatr1_n118), .D(oc8051_sfr1_oc8051_uatr1_n130), .Y(
        oc8051_sfr1_oc8051_uatr1_n122) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u140 ( .A(
        oc8051_sfr1_oc8051_uatr1_n42), .Y(oc8051_sfr1_oc8051_uatr1_n129) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u139 ( .A(descy), .B(
        oc8051_sfr1_oc8051_uatr1_n129), .Y(oc8051_sfr1_oc8051_uatr1_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u138 ( .A(
        oc8051_sfr1_oc8051_uatr1_n17), .Y(oc8051_sfr1_oc8051_uatr1_n116) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u137 ( .A0(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_), .A1(
        oc8051_sfr1_oc8051_uatr1_n122), .B0(oc8051_sfr1_oc8051_uatr1_n20), 
        .B1(wr_dat[2]), .C0(oc8051_sfr1_oc8051_uatr1_n116), .Y(
        oc8051_sfr1_oc8051_uatr1_n125) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u136 ( .A(oc8051_sfr1_scon_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n126) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u135 ( .A(
        oc8051_sfr1_oc8051_uatr1_n129), .B(oc8051_sfr1_oc8051_uatr1_n41), .Y(
        oc8051_sfr1_oc8051_uatr1_n21) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u134 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n21), .A1(wr_addr[0]), .A2(
        oc8051_sfr1_oc8051_uatr1_n28), .B0(oc8051_sfr1_oc8051_uatr1_n118), .Y(
        oc8051_sfr1_oc8051_uatr1_n128) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u133 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n122), .A1(oc8051_sfr1_oc8051_uatr1_n91), 
        .B0(oc8051_sfr1_oc8051_uatr1_n128), .Y(oc8051_sfr1_oc8051_uatr1_n127)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u132 ( .A(
        oc8051_sfr1_oc8051_uatr1_n125), .B(oc8051_sfr1_oc8051_uatr1_n126), 
        .S0(oc8051_sfr1_oc8051_uatr1_n127), .Y(oc8051_sfr1_oc8051_uatr1_n222)
         );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u131 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n20), .A1(wr_dat[0]), .B0(
        oc8051_sfr1_oc8051_uatr1_n116), .C0(oc8051_sfr1_oc8051_uatr1_n122), 
        .Y(oc8051_sfr1_oc8051_uatr1_n119) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u130 ( .A(
        oc8051_sfr1_oc8051_uatr1_n91), .B(oc8051_sfr1_oc8051_uatr1_n101), .C(
        oc8051_sfr1_scon_5_), .Y(oc8051_sfr1_oc8051_uatr1_n123) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u129 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n21), .A1(wr_addr[1]), .A2(wr_addr[0]), .B0(
        oc8051_sfr1_oc8051_uatr1_n118), .Y(oc8051_sfr1_oc8051_uatr1_n124) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u128 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n122), .A1(oc8051_sfr1_oc8051_uatr1_n123), 
        .B0(oc8051_sfr1_oc8051_uatr1_n124), .Y(oc8051_sfr1_oc8051_uatr1_n121)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u127 ( .A(
        oc8051_sfr1_oc8051_uatr1_n119), .B(oc8051_sfr1_oc8051_uatr1_n120), 
        .S0(oc8051_sfr1_oc8051_uatr1_n121), .Y(oc8051_sfr1_oc8051_uatr1_n223)
         );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u126 ( .A(wr_dat[1]), .B(
        oc8051_sfr1_oc8051_uatr1_n42), .S0(oc8051_sfr1_oc8051_uatr1_n118), .Y(
        oc8051_sfr1_oc8051_uatr1_n117) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u125 ( .A(
        oc8051_sfr1_oc8051_uatr1_n116), .B(oc8051_sfr1_oc8051_uatr1_n117), .Y(
        oc8051_sfr1_oc8051_uatr1_n112) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u124 ( .A(
        oc8051_sfr1_oc8051_uatr1_n198), .Y(oc8051_sfr1_oc8051_uatr1_n114) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u123 ( .A(
        oc8051_sfr1_oc8051_uatr1_n21), .B(wr_addr[1]), .C(
        oc8051_sfr1_oc8051_uatr1_n27), .Y(oc8051_sfr1_oc8051_uatr1_n115) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u122 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n42), .A1(oc8051_sfr1_oc8051_uatr1_n114), 
        .B0(oc8051_sfr1_oc8051_uatr1_n20), .C0(oc8051_sfr1_oc8051_uatr1_n115), 
        .Y(oc8051_sfr1_oc8051_uatr1_n113) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u121 ( .A(
        oc8051_sfr1_oc8051_uatr1_n112), .B(oc8051_sfr1_oc8051_uatr1_n180), 
        .S0(oc8051_sfr1_oc8051_uatr1_n113), .Y(oc8051_sfr1_oc8051_uatr1_n224)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u120 ( .A(
        oc8051_sfr1_oc8051_uatr1_n111), .Y(oc8051_sfr1_oc8051_uatr1_n110) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u119 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n109), .A1(oc8051_sfr1_oc8051_uatr1_n110), 
        .B0(oc8051_sfr1_oc8051_uatr1_rx_done), .C0(
        oc8051_sfr1_oc8051_uatr1_n204), .Y(oc8051_sfr1_oc8051_uatr1_n225) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u118 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n203), .A1(oc8051_sfr1_oc8051_uatr1_n107), 
        .B0(oc8051_sfr1_oc8051_uatr1_n204), .B1(oc8051_sfr1_oc8051_uatr1_n103), 
        .C0(oc8051_sfr1_oc8051_uatr1_n108), .Y(oc8051_sfr1_oc8051_uatr1_n226)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u117 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_sam_1_), .Y(oc8051_sfr1_oc8051_uatr1_n99)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u116 ( .A(
        oc8051_sfr1_oc8051_uatr1_rx_sam_0_), .Y(oc8051_sfr1_oc8051_uatr1_n95)
         );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u115 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n99), .A1(oc8051_sfr1_oc8051_uatr1_n95), .B0(
        oc8051_sfr1_oc8051_uatr1_n98), .C0(oc8051_sfr1_oc8051_uatr1_n106), .Y(
        oc8051_sfr1_oc8051_uatr1_n105) );
  AOI32_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u114 ( .A0(
        oc8051_sfr1_oc8051_uatr1_rx_sam_0_), .A1(oc8051_sfr1_oc8051_uatr1_n104), .A2(oc8051_sfr1_oc8051_uatr1_rx_sam_1_), .B0(rxd_i), .B1(
        oc8051_sfr1_oc8051_uatr1_n105), .Y(oc8051_sfr1_oc8051_uatr1_n102) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u113 ( .A(
        oc8051_sfr1_oc8051_uatr1_n101), .B(oc8051_sfr1_oc8051_uatr1_n102), 
        .S0(oc8051_sfr1_oc8051_uatr1_n103), .Y(oc8051_sfr1_oc8051_uatr1_n227)
         );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u112 ( .A(
        oc8051_sfr1_oc8051_uatr1_re_count_0_), .B(oc8051_sfr1_oc8051_uatr1_n98), .Y(oc8051_sfr1_oc8051_uatr1_n100) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u111 ( .A(
        oc8051_sfr1_oc8051_uatr1_n99), .B(oc8051_sfr1_oc8051_uatr1_n96), .S0(
        oc8051_sfr1_oc8051_uatr1_n100), .Y(oc8051_sfr1_oc8051_uatr1_n228) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u110 ( .A(
        oc8051_sfr1_oc8051_uatr1_re_count_3_), .B(oc8051_sfr1_oc8051_uatr1_n98), .Y(oc8051_sfr1_oc8051_uatr1_n97) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u109 ( .A(
        oc8051_sfr1_oc8051_uatr1_n95), .B(oc8051_sfr1_oc8051_uatr1_n96), .S0(
        oc8051_sfr1_oc8051_uatr1_n97), .Y(oc8051_sfr1_oc8051_uatr1_n229) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u108 ( .A(
        oc8051_sfr1_oc8051_uatr1_n94), .B(oc8051_sfr1_pcon[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n93) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u107 ( .A(
        oc8051_sfr1_oc8051_uatr1_smod_clk_re), .B(oc8051_sfr1_oc8051_uatr1_n93), .Y(oc8051_sfr1_oc8051_uatr1_n230) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u106 ( .A(
        oc8051_sfr1_oc8051_uatr1_n27), .B(oc8051_sfr1_oc8051_uatr1_n92), .Y(
        oc8051_sfr1_oc8051_uatr1_n61) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u105 ( .A(
        oc8051_sfr1_oc8051_uatr1_n61), .Y(oc8051_sfr1_oc8051_uatr1_n43) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u104 ( .A(
        oc8051_sfr1_oc8051_uatr1_trans), .B(oc8051_sfr1_oc8051_uatr1_n43), .Y(
        oc8051_sfr1_oc8051_uatr1_n11) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u103 ( .A(
        oc8051_sfr1_oc8051_uatr1_n11), .Y(oc8051_sfr1_oc8051_uatr1_n87) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u102 ( .A(
        oc8051_sfr1_oc8051_uatr1_n87), .B(oc8051_sfr1_oc8051_uatr1_n91), .C(
        oc8051_sfr1_oc8051_uatr1_shift_tr), .Y(oc8051_sfr1_oc8051_uatr1_n62)
         );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u101 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_), .B(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_), .C(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_), .Y(oc8051_sfr1_oc8051_uatr1_n88) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u100 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_7_), .Y(oc8051_sfr1_oc8051_uatr1_n75) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u99 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_), .Y(oc8051_sfr1_oc8051_uatr1_n77) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u98 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_6_), .Y(oc8051_sfr1_oc8051_uatr1_n73) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u97 ( .A(
        oc8051_sfr1_oc8051_uatr1_n75), .B(oc8051_sfr1_oc8051_uatr1_n77), .C(
        oc8051_sfr1_oc8051_uatr1_n73), .Y(oc8051_sfr1_oc8051_uatr1_n90) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u96 ( .A(
        oc8051_sfr1_oc8051_uatr1_n90), .B(oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_), .C(oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_), .Y(oc8051_sfr1_oc8051_uatr1_n89)
         );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u95 ( .A(
        oc8051_sfr1_oc8051_uatr1_n200), .B(oc8051_sfr1_oc8051_uatr1_n199), .C(
        oc8051_sfr1_oc8051_uatr1_n88), .D(oc8051_sfr1_oc8051_uatr1_n89), .Y(
        oc8051_sfr1_oc8051_uatr1_n46) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u94 ( .A(
        oc8051_sfr1_oc8051_uatr1_n62), .B(oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_), .C(oc8051_sfr1_oc8051_uatr1_n46), .Y(oc8051_sfr1_oc8051_uatr1_n15) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u93 ( .A(
        oc8051_sfr1_oc8051_uatr1_n15), .Y(oc8051_sfr1_oc8051_uatr1_n49) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u92 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_), .Y(oc8051_sfr1_oc8051_uatr1_n6)
         );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u91 ( .A(
        oc8051_sfr1_oc8051_uatr1_n49), .B(oc8051_sfr1_oc8051_uatr1_n6), .C(
        oc8051_sfr1_oc8051_uatr1_trans), .Y(oc8051_sfr1_oc8051_uatr1_n84) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u90 ( .A(
        oc8051_sfr1_oc8051_uatr1_n87), .B(oc8051_sfr1_oc8051_uatr1_n79), .C(
        oc8051_sfr1_pres_ow), .Y(oc8051_sfr1_oc8051_uatr1_n47) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u89 ( .A(
        oc8051_sfr1_oc8051_uatr1_n47), .Y(oc8051_sfr1_oc8051_uatr1_n13) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u88 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .Y(oc8051_sfr1_oc8051_uatr1_n86) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u87 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_2_), .Y(oc8051_sfr1_oc8051_uatr1_n53) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u86 ( .AN(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .B(oc8051_sfr1_oc8051_uatr1_n86), .C(oc8051_sfr1_oc8051_uatr1_n201), .D(oc8051_sfr1_oc8051_uatr1_n53), .Y(
        oc8051_sfr1_oc8051_uatr1_n48) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u85 ( .A(
        oc8051_sfr1_oc8051_uatr1_n62), .B(oc8051_sfr1_oc8051_uatr1_n48), .Y(
        oc8051_sfr1_oc8051_uatr1_n12) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u84 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n46), .A1(oc8051_sfr1_oc8051_uatr1_n13), .B0(
        oc8051_sfr1_oc8051_uatr1_n12), .Y(oc8051_sfr1_oc8051_uatr1_n83) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u83 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n61), .A1(oc8051_sfr1_oc8051_uatr1_trans), 
        .B0(oc8051_sfr1_oc8051_uatr1_n83), .Y(oc8051_sfr1_oc8051_uatr1_n85) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u82 ( .A(txd_o), .B(
        oc8051_sfr1_oc8051_uatr1_n84), .S0(oc8051_sfr1_oc8051_uatr1_n85), .Y(
        oc8051_sfr1_oc8051_uatr1_n231) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u81 ( .A(
        oc8051_sfr1_oc8051_uatr1_n83), .B(oc8051_sfr1_oc8051_uatr1_n43), .Y(
        oc8051_sfr1_oc8051_uatr1_n5) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u80 ( .B0(
        oc8051_sfr1_oc8051_uatr1_n47), .B1(oc8051_sfr1_oc8051_uatr1_n62), 
        .A0N(oc8051_sfr1_oc8051_uatr1_n5), .Y(oc8051_sfr1_oc8051_uatr1_n1) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u79 ( .A(oc8051_sfr1_scon_6_), 
        .B(oc8051_sfr1_scon_3_), .S0(oc8051_sfr1_scon_7_), .Y(
        oc8051_sfr1_oc8051_uatr1_n82) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u78 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n199), .A1(oc8051_sfr1_oc8051_uatr1_n1), .B0(
        oc8051_sfr1_oc8051_uatr1_n43), .B1(oc8051_sfr1_oc8051_uatr1_n82), .C0(
        oc8051_sfr1_oc8051_uatr1_n200), .C1(oc8051_sfr1_oc8051_uatr1_n5), .Y(
        oc8051_sfr1_oc8051_uatr1_n232) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u77 ( .A(
        oc8051_sfr1_oc8051_uatr1_n79), .B(oc8051_sfr1_oc8051_uatr1_n61), .Y(
        oc8051_sfr1_oc8051_uatr1_n3) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u76 ( .A(
        oc8051_sfr1_oc8051_uatr1_n5), .Y(oc8051_sfr1_oc8051_uatr1_n81) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u75 ( .A0(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_), .A1(
        oc8051_sfr1_oc8051_uatr1_n81), .B0(wr_dat[7]), .B1(
        oc8051_sfr1_oc8051_uatr1_n61), .Y(oc8051_sfr1_oc8051_uatr1_n80) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u74 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n200), .A1(oc8051_sfr1_oc8051_uatr1_n1), .B0(
        oc8051_sfr1_oc8051_uatr1_n3), .C0(oc8051_sfr1_oc8051_uatr1_n80), .Y(
        oc8051_sfr1_oc8051_uatr1_n233) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u73 ( .A(
        oc8051_sfr1_oc8051_uatr1_n43), .B(oc8051_sfr1_oc8051_uatr1_n79), .Y(
        oc8051_sfr1_oc8051_uatr1_n65) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u72 ( .A(
        oc8051_sfr1_oc8051_uatr1_n3), .Y(oc8051_sfr1_oc8051_uatr1_n66) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u71 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n65), .A1(wr_dat[6]), .B0(wr_dat[7]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n78) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u70 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n77), .B0(
        oc8051_sfr1_oc8051_uatr1_n5), .B1(oc8051_sfr1_oc8051_uatr1_n75), .C0(
        oc8051_sfr1_oc8051_uatr1_n78), .Y(oc8051_sfr1_oc8051_uatr1_n234) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u69 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n65), .A1(wr_dat[5]), .B0(wr_dat[6]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n76) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u68 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n75), .B0(
        oc8051_sfr1_oc8051_uatr1_n5), .B1(oc8051_sfr1_oc8051_uatr1_n73), .C0(
        oc8051_sfr1_oc8051_uatr1_n76), .Y(oc8051_sfr1_oc8051_uatr1_n235) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u67 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_), .Y(oc8051_sfr1_oc8051_uatr1_n71) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u66 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n65), .A1(wr_dat[4]), .B0(wr_dat[5]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n74) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u65 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n73), .B0(
        oc8051_sfr1_oc8051_uatr1_n5), .B1(oc8051_sfr1_oc8051_uatr1_n71), .C0(
        oc8051_sfr1_oc8051_uatr1_n74), .Y(oc8051_sfr1_oc8051_uatr1_n236) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u64 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_), .Y(oc8051_sfr1_oc8051_uatr1_n69) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u63 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n65), .A1(wr_dat[3]), .B0(wr_dat[4]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n72) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u62 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n71), .B0(
        oc8051_sfr1_oc8051_uatr1_n5), .B1(oc8051_sfr1_oc8051_uatr1_n69), .C0(
        oc8051_sfr1_oc8051_uatr1_n72), .Y(oc8051_sfr1_oc8051_uatr1_n237) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u61 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_), .Y(oc8051_sfr1_oc8051_uatr1_n67) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u60 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_uatr1_n65), .B0(wr_dat[3]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n70) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u59 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n69), .B0(
        oc8051_sfr1_oc8051_uatr1_n5), .B1(oc8051_sfr1_oc8051_uatr1_n67), .C0(
        oc8051_sfr1_oc8051_uatr1_n70), .Y(oc8051_sfr1_oc8051_uatr1_n238) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u58 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_), .Y(oc8051_sfr1_oc8051_uatr1_n63) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u57 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_uatr1_n65), .B0(wr_dat[2]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n68) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u56 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n67), .B0(
        oc8051_sfr1_oc8051_uatr1_n5), .B1(oc8051_sfr1_oc8051_uatr1_n63), .C0(
        oc8051_sfr1_oc8051_uatr1_n68), .Y(oc8051_sfr1_oc8051_uatr1_n239) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u55 ( .A(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_), .Y(oc8051_sfr1_oc8051_uatr1_n2)
         );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u54 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n65), .A1(wr_dat[0]), .B0(wr_dat[1]), .B1(
        oc8051_sfr1_oc8051_uatr1_n66), .Y(oc8051_sfr1_oc8051_uatr1_n64) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u53 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n63), .B0(
        oc8051_sfr1_oc8051_uatr1_n2), .B1(oc8051_sfr1_oc8051_uatr1_n5), .C0(
        oc8051_sfr1_oc8051_uatr1_n64), .Y(oc8051_sfr1_oc8051_uatr1_n240) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u52 ( .A(
        oc8051_sfr1_oc8051_uatr1_n43), .B(oc8051_sfr1_oc8051_uatr1_n62), .Y(
        oc8051_sfr1_oc8051_uatr1_n56) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u51 ( .A(
        oc8051_sfr1_oc8051_uatr1_n56), .B(oc8051_sfr1_oc8051_uatr1_n43), .C(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .Y(oc8051_sfr1_oc8051_uatr1_n57) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u50 ( .A(
        oc8051_sfr1_oc8051_uatr1_n57), .Y(oc8051_sfr1_oc8051_uatr1_n52) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u49 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .B(oc8051_sfr1_oc8051_uatr1_n52), .Y(oc8051_sfr1_oc8051_uatr1_n59) );
  OA21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u48 ( .A0(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .A1(
        oc8051_sfr1_oc8051_uatr1_n61), .B0(oc8051_sfr1_oc8051_uatr1_n56), .Y(
        oc8051_sfr1_oc8051_uatr1_n58) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u47 ( .A0(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .A1(
        oc8051_sfr1_oc8051_uatr1_n61), .B0(oc8051_sfr1_oc8051_uatr1_n58), .Y(
        oc8051_sfr1_oc8051_uatr1_n54) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u46 ( .A(
        oc8051_sfr1_oc8051_uatr1_n54), .Y(oc8051_sfr1_oc8051_uatr1_n60) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u45 ( .A(
        oc8051_sfr1_oc8051_uatr1_n59), .B(oc8051_sfr1_oc8051_uatr1_n60), .S0(
        oc8051_sfr1_oc8051_uatr1_tr_count_2_), .Y(
        oc8051_sfr1_oc8051_uatr1_n242) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u44 ( .A(
        oc8051_sfr1_oc8051_uatr1_n57), .B(oc8051_sfr1_oc8051_uatr1_n58), .S0(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .Y(
        oc8051_sfr1_oc8051_uatr1_n243) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u43 ( .A(
        oc8051_sfr1_oc8051_uatr1_n56), .B(oc8051_sfr1_oc8051_uatr1_n43), .Y(
        oc8051_sfr1_oc8051_uatr1_n55) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u42 ( .A(
        oc8051_sfr1_oc8051_uatr1_n55), .B(oc8051_sfr1_oc8051_uatr1_n56), .S0(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_), .Y(
        oc8051_sfr1_oc8051_uatr1_n244) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u41 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n43), .A1(oc8051_sfr1_oc8051_uatr1_n53), .B0(
        oc8051_sfr1_oc8051_uatr1_n54), .Y(oc8051_sfr1_oc8051_uatr1_n50) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u40 ( .A(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_), .B(oc8051_sfr1_oc8051_uatr1_n52), .C(oc8051_sfr1_oc8051_uatr1_tr_count_2_), .Y(oc8051_sfr1_oc8051_uatr1_n51)
         );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u39 ( .A(
        oc8051_sfr1_oc8051_uatr1_n50), .B(oc8051_sfr1_oc8051_uatr1_n51), .S0(
        oc8051_sfr1_oc8051_uatr1_n201), .Y(oc8051_sfr1_oc8051_uatr1_n245) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u38 ( .A(
        oc8051_sfr1_oc8051_uatr1_trans), .Y(oc8051_sfr1_oc8051_uatr1_n44) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u37 ( .A(
        oc8051_sfr1_oc8051_uatr1_n48), .B(oc8051_sfr1_oc8051_uatr1_n49), .Y(
        oc8051_sfr1_oc8051_uatr1_n45) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u36 ( .A(
        oc8051_sfr1_oc8051_uatr1_n46), .B(oc8051_sfr1_oc8051_uatr1_n47), .Y(
        oc8051_sfr1_oc8051_uatr1_n14) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u35 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n44), .A1(oc8051_sfr1_oc8051_uatr1_n45), .A2(
        oc8051_sfr1_oc8051_uatr1_n14), .B0(oc8051_sfr1_oc8051_uatr1_n43), .Y(
        oc8051_sfr1_oc8051_uatr1_n246) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u34 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n43), .A1(oc8051_sfr1_oc8051_uatr1_n40), .B0(
        oc8051_sfr1_oc8051_uatr1_n199), .B1(oc8051_sfr1_oc8051_uatr1_n5), .Y(
        oc8051_sfr1_oc8051_uatr1_n247) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u33 ( .A(
        oc8051_sfr1_oc8051_uatr1_n41), .B(oc8051_sfr1_oc8051_uatr1_n42), .Y(
        oc8051_sfr1_oc8051_uatr1_n29) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u32 ( .A(
        oc8051_sfr1_oc8051_uatr1_n29), .B(oc8051_sfr1_oc8051_uatr1_n22), .Y(
        oc8051_sfr1_oc8051_uatr1_n37) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u31 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n37), .B(oc8051_sfr1_oc8051_uatr1_n40), .Y(
        oc8051_sfr1_oc8051_uatr1_n39) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u30 ( .A(
        oc8051_sfr1_oc8051_uatr1_n39), .B(wr_dat[7]), .S0(
        oc8051_sfr1_oc8051_uatr1_n20), .Y(oc8051_sfr1_oc8051_uatr1_n38) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u29 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n17), .A1(oc8051_sfr1_oc8051_uatr1_n37), .B0(
        oc8051_sfr1_oc8051_uatr1_n38), .Y(oc8051_sfr1_oc8051_uatr1_n248) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u28 ( .A(wr_addr[1]), .B(
        oc8051_sfr1_oc8051_uatr1_n27), .C(oc8051_sfr1_oc8051_uatr1_n29), .Y(
        oc8051_sfr1_oc8051_uatr1_n33) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u27 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n33), .B(oc8051_sfr1_oc8051_uatr1_n36), .Y(
        oc8051_sfr1_oc8051_uatr1_n35) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u26 ( .A(
        oc8051_sfr1_oc8051_uatr1_n35), .B(wr_dat[6]), .S0(
        oc8051_sfr1_oc8051_uatr1_n20), .Y(oc8051_sfr1_oc8051_uatr1_n34) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u25 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n17), .A1(oc8051_sfr1_oc8051_uatr1_n33), .B0(
        oc8051_sfr1_oc8051_uatr1_n34), .Y(oc8051_sfr1_oc8051_uatr1_n249) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u24 ( .A(
        oc8051_sfr1_oc8051_uatr1_n30), .B(oc8051_sfr1_scon_5_), .Y(
        oc8051_sfr1_oc8051_uatr1_n32) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u23 ( .A(
        oc8051_sfr1_oc8051_uatr1_n32), .B(wr_dat[5]), .S0(
        oc8051_sfr1_oc8051_uatr1_n20), .Y(oc8051_sfr1_oc8051_uatr1_n31) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u22 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n17), .A1(oc8051_sfr1_oc8051_uatr1_n30), .B0(
        oc8051_sfr1_oc8051_uatr1_n31), .Y(oc8051_sfr1_oc8051_uatr1_n250) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u21 ( .A(
        oc8051_sfr1_oc8051_uatr1_n27), .B(oc8051_sfr1_oc8051_uatr1_n28), .C(
        oc8051_sfr1_oc8051_uatr1_n29), .Y(oc8051_sfr1_oc8051_uatr1_n23) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u20 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n23), .B(oc8051_sfr1_oc8051_uatr1_n26), .Y(
        oc8051_sfr1_oc8051_uatr1_n25) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u19 ( .A(
        oc8051_sfr1_oc8051_uatr1_n25), .B(wr_dat[4]), .S0(
        oc8051_sfr1_oc8051_uatr1_n20), .Y(oc8051_sfr1_oc8051_uatr1_n24) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u18 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n17), .A1(oc8051_sfr1_oc8051_uatr1_n23), .B0(
        oc8051_sfr1_oc8051_uatr1_n24), .Y(oc8051_sfr1_oc8051_uatr1_n251) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u17 ( .AN(
        oc8051_sfr1_oc8051_uatr1_n21), .B(oc8051_sfr1_oc8051_uatr1_n22), .Y(
        oc8051_sfr1_oc8051_uatr1_n16) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u16 ( .A(
        oc8051_sfr1_oc8051_uatr1_n16), .B(oc8051_sfr1_scon_3_), .Y(
        oc8051_sfr1_oc8051_uatr1_n19) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u15 ( .A(
        oc8051_sfr1_oc8051_uatr1_n19), .B(wr_dat[3]), .S0(
        oc8051_sfr1_oc8051_uatr1_n20), .Y(oc8051_sfr1_oc8051_uatr1_n18) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u14 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n16), .A1(oc8051_sfr1_oc8051_uatr1_n17), .B0(
        oc8051_sfr1_oc8051_uatr1_n18), .Y(oc8051_sfr1_oc8051_uatr1_n252) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u13 ( .A(
        oc8051_sfr1_oc8051_uatr1_n14), .B(oc8051_sfr1_oc8051_uatr1_n15), .Y(
        oc8051_sfr1_oc8051_uatr1_n9) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u12 ( .A(
        oc8051_sfr1_oc8051_uatr1_n11), .B(oc8051_sfr1_oc8051_uatr1_n12), .C(
        oc8051_sfr1_oc8051_uatr1_n13), .Y(oc8051_sfr1_oc8051_uatr1_n10) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u11 ( .A(
        oc8051_sfr1_oc8051_uatr1_n9), .B(oc8051_sfr1_oc8051_uatr1_n198), .S0(
        oc8051_sfr1_oc8051_uatr1_n10), .Y(oc8051_sfr1_oc8051_uatr1_n253) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_uatr1_u10 ( .A(
        oc8051_sfr1_oc8051_uatr1_n8), .B(oc8051_sfr1_pcon[7]), .Y(
        oc8051_sfr1_oc8051_uatr1_n7) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u9 ( .A(
        oc8051_sfr1_oc8051_uatr1_smod_clk_tr), .B(oc8051_sfr1_oc8051_uatr1_n7), 
        .Y(oc8051_sfr1_oc8051_uatr1_n254) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u8 ( .A(wb_rst_i), .Y(
        oc8051_sfr1_oc8051_uatr1_n172) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u7 ( .A(
        oc8051_sfr1_oc8051_uatr1_n180), .Y(oc8051_sfr1_scon_1_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_uatr1_u6 ( .A(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_uatr1_n4) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u5 ( .A0(
        oc8051_sfr1_oc8051_uatr1_n1), .A1(oc8051_sfr1_oc8051_uatr1_n2), .B0(
        oc8051_sfr1_oc8051_uatr1_n3), .B1(oc8051_sfr1_oc8051_uatr1_n4), .C0(
        oc8051_sfr1_oc8051_uatr1_n5), .C1(oc8051_sfr1_oc8051_uatr1_n6), .Y(
        oc8051_sfr1_oc8051_uatr1_n170) );
  NAND3_X0P5M_A12TS oc8051_sfr1_oc8051_uatr1_u4 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_uatr1_n28), .C(oc8051_sfr1_oc8051_uatr1_n29), .Y(
        oc8051_sfr1_oc8051_uatr1_n30) );
  AND4_X0P7M_A12TS oc8051_sfr1_oc8051_uatr1_u3 ( .A(
        oc8051_sfr1_oc8051_uatr1_n22), .B(oc8051_sfr1_oc8051_uatr1_n132), .C(
        wr_addr[2]), .D(oc8051_sfr1_oc8051_uatr1_n162), .Y(
        oc8051_sfr1_oc8051_uatr1_n161) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n224), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n180) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tx_done_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n253), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n198) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_9_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n232), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n200) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_10_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n247), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n199) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n245), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n201) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rx_done_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n225), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_uatr1_n172), .Q(oc8051_sfr1_oc8051_uatr1_rx_done)
         );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n215), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n203) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n214), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n202) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n226), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n204) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_uatr1_t1_ow_buf_reg ( .D(
        oc8051_sfr1_tf1), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_uatr1_n205) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n248), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n251), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n243), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_tr_count_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n219), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n197), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n244), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_tr_count_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n218), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n249), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_trans_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n246), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_trans) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n223), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_receive_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n221), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_receive) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n252), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n250), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_tr_count_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n242), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_tr_count_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n216), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_re_count_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n217), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_re_count_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_scon_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n222), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_scon_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_smod_clk_tr_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n254), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_smod_clk_tr) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_smod_clk_re_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n230), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_smod_clk_re) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rx_sam_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n228), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_rx_sam_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_11_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n227), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_11_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n239), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n237), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_8_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n233), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_8_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rx_sam_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n229), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_rx_sam_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n240), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_shift_re_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n269), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_shift_re) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n170), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n238), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n236), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n213), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n212), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n211), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n210), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n209), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_8_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n207), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_8_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_9_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n208), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_9_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_reg_10_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n206), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_rxd_tmp_10_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n181), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n182), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n183), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n184), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n185), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n186), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n187), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_rxd_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n188), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_sbuf[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_0_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n190), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_1_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n191), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_2_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n192), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_3_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n193), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_4_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n194), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_5_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n195), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_pcon_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n196), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_pcon[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_6_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n235), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_sbuf_txd_reg_7_ ( .D(
        oc8051_sfr1_oc8051_uatr1_n234), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_sbuf_txd_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_shift_tr_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n174), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_uatr1_shift_tr) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_rxd_r_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n220), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_uatr1_n172), .Q(oc8051_sfr1_oc8051_uatr1_rxd_r) );
  DFFSQ_X1M_A12TS oc8051_sfr1_oc8051_uatr1_txd_reg ( .D(
        oc8051_sfr1_oc8051_uatr1_n231), .CK(wb_clk_i), .SN(
        oc8051_sfr1_oc8051_uatr1_n172), .Q(txd_o) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u244 ( .A(oc8051_sfr1_oc8051_int1_n8), .Y(int_src[5]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u243 ( .A(oc8051_sfr1_oc8051_int1_n7), .Y(int_src[4]) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u242 ( .A(int_src[5]), .B(
        int_src[4]), .Y(oc8051_sfr1_oc8051_int1_n209) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u241 ( .A(
        oc8051_sfr1_oc8051_int1_n4), .B(oc8051_sfr1_oc8051_int1_n5), .C(
        oc8051_sfr1_oc8051_int1_n209), .D(oc8051_sfr1_oc8051_int1_n6), .Y(intr) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u240 ( .A(reti), .B(
        oc8051_sfr1_oc8051_int1_int_proc), .Y(oc8051_sfr1_oc8051_int1_n154) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u239 ( .A(oc8051_sfr1_ie_0_), .B(
        oc8051_sfr1_ip_0_), .C(oc8051_sfr1_tcon_1_), .Y(
        oc8051_sfr1_oc8051_int1_n183) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u238 ( .A(oc8051_sfr1_tcon_5_), 
        .B(oc8051_sfr1_ie_1_), .Y(oc8051_sfr1_oc8051_int1_n186) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u237 ( .A(
        oc8051_sfr1_oc8051_int1_n186), .Y(oc8051_sfr1_oc8051_int1_n181) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u236 ( .A(
        oc8051_sfr1_oc8051_int1_n181), .B(oc8051_sfr1_ip_1_), .Y(
        oc8051_sfr1_oc8051_int1_n184) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u235 ( .A(oc8051_sfr1_ie_2_), .B(
        oc8051_sfr1_ip_2_), .C(oc8051_sfr1_tcon_3_), .Y(
        oc8051_sfr1_oc8051_int1_n208) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u234 ( .A(
        oc8051_sfr1_oc8051_int1_n183), .B(oc8051_sfr1_oc8051_int1_n184), .C(
        oc8051_sfr1_oc8051_int1_n208), .Y(oc8051_sfr1_oc8051_int1_n200) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u233 ( .A(oc8051_sfr1_tcon_7_), 
        .B(oc8051_sfr1_ie_3_), .Y(oc8051_sfr1_oc8051_int1_n195) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u232 ( .A(oc8051_sfr1_ip_3_), .Y(
        oc8051_sfr1_oc8051_int1_n27) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u231 ( .A(
        oc8051_sfr1_oc8051_int1_n195), .B(oc8051_sfr1_oc8051_int1_n27), .Y(
        oc8051_sfr1_oc8051_int1_n201) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u230 ( .AN(
        oc8051_sfr1_oc8051_int1_n200), .B(oc8051_sfr1_oc8051_int1_n201), .Y(
        oc8051_sfr1_oc8051_int1_n194) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u229 ( .A(oc8051_sfr1_tc2_int), .Y(
        oc8051_sfr1_oc8051_int1_n197) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u228 ( .A(oc8051_sfr1_ie_5_), .Y(
        oc8051_sfr1_oc8051_int1_n66) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u227 ( .A(oc8051_sfr1_ie_4_), .B(
        oc8051_sfr1_ip_4_), .C(oc8051_sfr1_uart_int), .Y(
        oc8051_sfr1_oc8051_int1_n193) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u226 ( .A0(
        oc8051_sfr1_oc8051_int1_n197), .A1(oc8051_sfr1_oc8051_int1_n9), .A2(
        oc8051_sfr1_oc8051_int1_n66), .B0(oc8051_sfr1_oc8051_int1_n193), .Y(
        oc8051_sfr1_oc8051_int1_n205) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u225 ( .A(oc8051_sfr1_ie_7_), .Y(
        oc8051_sfr1_oc8051_int1_n55) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u224 ( .A(
        oc8051_sfr1_oc8051_int1_n52), .B(oc8051_sfr1_oc8051_int1_n53), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n207)
         );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u223 ( .A0(
        oc8051_sfr1_oc8051_int1_n55), .A1(oc8051_sfr1_oc8051_int1_n207), .B0(
        oc8051_sfr1_oc8051_int1_int_proc), .Y(oc8051_sfr1_oc8051_int1_n206) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u222 ( .A1N(
        oc8051_sfr1_oc8051_int1_n194), .A0(oc8051_sfr1_oc8051_int1_n205), .B0(
        oc8051_sfr1_oc8051_int1_n206), .Y(oc8051_sfr1_oc8051_int1_n202) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u221 ( .A(
        oc8051_sfr1_oc8051_int1_n154), .B(oc8051_sfr1_oc8051_int1_n202), .Y(
        oc8051_sfr1_oc8051_int1_n151) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u220 ( .A(
        oc8051_sfr1_oc8051_int1_n151), .Y(oc8051_sfr1_oc8051_int1_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u219 ( .A(
        oc8051_sfr1_oc8051_int1_n195), .Y(oc8051_sfr1_oc8051_int1_n204) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u218 ( .A(oc8051_sfr1_ie_2_), .Y(
        oc8051_sfr1_oc8051_int1_n75) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u217 ( .A(oc8051_sfr1_tcon_3_), .Y(
        oc8051_sfr1_oc8051_int1_n143) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u216 ( .A(oc8051_sfr1_tcon_1_), 
        .B(oc8051_sfr1_ie_0_), .Y(oc8051_sfr1_oc8051_int1_n188) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u215 ( .A0(
        oc8051_sfr1_oc8051_int1_n75), .A1(oc8051_sfr1_oc8051_int1_n143), .B0(
        oc8051_sfr1_oc8051_int1_n186), .C0(oc8051_sfr1_oc8051_int1_n188), .Y(
        oc8051_sfr1_oc8051_int1_n191) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u214 ( .A0(oc8051_sfr1_ie_4_), 
        .A1(oc8051_sfr1_uart_int), .B0(oc8051_sfr1_oc8051_int1_n204), .C0(
        oc8051_sfr1_oc8051_int1_n191), .Y(oc8051_sfr1_oc8051_int1_n198) );
  OA21A1OI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u213 ( .A0(
        oc8051_sfr1_oc8051_int1_n66), .A1(oc8051_sfr1_oc8051_int1_n197), .B0(
        oc8051_sfr1_oc8051_int1_n198), .C0(oc8051_sfr1_oc8051_int1_int_proc), 
        .Y(oc8051_sfr1_oc8051_int1_n203) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u212 ( .A(
        oc8051_sfr1_oc8051_int1_n159), .B(oc8051_sfr1_ie_7_), .C(
        oc8051_sfr1_oc8051_int1_n203), .Y(oc8051_sfr1_oc8051_int1_n179) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u211 ( .A(
        oc8051_sfr1_oc8051_int1_n154), .Y(oc8051_sfr1_oc8051_int1_n155) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u210 ( .A(
        oc8051_sfr1_oc8051_int1_n202), .B(oc8051_sfr1_oc8051_int1_n155), .Y(
        oc8051_sfr1_oc8051_int1_n162) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u209 ( .A(
        oc8051_sfr1_oc8051_int1_n162), .B(oc8051_sfr1_oc8051_int1_n200), .C(
        oc8051_sfr1_oc8051_int1_n201), .Y(oc8051_sfr1_oc8051_int1_n199) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u208 ( .A0(
        oc8051_sfr1_oc8051_int1_n179), .A1(oc8051_sfr1_oc8051_int1_n195), .A2(
        oc8051_sfr1_oc8051_int1_n191), .B0(oc8051_sfr1_oc8051_int1_n199), .Y(
        oc8051_sfr1_oc8051_int1_n167) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u207 ( .A(
        oc8051_sfr1_oc8051_int1_n167), .Y(oc8051_sfr1_oc8051_int1_n170) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u206 ( .A(
        oc8051_sfr1_oc8051_int1_n179), .Y(oc8051_sfr1_oc8051_int1_n160) );
  AOI32_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u205 ( .A0(
        oc8051_sfr1_oc8051_int1_n194), .A1(oc8051_sfr1_oc8051_int1_n193), .A2(
        oc8051_sfr1_oc8051_int1_n162), .B0(oc8051_sfr1_oc8051_int1_n160), .B1(
        oc8051_sfr1_oc8051_int1_n198), .Y(oc8051_sfr1_oc8051_int1_n196) );
  OR3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u204 ( .A(
        oc8051_sfr1_oc8051_int1_n196), .B(oc8051_sfr1_oc8051_int1_n66), .C(
        oc8051_sfr1_oc8051_int1_n197), .Y(oc8051_sfr1_oc8051_int1_n165) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u203 ( .A(oc8051_sfr1_ie_4_), .B(
        oc8051_sfr1_oc8051_int1_n195), .C(oc8051_sfr1_uart_int), .Y(
        oc8051_sfr1_oc8051_int1_n190) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u202 ( .AN(
        oc8051_sfr1_oc8051_int1_n193), .B(oc8051_sfr1_oc8051_int1_n162), .C(
        oc8051_sfr1_oc8051_int1_n194), .Y(oc8051_sfr1_oc8051_int1_n192) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u201 ( .A0(
        oc8051_sfr1_oc8051_int1_n190), .A1(oc8051_sfr1_oc8051_int1_n191), .A2(
        oc8051_sfr1_oc8051_int1_n179), .B0(oc8051_sfr1_oc8051_int1_n192), .Y(
        oc8051_sfr1_oc8051_int1_n189) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u200 ( .A(
        oc8051_sfr1_oc8051_int1_n189), .Y(oc8051_sfr1_oc8051_int1_n171) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u199 ( .A(
        oc8051_sfr1_oc8051_int1_n170), .B(oc8051_sfr1_oc8051_int1_n165), .C(
        oc8051_sfr1_oc8051_int1_n171), .Y(oc8051_sfr1_oc8051_int1_n117) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u198 ( .A(
        oc8051_sfr1_oc8051_int1_int_dept_1_), .B(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n152)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u197 ( .A(
        oc8051_sfr1_oc8051_int1_n188), .Y(oc8051_sfr1_oc8051_int1_n180) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u196 ( .AN(
        oc8051_sfr1_oc8051_int1_n184), .B(oc8051_sfr1_oc8051_int1_n162), .C(
        oc8051_sfr1_oc8051_int1_n183), .Y(oc8051_sfr1_oc8051_int1_n187) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u195 ( .A0(
        oc8051_sfr1_oc8051_int1_n179), .A1(oc8051_sfr1_oc8051_int1_n180), .A2(
        oc8051_sfr1_oc8051_int1_n186), .B0(oc8051_sfr1_oc8051_int1_n187), .Y(
        oc8051_sfr1_oc8051_int1_n168) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u194 ( .A(
        oc8051_sfr1_oc8051_int1_n168), .Y(oc8051_sfr1_oc8051_int1_n177) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u193 ( .A(
        oc8051_sfr1_oc8051_int1_n183), .Y(oc8051_sfr1_oc8051_int1_n185) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u192 ( .A0(
        oc8051_sfr1_oc8051_int1_n160), .A1(oc8051_sfr1_oc8051_int1_n180), .B0(
        oc8051_sfr1_oc8051_int1_n162), .B1(oc8051_sfr1_oc8051_int1_n185), .Y(
        oc8051_sfr1_oc8051_int1_n175) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u191 ( .A(
        oc8051_sfr1_oc8051_int1_n162), .B(oc8051_sfr1_ip_2_), .C(
        oc8051_sfr1_oc8051_int1_n183), .D(oc8051_sfr1_oc8051_int1_n184), .Y(
        oc8051_sfr1_oc8051_int1_n182) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u190 ( .A0(
        oc8051_sfr1_oc8051_int1_n179), .A1(oc8051_sfr1_oc8051_int1_n180), .A2(
        oc8051_sfr1_oc8051_int1_n181), .B0(oc8051_sfr1_oc8051_int1_n182), .Y(
        oc8051_sfr1_oc8051_int1_n178) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u189 ( .A(oc8051_sfr1_ie_2_), .B(
        oc8051_sfr1_oc8051_int1_n178), .C(oc8051_sfr1_tcon_3_), .Y(
        oc8051_sfr1_oc8051_int1_n169) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u188 ( .A(
        oc8051_sfr1_oc8051_int1_n117), .B(oc8051_sfr1_oc8051_int1_n177), .C(
        oc8051_sfr1_oc8051_int1_n175), .D(oc8051_sfr1_oc8051_int1_n169), .Y(
        oc8051_sfr1_oc8051_int1_n172) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u187 ( .A(
        oc8051_sfr1_oc8051_int1_n152), .B(oc8051_sfr1_oc8051_int1_n172), .Y(
        oc8051_sfr1_oc8051_int1_n174) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u186 ( .A(
        oc8051_sfr1_oc8051_int1_n47), .B(oc8051_sfr1_oc8051_int1_n117), .S0(
        oc8051_sfr1_oc8051_int1_n174), .Y(oc8051_sfr1_oc8051_int1_n235) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u185 ( .A(
        oc8051_sfr1_oc8051_int1_n169), .B(oc8051_sfr1_oc8051_int1_n165), .C(
        oc8051_sfr1_oc8051_int1_n177), .Y(oc8051_sfr1_oc8051_int1_n176) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u184 ( .A(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n157)
         );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u183 ( .A(
        oc8051_sfr1_oc8051_int1_n157), .B(oc8051_sfr1_oc8051_int1_int_dept_1_), 
        .Y(oc8051_sfr1_oc8051_int1_n153) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u182 ( .A(
        oc8051_sfr1_oc8051_int1_n153), .B(oc8051_sfr1_oc8051_int1_n172), .Y(
        oc8051_sfr1_oc8051_int1_n118) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u181 ( .A(
        oc8051_sfr1_oc8051_int1_n45), .B(oc8051_sfr1_oc8051_int1_n176), .S0(
        oc8051_sfr1_oc8051_int1_n118), .Y(oc8051_sfr1_oc8051_int1_n236) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u180 ( .A(
        oc8051_sfr1_oc8051_int1_n48), .B(oc8051_sfr1_oc8051_int1_n176), .S0(
        oc8051_sfr1_oc8051_int1_n174), .Y(oc8051_sfr1_oc8051_int1_n237) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u179 ( .A(
        oc8051_sfr1_oc8051_int1_n171), .B(oc8051_sfr1_oc8051_int1_n169), .C(
        oc8051_sfr1_oc8051_int1_n175), .Y(oc8051_sfr1_oc8051_int1_n173) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u178 ( .A(
        oc8051_sfr1_oc8051_int1_n46), .B(oc8051_sfr1_oc8051_int1_n173), .S0(
        oc8051_sfr1_oc8051_int1_n118), .Y(oc8051_sfr1_oc8051_int1_n238) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u177 ( .A(
        oc8051_sfr1_oc8051_int1_n49), .B(oc8051_sfr1_oc8051_int1_n173), .S0(
        oc8051_sfr1_oc8051_int1_n174), .Y(oc8051_sfr1_oc8051_int1_n239) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u176 ( .AN(
        oc8051_sfr1_oc8051_int1_n172), .B(oc8051_sfr1_oc8051_int1_n151), .Y(
        oc8051_sfr1_oc8051_int1_n164) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u175 ( .A0(
        oc8051_sfr1_oc8051_int1_n8), .A1(oc8051_sfr1_oc8051_int1_n164), .B0(
        oc8051_sfr1_oc8051_int1_n165), .C0(oc8051_sfr1_oc8051_int1_n171), .Y(
        oc8051_sfr1_oc8051_int1_n240) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u174 ( .A0(
        oc8051_sfr1_oc8051_int1_n7), .A1(oc8051_sfr1_oc8051_int1_n164), .B0(
        oc8051_sfr1_oc8051_int1_n169), .C0(oc8051_sfr1_oc8051_int1_n170), .Y(
        oc8051_sfr1_oc8051_int1_n241) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u173 ( .A(
        oc8051_sfr1_oc8051_int1_n167), .B(oc8051_sfr1_oc8051_int1_n168), .Y(
        oc8051_sfr1_oc8051_int1_n166) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u172 ( .A0(
        oc8051_sfr1_oc8051_int1_n6), .A1(oc8051_sfr1_oc8051_int1_n164), .B0(
        oc8051_sfr1_oc8051_int1_n165), .C0(oc8051_sfr1_oc8051_int1_n166), .Y(
        oc8051_sfr1_oc8051_int1_n242) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u171 ( .A(
        oc8051_sfr1_oc8051_int1_n160), .B(oc8051_sfr1_oc8051_int1_n162), .Y(
        oc8051_sfr1_oc8051_int1_n156) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u170 ( .A0(
        oc8051_sfr1_oc8051_int1_n5), .A1(oc8051_sfr1_oc8051_int1_n164), .B0(
        oc8051_sfr1_oc8051_int1_n156), .Y(oc8051_sfr1_oc8051_int1_n243) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u169 ( .A0(
        oc8051_sfr1_oc8051_int1_n4), .A1(oc8051_sfr1_oc8051_int1_n164), .B0(
        oc8051_sfr1_oc8051_int1_n156), .Y(oc8051_sfr1_oc8051_int1_n244) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u168 ( .A(
        oc8051_sfr1_oc8051_int1_n153), .B(oc8051_sfr1_oc8051_int1_n162), .Y(
        oc8051_sfr1_oc8051_int1_n163) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u167 ( .A0(
        oc8051_sfr1_oc8051_int1_n153), .A1(oc8051_sfr1_oc8051_int1_n160), .B0(
        oc8051_sfr1_oc8051_int1_n52), .C0(oc8051_sfr1_oc8051_int1_n163), .Y(
        oc8051_sfr1_oc8051_int1_n245) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u166 ( .A(
        oc8051_sfr1_oc8051_int1_n152), .B(oc8051_sfr1_oc8051_int1_n162), .Y(
        oc8051_sfr1_oc8051_int1_n161) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u165 ( .A0(
        oc8051_sfr1_oc8051_int1_n152), .A1(oc8051_sfr1_oc8051_int1_n160), .B0(
        oc8051_sfr1_oc8051_int1_n53), .C0(oc8051_sfr1_oc8051_int1_n161), .Y(
        oc8051_sfr1_oc8051_int1_n246) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u164 ( .A(
        oc8051_sfr1_oc8051_int1_n159), .B(oc8051_sfr1_oc8051_int1_n157), .Y(
        oc8051_sfr1_oc8051_int1_n158) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u163 ( .A(
        oc8051_sfr1_oc8051_int1_n156), .B(oc8051_sfr1_oc8051_int1_n154), .Y(
        oc8051_sfr1_oc8051_int1_n147) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u162 ( .A(
        oc8051_sfr1_oc8051_int1_n157), .B(oc8051_sfr1_oc8051_int1_n158), .S0(
        oc8051_sfr1_oc8051_int1_n147), .Y(oc8051_sfr1_oc8051_int1_n247) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u161 ( .A(
        oc8051_sfr1_oc8051_int1_int_proc), .Y(oc8051_sfr1_oc8051_int1_n107) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u160 ( .A0(
        oc8051_sfr1_oc8051_int1_n155), .A1(oc8051_sfr1_oc8051_int1_n153), .B0(
        oc8051_sfr1_oc8051_int1_n107), .C0(oc8051_sfr1_oc8051_int1_n156), .Y(
        oc8051_sfr1_oc8051_int1_n248) );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u159 ( .A(
        oc8051_sfr1_oc8051_int1_n154), .B(oc8051_sfr1_oc8051_int1_int_dept_0_), 
        .Y(oc8051_sfr1_oc8051_int1_n149) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u158 ( .A(
        oc8051_sfr1_oc8051_int1_n152), .B(oc8051_sfr1_oc8051_int1_n153), .S0(
        oc8051_sfr1_oc8051_int1_n154), .Y(oc8051_sfr1_oc8051_int1_n150) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u157 ( .A0(
        oc8051_sfr1_oc8051_int1_n149), .A1(oc8051_sfr1_oc8051_int1_int_dept_1_), .B0(oc8051_sfr1_oc8051_int1_n150), .C0(oc8051_sfr1_oc8051_int1_n151), .Y(
        oc8051_sfr1_oc8051_int1_n148) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u156 ( .A1N(
        oc8051_sfr1_oc8051_int1_int_dept_1_), .A0(oc8051_sfr1_oc8051_int1_n147), .B0(oc8051_sfr1_oc8051_int1_n148), .Y(oc8051_sfr1_oc8051_int1_n249) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u155 ( .A(
        oc8051_sfr1_oc8051_int1_n46), .B(oc8051_sfr1_oc8051_int1_n49), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n146)
         );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u154 ( .A(
        oc8051_sfr1_oc8051_int1_n146), .B(oc8051_sfr1_oc8051_int1_int_proc), 
        .Y(oc8051_sfr1_oc8051_int1_n110) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u153 ( .A(
        oc8051_sfr1_oc8051_int1_n43), .B(oc8051_sfr1_oc8051_int1_n47), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n111)
         );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u152 ( .A(int_ack), .Y(
        oc8051_sfr1_oc8051_int1_n108) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u151 ( .A(
        oc8051_sfr1_oc8051_int1_n111), .B(oc8051_sfr1_oc8051_int1_n108), .Y(
        oc8051_sfr1_oc8051_int1_n133) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u150 ( .A(
        oc8051_sfr1_oc8051_int1_n133), .Y(oc8051_sfr1_oc8051_int1_n125) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u149 ( .A(
        oc8051_sfr1_oc8051_int1_n45), .B(oc8051_sfr1_oc8051_int1_n48), .S0(
        oc8051_sfr1_oc8051_int1_int_dept_0_), .Y(oc8051_sfr1_oc8051_int1_n145)
         );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u148 ( .A(
        oc8051_sfr1_oc8051_int1_n145), .B(oc8051_sfr1_oc8051_int1_int_proc), 
        .Y(oc8051_sfr1_oc8051_int1_n109) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u147 ( .A(wr_addr[4]), .B(
        wr_addr[6]), .C(wr_addr[5]), .Y(oc8051_sfr1_oc8051_int1_n144) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u146 ( .A(wr_addr[7]), .B(n_5_net_), 
        .C(wr_addr[3]), .D(oc8051_sfr1_oc8051_int1_n144), .Y(
        oc8051_sfr1_oc8051_int1_n141) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u145 ( .A(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_int1_n44) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u144 ( .AN(
        oc8051_sfr1_oc8051_int1_n141), .B(oc8051_sfr1_oc8051_int1_n44), .Y(
        oc8051_sfr1_oc8051_int1_n113) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u143 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_int1_n115) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u142 ( .A(
        oc8051_sfr1_oc8051_int1_n115), .B(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_int1_n29) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u141 ( .A(
        oc8051_sfr1_oc8051_int1_n113), .B(oc8051_sfr1_oc8051_int1_n29), .Y(
        oc8051_sfr1_oc8051_int1_n94) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u140 ( .AN(
        oc8051_sfr1_oc8051_int1_n94), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n137) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u139 ( .A0(
        oc8051_sfr1_oc8051_int1_n110), .A1(oc8051_sfr1_oc8051_int1_n125), .A2(
        oc8051_sfr1_oc8051_int1_n109), .B0(oc8051_sfr1_oc8051_int1_n137), .Y(
        oc8051_sfr1_oc8051_int1_n142) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u138 ( .A(oc8051_sfr1_tcon_2_), .Y(
        oc8051_sfr1_oc8051_int1_n139) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u137 ( .A(
        oc8051_sfr1_oc8051_int1_n142), .B(oc8051_sfr1_oc8051_int1_n139), .C(
        oc8051_sfr1_oc8051_int1_n143), .Y(oc8051_sfr1_oc8051_int1_n140) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u136 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n38) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u135 ( .A(wr_addr[2]), .B(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_int1_n36) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u134 ( .A(
        oc8051_sfr1_oc8051_int1_n38), .B(oc8051_sfr1_oc8051_int1_n44), .C(
        oc8051_sfr1_oc8051_int1_n36), .Y(oc8051_sfr1_oc8051_int1_n84) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u133 ( .A(
        oc8051_sfr1_oc8051_int1_n141), .B(oc8051_sfr1_oc8051_int1_n84), .Y(
        oc8051_sfr1_oc8051_int1_n116) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u132 ( .A(
        oc8051_sfr1_oc8051_int1_n116), .Y(oc8051_sfr1_oc8051_int1_n90) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u131 ( .A(
        oc8051_sfr1_oc8051_int1_n140), .B(wr_dat[3]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n134) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u130 ( .A(
        oc8051_sfr1_oc8051_int1_ie1_buff), .B(oc8051_sfr1_oc8051_int1_n139), 
        .Y(oc8051_sfr1_oc8051_int1_n138) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u129 ( .A(
        oc8051_sfr1_oc8051_int1_n138), .B(int1_i), .C(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n136) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u128 ( .A(descy), .B(
        oc8051_sfr1_oc8051_int1_n136), .S0(oc8051_sfr1_oc8051_int1_n137), .Y(
        oc8051_sfr1_oc8051_int1_n135) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u127 ( .A(
        oc8051_sfr1_oc8051_int1_n134), .B(oc8051_sfr1_oc8051_int1_n135), .Y(
        oc8051_sfr1_oc8051_int1_n250) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u126 ( .A(
        oc8051_sfr1_oc8051_int1_n110), .Y(oc8051_sfr1_oc8051_int1_n124) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u125 ( .A(
        oc8051_sfr1_oc8051_int1_n113), .B(oc8051_sfr1_oc8051_int1_n36), .Y(
        oc8051_sfr1_oc8051_int1_n97) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u124 ( .A(
        oc8051_sfr1_oc8051_int1_n97), .B(oc8051_sfr1_oc8051_int1_n38), .Y(
        oc8051_sfr1_oc8051_int1_n129) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u123 ( .A0(
        oc8051_sfr1_oc8051_int1_n124), .A1(oc8051_sfr1_oc8051_int1_n109), .A2(
        oc8051_sfr1_oc8051_int1_n133), .B0(oc8051_sfr1_oc8051_int1_n129), .Y(
        oc8051_sfr1_oc8051_int1_n132) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u122 ( .A(
        oc8051_sfr1_oc8051_int1_n132), .B(oc8051_sfr1_tcon_0_), .C(
        oc8051_sfr1_tcon_1_), .Y(oc8051_sfr1_oc8051_int1_n131) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u121 ( .A(
        oc8051_sfr1_oc8051_int1_n131), .B(wr_dat[1]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n126) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u120 ( .AN(oc8051_sfr1_tcon_0_), 
        .B(oc8051_sfr1_oc8051_int1_ie0_buff), .Y(oc8051_sfr1_oc8051_int1_n130)
         );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u119 ( .A(
        oc8051_sfr1_oc8051_int1_n130), .B(int0_i), .C(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n128) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u118 ( .A(
        oc8051_sfr1_oc8051_int1_n128), .B(descy), .S0(
        oc8051_sfr1_oc8051_int1_n129), .Y(oc8051_sfr1_oc8051_int1_n127) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u117 ( .A(
        oc8051_sfr1_oc8051_int1_n126), .B(oc8051_sfr1_oc8051_int1_n127), .Y(
        oc8051_sfr1_oc8051_int1_n251) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u116 ( .A0(
        oc8051_sfr1_oc8051_int1_n109), .A1(oc8051_sfr1_oc8051_int1_n124), .A2(
        oc8051_sfr1_oc8051_int1_n125), .B0(oc8051_sfr1_tcon_5_), .Y(
        oc8051_sfr1_oc8051_int1_n123) );
  OAI2XB1_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u115 ( .A1N(oc8051_sfr1_tf0), 
        .A0(oc8051_sfr1_oc8051_int1_tf0_buff), .B0(
        oc8051_sfr1_oc8051_int1_n123), .Y(oc8051_sfr1_oc8051_int1_n121) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u114 ( .A(wr_addr[2]), .Y(
        oc8051_sfr1_oc8051_int1_n114) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u113 ( .A(
        oc8051_sfr1_oc8051_int1_n114), .B(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_int1_n21) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u112 ( .A(
        oc8051_sfr1_oc8051_int1_n113), .B(oc8051_sfr1_oc8051_int1_n21), .Y(
        oc8051_sfr1_oc8051_int1_n91) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u111 ( .A(
        oc8051_sfr1_oc8051_int1_n38), .B(oc8051_sfr1_oc8051_int1_n91), .Y(
        oc8051_sfr1_oc8051_int1_n122) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u110 ( .A(
        oc8051_sfr1_oc8051_int1_n121), .B(descy), .S0(
        oc8051_sfr1_oc8051_int1_n122), .Y(oc8051_sfr1_oc8051_int1_n119) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u109 ( .A(
        oc8051_sfr1_oc8051_int1_n119), .B(oc8051_sfr1_oc8051_int1_n120), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n252) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u108 ( .A(
        oc8051_sfr1_oc8051_int1_n43), .B(oc8051_sfr1_oc8051_int1_n117), .S0(
        oc8051_sfr1_oc8051_int1_n118), .Y(oc8051_sfr1_oc8051_int1_n253) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u107 ( .AN(
        oc8051_sfr1_oc8051_int1_tf1_buff), .B(oc8051_sfr1_oc8051_int1_n116), 
        .C(oc8051_sfr1_tf1), .Y(oc8051_sfr1_oc8051_int1_n112) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u106 ( .A(descy), .Y(
        oc8051_sfr1_oc8051_int1_n86) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u105 ( .A(
        oc8051_sfr1_oc8051_int1_n114), .B(oc8051_sfr1_oc8051_int1_n115), .Y(
        oc8051_sfr1_oc8051_int1_n11) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u104 ( .A(
        oc8051_sfr1_oc8051_int1_n113), .B(oc8051_sfr1_oc8051_int1_n11), .Y(
        oc8051_sfr1_oc8051_int1_n87) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u103 ( .A(
        oc8051_sfr1_oc8051_int1_n87), .B(oc8051_sfr1_oc8051_int1_n38), .Y(
        oc8051_sfr1_oc8051_int1_n104) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u102 ( .A(
        oc8051_sfr1_oc8051_int1_n112), .B(oc8051_sfr1_oc8051_int1_n86), .S0(
        oc8051_sfr1_oc8051_int1_n104), .Y(oc8051_sfr1_oc8051_int1_n100) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u101 ( .A(oc8051_sfr1_tcon_7_), .Y(
        oc8051_sfr1_oc8051_int1_n103) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u100 ( .A(
        oc8051_sfr1_oc8051_int1_n109), .B(oc8051_sfr1_oc8051_int1_n110), .C(
        oc8051_sfr1_oc8051_int1_n111), .Y(oc8051_sfr1_oc8051_int1_n106) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u99 ( .A(
        oc8051_sfr1_oc8051_int1_n106), .B(oc8051_sfr1_oc8051_int1_n107), .C(
        oc8051_sfr1_oc8051_int1_n108), .Y(oc8051_sfr1_oc8051_int1_n105) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u98 ( .A(
        oc8051_sfr1_oc8051_int1_n103), .B(oc8051_sfr1_oc8051_int1_n104), .C(
        oc8051_sfr1_oc8051_int1_n105), .Y(oc8051_sfr1_oc8051_int1_n102) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u97 ( .A(
        oc8051_sfr1_oc8051_int1_n102), .B(wr_dat[7]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n101) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u96 ( .AN(
        oc8051_sfr1_oc8051_int1_n100), .B(oc8051_sfr1_oc8051_int1_n101), .Y(
        oc8051_sfr1_oc8051_int1_n254) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u95 ( .A(
        oc8051_sfr1_oc8051_int1_n97), .B(oc8051_sfr1_tcon_0_), .Y(
        oc8051_sfr1_oc8051_int1_n99) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u94 ( .A(
        oc8051_sfr1_oc8051_int1_n99), .B(wr_dat[0]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n98) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u93 ( .A0(
        oc8051_sfr1_oc8051_int1_n86), .A1(oc8051_sfr1_oc8051_int1_n97), .B0(
        oc8051_sfr1_oc8051_int1_n98), .Y(oc8051_sfr1_oc8051_int1_n255) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u92 ( .A(
        oc8051_sfr1_oc8051_int1_n94), .B(oc8051_sfr1_tcon_2_), .Y(
        oc8051_sfr1_oc8051_int1_n96) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u91 ( .A(
        oc8051_sfr1_oc8051_int1_n96), .B(wr_dat[2]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n95) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u90 ( .A0(
        oc8051_sfr1_oc8051_int1_n86), .A1(oc8051_sfr1_oc8051_int1_n94), .B0(
        oc8051_sfr1_oc8051_int1_n95), .Y(oc8051_sfr1_oc8051_int1_n256) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u89 ( .A(oc8051_sfr1_tr0), .B(
        oc8051_sfr1_oc8051_int1_n91), .Y(oc8051_sfr1_oc8051_int1_n93) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u88 ( .A(
        oc8051_sfr1_oc8051_int1_n93), .B(wr_dat[4]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n92) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u87 ( .A0(
        oc8051_sfr1_oc8051_int1_n86), .A1(oc8051_sfr1_oc8051_int1_n91), .B0(
        oc8051_sfr1_oc8051_int1_n92), .Y(oc8051_sfr1_oc8051_int1_n257) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u86 ( .A(oc8051_sfr1_tr1), .B(
        oc8051_sfr1_oc8051_int1_n87), .Y(oc8051_sfr1_oc8051_int1_n89) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u85 ( .A(
        oc8051_sfr1_oc8051_int1_n89), .B(wr_dat[6]), .S0(
        oc8051_sfr1_oc8051_int1_n90), .Y(oc8051_sfr1_oc8051_int1_n88) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u84 ( .A0(
        oc8051_sfr1_oc8051_int1_n86), .A1(oc8051_sfr1_oc8051_int1_n87), .B0(
        oc8051_sfr1_oc8051_int1_n88), .Y(oc8051_sfr1_oc8051_int1_n258) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u83 ( .A(wr_addr[6]), .Y(
        oc8051_sfr1_oc8051_int1_n85) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u82 ( .A(
        oc8051_sfr1_oc8051_int1_n85), .B(wr_addr[7]), .C(wr_addr[5]), .D(
        n_5_net_), .Y(oc8051_sfr1_oc8051_int1_n50) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u81 ( .AN(wr_addr[4]), .B(
        oc8051_sfr1_oc8051_int1_n84), .C(wr_addr[3]), .D(
        oc8051_sfr1_oc8051_int1_n50), .Y(oc8051_sfr1_oc8051_int1_n63) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u80 ( .A(oc8051_sfr1_oc8051_int1_n63), .Y(oc8051_sfr1_oc8051_int1_n58) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u79 ( .A(wr_addr[3]), .B(
        oc8051_sfr1_oc8051_int1_n50), .C(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_int1_n42) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u78 ( .AN(
        oc8051_sfr1_oc8051_int1_n42), .B(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_int1_n80) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u77 ( .A(
        oc8051_sfr1_oc8051_int1_n80), .B(descy), .Y(
        oc8051_sfr1_oc8051_int1_n64) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u76 ( .A(oc8051_sfr1_oc8051_int1_n64), .Y(oc8051_sfr1_oc8051_int1_n59) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u75 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[0]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n81) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u74 ( .A(oc8051_sfr1_ie_0_), .Y(
        oc8051_sfr1_oc8051_int1_n82) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u73 ( .AN(
        oc8051_sfr1_oc8051_int1_n80), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n62) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u72 ( .A0(
        oc8051_sfr1_oc8051_int1_n62), .A1(oc8051_sfr1_oc8051_int1_n36), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n83) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u71 ( .A(
        oc8051_sfr1_oc8051_int1_n81), .B(oc8051_sfr1_oc8051_int1_n82), .S0(
        oc8051_sfr1_oc8051_int1_n83), .Y(oc8051_sfr1_oc8051_int1_n259) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u70 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[1]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n77) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u69 ( .A(oc8051_sfr1_ie_1_), .Y(
        oc8051_sfr1_oc8051_int1_n78) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u68 ( .AN(
        oc8051_sfr1_oc8051_int1_n80), .B(oc8051_sfr1_oc8051_int1_n38), .Y(
        oc8051_sfr1_oc8051_int1_n57) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u67 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n36), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n79) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u66 ( .A(
        oc8051_sfr1_oc8051_int1_n77), .B(oc8051_sfr1_oc8051_int1_n78), .S0(
        oc8051_sfr1_oc8051_int1_n79), .Y(oc8051_sfr1_oc8051_int1_n260) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u65 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[2]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n74) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u64 ( .A0(
        oc8051_sfr1_oc8051_int1_n62), .A1(oc8051_sfr1_oc8051_int1_n29), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n76) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u63 ( .A(
        oc8051_sfr1_oc8051_int1_n74), .B(oc8051_sfr1_oc8051_int1_n75), .S0(
        oc8051_sfr1_oc8051_int1_n76), .Y(oc8051_sfr1_oc8051_int1_n261) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u62 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[3]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n71) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u61 ( .A(oc8051_sfr1_ie_3_), .Y(
        oc8051_sfr1_oc8051_int1_n72) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u60 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n29), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n73) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u59 ( .A(
        oc8051_sfr1_oc8051_int1_n71), .B(oc8051_sfr1_oc8051_int1_n72), .S0(
        oc8051_sfr1_oc8051_int1_n73), .Y(oc8051_sfr1_oc8051_int1_n262) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u58 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[4]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n68) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u57 ( .A(oc8051_sfr1_ie_4_), .Y(
        oc8051_sfr1_oc8051_int1_n69) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u56 ( .A0(
        oc8051_sfr1_oc8051_int1_n62), .A1(oc8051_sfr1_oc8051_int1_n21), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n70) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u55 ( .A(
        oc8051_sfr1_oc8051_int1_n68), .B(oc8051_sfr1_oc8051_int1_n69), .S0(
        oc8051_sfr1_oc8051_int1_n70), .Y(oc8051_sfr1_oc8051_int1_n263) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u54 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[5]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n65) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u53 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n21), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n67) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u52 ( .A(
        oc8051_sfr1_oc8051_int1_n65), .B(oc8051_sfr1_oc8051_int1_n66), .S0(
        oc8051_sfr1_oc8051_int1_n67), .Y(oc8051_sfr1_oc8051_int1_n264) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u51 ( .A(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_int1_n18) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u50 ( .A0(
        oc8051_sfr1_oc8051_int1_n18), .A1(oc8051_sfr1_oc8051_int1_n63), .B0(
        oc8051_sfr1_oc8051_int1_n64), .Y(oc8051_sfr1_oc8051_int1_n60) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u49 ( .A0(
        oc8051_sfr1_oc8051_int1_n62), .A1(oc8051_sfr1_oc8051_int1_n11), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n61) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u48 ( .A(
        oc8051_sfr1_oc8051_int1_n60), .B(oc8051_sfr1_ie_6_), .S0(
        oc8051_sfr1_oc8051_int1_n61), .Y(oc8051_sfr1_oc8051_int1_n265) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u47 ( .A0(
        oc8051_sfr1_oc8051_int1_n58), .A1(wr_dat[7]), .B0(
        oc8051_sfr1_oc8051_int1_n59), .Y(oc8051_sfr1_oc8051_int1_n54) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u46 ( .A0(
        oc8051_sfr1_oc8051_int1_n57), .A1(oc8051_sfr1_oc8051_int1_n11), .B0(
        oc8051_sfr1_oc8051_int1_n58), .Y(oc8051_sfr1_oc8051_int1_n56) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u45 ( .A(
        oc8051_sfr1_oc8051_int1_n54), .B(oc8051_sfr1_oc8051_int1_n55), .S0(
        oc8051_sfr1_oc8051_int1_n56), .Y(oc8051_sfr1_oc8051_int1_n266) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u44 ( .A(
        oc8051_sfr1_oc8051_int1_n11), .B(wr_addr[4]), .C(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n51) );
  NAND4B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u43 ( .AN(wr_addr[3]), .B(
        oc8051_sfr1_oc8051_int1_n44), .C(oc8051_sfr1_oc8051_int1_n50), .D(
        oc8051_sfr1_oc8051_int1_n51), .Y(oc8051_sfr1_oc8051_int1_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u42 ( .A(oc8051_sfr1_oc8051_int1_n17), .Y(oc8051_sfr1_oc8051_int1_n12) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u41 ( .A(
        oc8051_sfr1_oc8051_int1_n42), .B(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_int1_n37) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_int1_u40 ( .A(descy), .B(
        oc8051_sfr1_oc8051_int1_n37), .Y(oc8051_sfr1_oc8051_int1_n13) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u39 ( .A(oc8051_sfr1_oc8051_int1_n13), .Y(oc8051_sfr1_oc8051_int1_n22) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u38 ( .A0(wr_dat[0]), .A1(
        oc8051_sfr1_oc8051_int1_n12), .B0(oc8051_sfr1_oc8051_int1_n22), .Y(
        oc8051_sfr1_oc8051_int1_n39) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u37 ( .A(oc8051_sfr1_ip_0_), .Y(
        oc8051_sfr1_oc8051_int1_n40) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u36 ( .AN(
        oc8051_sfr1_oc8051_int1_n37), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_int1_n16) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u35 ( .A0(
        oc8051_sfr1_oc8051_int1_n36), .A1(oc8051_sfr1_oc8051_int1_n16), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n41) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u34 ( .A(
        oc8051_sfr1_oc8051_int1_n39), .B(oc8051_sfr1_oc8051_int1_n40), .S0(
        oc8051_sfr1_oc8051_int1_n41), .Y(oc8051_sfr1_oc8051_int1_n267) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u33 ( .A0(wr_dat[1]), .A1(
        oc8051_sfr1_oc8051_int1_n12), .B0(oc8051_sfr1_oc8051_int1_n22), .Y(
        oc8051_sfr1_oc8051_int1_n33) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u32 ( .A(oc8051_sfr1_ip_1_), .Y(
        oc8051_sfr1_oc8051_int1_n34) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u31 ( .AN(
        oc8051_sfr1_oc8051_int1_n37), .B(oc8051_sfr1_oc8051_int1_n38), .Y(
        oc8051_sfr1_oc8051_int1_n10) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u30 ( .A0(
        oc8051_sfr1_oc8051_int1_n36), .A1(oc8051_sfr1_oc8051_int1_n10), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n35) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u29 ( .A(
        oc8051_sfr1_oc8051_int1_n33), .B(oc8051_sfr1_oc8051_int1_n34), .S0(
        oc8051_sfr1_oc8051_int1_n35), .Y(oc8051_sfr1_oc8051_int1_n268) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u28 ( .A0(wr_dat[2]), .A1(
        oc8051_sfr1_oc8051_int1_n12), .B0(oc8051_sfr1_oc8051_int1_n22), .Y(
        oc8051_sfr1_oc8051_int1_n30) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u27 ( .A(oc8051_sfr1_ip_2_), .Y(
        oc8051_sfr1_oc8051_int1_n31) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u26 ( .A0(
        oc8051_sfr1_oc8051_int1_n29), .A1(oc8051_sfr1_oc8051_int1_n16), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n32) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u25 ( .A(
        oc8051_sfr1_oc8051_int1_n30), .B(oc8051_sfr1_oc8051_int1_n31), .S0(
        oc8051_sfr1_oc8051_int1_n32), .Y(oc8051_sfr1_oc8051_int1_n269) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u24 ( .A0(wr_dat[3]), .A1(
        oc8051_sfr1_oc8051_int1_n12), .B0(oc8051_sfr1_oc8051_int1_n22), .Y(
        oc8051_sfr1_oc8051_int1_n26) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u23 ( .A0(
        oc8051_sfr1_oc8051_int1_n29), .A1(oc8051_sfr1_oc8051_int1_n10), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n28) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u22 ( .A(
        oc8051_sfr1_oc8051_int1_n26), .B(oc8051_sfr1_oc8051_int1_n27), .S0(
        oc8051_sfr1_oc8051_int1_n28), .Y(oc8051_sfr1_oc8051_int1_n270) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u21 ( .A0(wr_dat[4]), .A1(
        oc8051_sfr1_oc8051_int1_n12), .B0(oc8051_sfr1_oc8051_int1_n22), .Y(
        oc8051_sfr1_oc8051_int1_n23) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u20 ( .A(oc8051_sfr1_ip_4_), .Y(
        oc8051_sfr1_oc8051_int1_n24) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u19 ( .A0(
        oc8051_sfr1_oc8051_int1_n21), .A1(oc8051_sfr1_oc8051_int1_n16), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n25) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u18 ( .A(
        oc8051_sfr1_oc8051_int1_n23), .B(oc8051_sfr1_oc8051_int1_n24), .S0(
        oc8051_sfr1_oc8051_int1_n25), .Y(oc8051_sfr1_oc8051_int1_n271) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u17 ( .A0(wr_dat[5]), .A1(
        oc8051_sfr1_oc8051_int1_n12), .B0(oc8051_sfr1_oc8051_int1_n22), .Y(
        oc8051_sfr1_oc8051_int1_n19) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u16 ( .A0(
        oc8051_sfr1_oc8051_int1_n21), .A1(oc8051_sfr1_oc8051_int1_n10), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n20) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u15 ( .A(
        oc8051_sfr1_oc8051_int1_n19), .B(oc8051_sfr1_oc8051_int1_n9), .S0(
        oc8051_sfr1_oc8051_int1_n20), .Y(oc8051_sfr1_oc8051_int1_n272) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u14 ( .A0(
        oc8051_sfr1_oc8051_int1_n17), .A1(oc8051_sfr1_oc8051_int1_n18), .B0(
        oc8051_sfr1_oc8051_int1_n13), .Y(oc8051_sfr1_oc8051_int1_n14) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u13 ( .A0(
        oc8051_sfr1_oc8051_int1_n16), .A1(oc8051_sfr1_oc8051_int1_n11), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n15) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u12 ( .A(
        oc8051_sfr1_oc8051_int1_n14), .B(oc8051_sfr1_ip_6_), .S0(
        oc8051_sfr1_oc8051_int1_n15), .Y(oc8051_sfr1_oc8051_int1_n273) );
  AO1B2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u11 ( .B0(
        oc8051_sfr1_oc8051_int1_n12), .B1(wr_dat[7]), .A0N(
        oc8051_sfr1_oc8051_int1_n13), .Y(oc8051_sfr1_oc8051_int1_n2) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u10 ( .A0(
        oc8051_sfr1_oc8051_int1_n10), .A1(oc8051_sfr1_oc8051_int1_n11), .B0(
        oc8051_sfr1_oc8051_int1_n12), .Y(oc8051_sfr1_oc8051_int1_n3) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u9 ( .A(oc8051_sfr1_oc8051_int1_n2), 
        .B(oc8051_sfr1_ip_7_), .S0(oc8051_sfr1_oc8051_int1_n3), .Y(
        oc8051_sfr1_oc8051_int1_n274) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u8 ( .A(oc8051_sfr1_oc8051_int1_n4), 
        .Y(int_src[0]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u7 ( .A(oc8051_sfr1_oc8051_int1_n5), 
        .Y(int_src[1]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u6 ( .A(oc8051_sfr1_oc8051_int1_n6), 
        .Y(int_src[3]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_int1_u5 ( .A(oc8051_sfr1_oc8051_int1_n9), 
        .Y(oc8051_sfr1_ip_5_) );
  INV_X0P5M_A12TS oc8051_sfr1_oc8051_int1_u4 ( .A(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_int1_n120) );
  TIELO_X1M_A12TS oc8051_sfr1_oc8051_int1_u3 ( .Y(
        oc8051_sfr1_oc8051_int1_int_vec_2_) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_5_ ( .D(
        oc8051_sfr1_oc8051_int1_n272), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n9) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n244), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n4) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n242), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n6) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n243), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n5) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_0__1_ ( .D(
        oc8051_sfr1_oc8051_int1_n237), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n48) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_0__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n239), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n49) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_0__2_ ( .D(
        oc8051_sfr1_oc8051_int1_n235), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n47) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_1__1_ ( .D(
        oc8051_sfr1_oc8051_int1_n236), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n45) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_1__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n238), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n46) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_isrc_reg_1__2_ ( .D(
        oc8051_sfr1_oc8051_int1_n253), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n43) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_4_ ( .D(
        oc8051_sfr1_oc8051_int1_n241), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n7) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_vec_reg_5_ ( .D(
        oc8051_sfr1_oc8051_int1_n240), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n8) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_lev_reg_0__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n246), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n53) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_int1_int_lev_reg_1__0_ ( .D(
        oc8051_sfr1_oc8051_int1_n245), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_int1_n52) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_dept_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n247), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_dept_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_4_ ( .D(
        oc8051_sfr1_oc8051_int1_n263), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_proc_reg ( .D(
        oc8051_sfr1_oc8051_int1_n248), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_proc) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_2_ ( .D(
        oc8051_sfr1_oc8051_int1_n261), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_ie1_reg ( .D(
        oc8051_sfr1_oc8051_int1_n250), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n259), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_2_ ( .D(
        oc8051_sfr1_oc8051_int1_n269), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_ie0_reg ( .D(
        oc8051_sfr1_oc8051_int1_n251), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n258), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tr1) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n255), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_tf1_reg ( .D(
        oc8051_sfr1_oc8051_int1_n254), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n268), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_0_ ( .D(
        oc8051_sfr1_oc8051_int1_n267), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_4_ ( .D(
        oc8051_sfr1_oc8051_int1_n271), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_4_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n260), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n262), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_7_ ( .D(
        oc8051_sfr1_oc8051_int1_n266), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_tf0_reg ( .D(
        oc8051_sfr1_oc8051_int1_n252), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n256), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tcon_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_int_dept_reg_1_ ( .D(
        oc8051_sfr1_oc8051_int1_n249), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_int1_int_dept_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tcon_s_reg_2_ ( .D(
        oc8051_sfr1_oc8051_int1_n257), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tr0) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_5_ ( .D(
        oc8051_sfr1_oc8051_int1_n264), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_5_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_3_ ( .D(
        oc8051_sfr1_oc8051_int1_n270), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_6_ ( .D(
        oc8051_sfr1_oc8051_int1_n273), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie_reg_6_ ( .D(
        oc8051_sfr1_oc8051_int1_n265), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ie_6_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ip_reg_7_ ( .D(
        oc8051_sfr1_oc8051_int1_n274), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_ip_7_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie1_buff_reg ( .D(int1_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_ie1_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_ie0_buff_reg ( .D(int0_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_ie0_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tf0_buff_reg ( .D(oc8051_sfr1_tf0), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_tf0_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_int1_tf1_buff_reg ( .D(oc8051_sfr1_tf1), 
        .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_int1_tf1_buff) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u245 ( .A(oc8051_sfr1_tmod[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u244 ( .A(oc8051_sfr1_tmod[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n79) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u243 ( .A(
        oc8051_sfr1_oc8051_tc1_n159), .B(oc8051_sfr1_oc8051_tc1_n79), .Y(
        oc8051_sfr1_oc8051_tc1_n20) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u242 ( .A(oc8051_sfr1_pres_ow), .B(
        oc8051_sfr1_oc8051_tc1_n20), .C(oc8051_sfr1_tr1), .Y(
        oc8051_sfr1_oc8051_tc1_n16) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u241 ( .A(oc8051_sfr1_tmod[0]), .B(
        oc8051_sfr1_tmod[1]), .Y(oc8051_sfr1_oc8051_tc1_n28) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u240 ( .A(oc8051_sfr1_tmod[3]), .B(
        int0_i), .Y(oc8051_sfr1_oc8051_tc1_n162) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u239 ( .A(oc8051_sfr1_pres_ow), .Y(
        oc8051_sfr1_oc8051_tc1_n154) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u238 ( .AN(t0_i), .B(
        oc8051_sfr1_oc8051_tc1_t0_buff), .Y(oc8051_sfr1_oc8051_tc1_n164) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u237 ( .A(
        oc8051_sfr1_oc8051_tc1_n154), .B(oc8051_sfr1_oc8051_tc1_n164), .S0(
        oc8051_sfr1_tmod[2]), .Y(oc8051_sfr1_oc8051_tc1_n163) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u236 ( .A(oc8051_sfr1_tr0), .B(
        oc8051_sfr1_oc8051_tc1_n162), .C(oc8051_sfr1_oc8051_tc1_n163), .Y(
        oc8051_sfr1_oc8051_tc1_n75) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u235 ( .A(oc8051_sfr1_oc8051_tc1_n75), 
        .Y(oc8051_sfr1_oc8051_tc1_n69) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u234 ( .A(
        oc8051_sfr1_oc8051_tc1_n28), .B(oc8051_sfr1_oc8051_tc1_n69), .Y(
        oc8051_sfr1_oc8051_tc1_n161) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u233 ( .A(
        oc8051_sfr1_oc8051_tc1_n159), .B(oc8051_sfr1_tmod[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n27) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u232 ( .A(
        oc8051_sfr1_oc8051_tc1_n27), .B(oc8051_sfr1_oc8051_tc1_n69), .Y(
        oc8051_sfr1_oc8051_tc1_n66) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u231 ( .A(
        oc8051_sfr1_oc8051_tc1_n161), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_n42) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u230 ( .A(oc8051_sfr1_tl0[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n43) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u229 ( .A0(
        oc8051_sfr1_oc8051_tc1_n223), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n43), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_0) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u228 ( .A(oc8051_sfr1_tl0[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n49) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u227 ( .A0(
        oc8051_sfr1_oc8051_tc1_n222), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n49), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_1) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u226 ( .A0(
        oc8051_sfr1_oc8051_tc1_n218), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n221), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_10) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u225 ( .A0(
        oc8051_sfr1_oc8051_tc1_n217), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n220), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_11) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u224 ( .A0(
        oc8051_sfr1_oc8051_tc1_n216), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n219), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_12) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u223 ( .A(
        oc8051_sfr1_oc8051_tc1_n218), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_13) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u222 ( .A(
        oc8051_sfr1_oc8051_tc1_n217), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_14) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u221 ( .A(
        oc8051_sfr1_oc8051_tc1_n216), .B(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_15) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u220 ( .A(oc8051_sfr1_tl0[2]), .Y(
        oc8051_sfr1_oc8051_tc1_n52) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u219 ( .A0(
        oc8051_sfr1_oc8051_tc1_n221), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n52), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_2) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u218 ( .A(oc8051_sfr1_tl0[3]), .Y(
        oc8051_sfr1_oc8051_tc1_n55) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u217 ( .A0(
        oc8051_sfr1_oc8051_tc1_n220), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n55), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_3) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u216 ( .A(oc8051_sfr1_tl0[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n58) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u215 ( .A0(
        oc8051_sfr1_oc8051_tc1_n219), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n42), .B1(oc8051_sfr1_oc8051_tc1_n58), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_4) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u214 ( .A(oc8051_sfr1_tl0[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n61) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u213 ( .A0(
        oc8051_sfr1_oc8051_tc1_n223), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n61), .B1(oc8051_sfr1_oc8051_tc1_n66), .C0(
        oc8051_sfr1_oc8051_tc1_n218), .C1(oc8051_sfr1_oc8051_tc1_n16), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_5) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u212 ( .A(oc8051_sfr1_tl0[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n64) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u211 ( .A0(
        oc8051_sfr1_oc8051_tc1_n222), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n64), .B1(oc8051_sfr1_oc8051_tc1_n66), .C0(
        oc8051_sfr1_oc8051_tc1_n217), .C1(oc8051_sfr1_oc8051_tc1_n16), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_6) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u210 ( .A(oc8051_sfr1_tl0[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n1) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u209 ( .A0(
        oc8051_sfr1_oc8051_tc1_n221), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n1), .B1(oc8051_sfr1_oc8051_tc1_n66), .C0(
        oc8051_sfr1_oc8051_tc1_n216), .C1(oc8051_sfr1_oc8051_tc1_n16), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_7) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u208 ( .A0(
        oc8051_sfr1_oc8051_tc1_n220), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n223), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_8) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u207 ( .A0(
        oc8051_sfr1_oc8051_tc1_n219), .A1(oc8051_sfr1_oc8051_tc1_n161), .B0(
        oc8051_sfr1_oc8051_tc1_n222), .B1(oc8051_sfr1_oc8051_tc1_n66), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_9) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u206 ( .A(oc8051_sfr1_th1[5]), .B(
        oc8051_sfr1_th1[2]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_10) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u205 ( .A(oc8051_sfr1_th1[6]), .B(
        oc8051_sfr1_th1[3]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_11) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u204 ( .A(oc8051_sfr1_th1[7]), .B(
        oc8051_sfr1_th1[4]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_12) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u203 ( .A(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n120) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u202 ( .A(oc8051_sfr1_th1[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n140) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u201 ( .A(
        oc8051_sfr1_oc8051_tc1_n120), .B(oc8051_sfr1_oc8051_tc1_n140), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_13) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u200 ( .A(oc8051_sfr1_th1[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n113) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u199 ( .A(
        oc8051_sfr1_oc8051_tc1_n120), .B(oc8051_sfr1_oc8051_tc1_n113), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_14) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u198 ( .A(oc8051_sfr1_th1[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n87) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u197 ( .A(oc8051_sfr1_oc8051_tc1_n87), .B(oc8051_sfr1_oc8051_tc1_n120), .Y(oc8051_sfr1_oc8051_tc1_u3_u8_z_15) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u196 ( .A(oc8051_sfr1_th1[0]), .B(
        oc8051_sfr1_tl1[5]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_5) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u195 ( .A(oc8051_sfr1_th1[1]), .B(
        oc8051_sfr1_tl1[6]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_6) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u194 ( .A(oc8051_sfr1_th1[2]), .B(
        oc8051_sfr1_tl1[7]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_7) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u193 ( .A(oc8051_sfr1_th1[3]), .B(
        oc8051_sfr1_th1[0]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_8) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u192 ( .A(oc8051_sfr1_th1[4]), .B(
        oc8051_sfr1_th1[1]), .S0(oc8051_sfr1_tmod[4]), .Y(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_9) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u191 ( .A(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n26) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u190 ( .AN(n_5_net_), .B(
        oc8051_sfr1_wr_bit_r), .Y(oc8051_sfr1_oc8051_tc1_n157) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u189 ( .A(wr_addr[4]), .B(wr_addr[6]), .C(wr_addr[5]), .Y(oc8051_sfr1_oc8051_tc1_n160) );
  AND3_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u188 ( .A(wr_addr[7]), .B(wr_addr[3]), .C(oc8051_sfr1_oc8051_tc1_n160), .Y(oc8051_sfr1_oc8051_tc1_n156) );
  NAND3B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u187 ( .AN(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_tc1_n157), .C(oc8051_sfr1_oc8051_tc1_n156), .Y(
        oc8051_sfr1_oc8051_tc1_n80) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u186 ( .A(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n83) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u185 ( .A(oc8051_sfr1_oc8051_tc1_n80), .B(wr_addr[1]), .C(oc8051_sfr1_oc8051_tc1_n83), .Y(
        oc8051_sfr1_oc8051_tc1_n158) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u184 ( .A(
        oc8051_sfr1_oc8051_tc1_n159), .B(oc8051_sfr1_oc8051_tc1_n26), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n224) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u183 ( .A(
        oc8051_sfr1_oc8051_tc1_n79), .B(oc8051_sfr1_oc8051_tc1_n30), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n225) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u182 ( .A(oc8051_sfr1_tmod[2]), .B(
        wr_dat[2]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n226) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u181 ( .A(oc8051_sfr1_tmod[3]), .B(
        wr_dat[3]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n227) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u180 ( .A(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n36) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u179 ( .A(
        oc8051_sfr1_oc8051_tc1_n120), .B(oc8051_sfr1_oc8051_tc1_n36), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n228) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u178 ( .A(oc8051_sfr1_tmod[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n92) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u177 ( .A(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n38) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u176 ( .A(
        oc8051_sfr1_oc8051_tc1_n92), .B(oc8051_sfr1_oc8051_tc1_n38), .S0(
        oc8051_sfr1_oc8051_tc1_n158), .Y(oc8051_sfr1_oc8051_tc1_n229) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u175 ( .A(oc8051_sfr1_tmod[6]), .B(
        wr_dat[6]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n230) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u174 ( .A(oc8051_sfr1_tmod[7]), .B(
        wr_dat[7]), .S0(oc8051_sfr1_oc8051_tc1_n158), .Y(
        oc8051_sfr1_oc8051_tc1_n231) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u173 ( .A(wr_addr[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n81) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u172 ( .A(oc8051_sfr1_oc8051_tc1_n81), .B(oc8051_sfr1_oc8051_tc1_n80), .C(oc8051_sfr1_oc8051_tc1_n83), .Y(
        oc8051_sfr1_oc8051_tc1_n90) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u171 ( .A(wr_addr[2]), .B(
        oc8051_sfr1_oc8051_tc1_n156), .C(oc8051_sfr1_oc8051_tc1_n157), .D(
        oc8051_sfr1_oc8051_tc1_n81), .Y(oc8051_sfr1_oc8051_tc1_n82) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u170 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_tc1_n82), .Y(oc8051_sfr1_oc8051_tc1_n114) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u169 ( .A(oc8051_sfr1_oc8051_tc1_n114), .Y(oc8051_sfr1_oc8051_tc1_n99) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u168 ( .A(oc8051_sfr1_oc8051_tc1_n90), .B(oc8051_sfr1_oc8051_tc1_n99), .Y(oc8051_sfr1_oc8051_tc1_n119) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u167 ( .A(oc8051_sfr1_oc8051_tc1_n90), 
        .Y(oc8051_sfr1_oc8051_tc1_n125) );
  NAND2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u166 ( .AN(t1_i), .B(
        oc8051_sfr1_oc8051_tc1_t1_buff), .Y(oc8051_sfr1_oc8051_tc1_n155) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u165 ( .A(
        oc8051_sfr1_oc8051_tc1_n154), .B(oc8051_sfr1_oc8051_tc1_n155), .S0(
        oc8051_sfr1_tmod[6]), .Y(oc8051_sfr1_oc8051_tc1_n152) );
  AOI21B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u164 ( .A0(oc8051_sfr1_tmod[7]), 
        .A1(int1_i), .B0N(oc8051_sfr1_tr1), .Y(oc8051_sfr1_oc8051_tc1_n153) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u163 ( .A(
        oc8051_sfr1_oc8051_tc1_n152), .B(oc8051_sfr1_oc8051_tc1_n119), .C(
        oc8051_sfr1_oc8051_tc1_n153), .Y(oc8051_sfr1_oc8051_tc1_n122) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u162 ( .A(
        oc8051_sfr1_oc8051_tc1_n125), .B(oc8051_sfr1_oc8051_tc1_n122), .Y(
        oc8051_sfr1_oc8051_tc1_n124) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u161 ( .A(
        oc8051_sfr1_oc8051_tc1_n119), .B(oc8051_sfr1_oc8051_tc1_n124), .Y(
        oc8051_sfr1_oc8051_tc1_n138) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u160 ( .A(oc8051_sfr1_oc8051_tc1_n174), .Y(oc8051_sfr1_oc8051_tc1_n110) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u159 ( .A(oc8051_sfr1_tmod[5]), .B(
        oc8051_sfr1_oc8051_tc1_n110), .Y(oc8051_sfr1_oc8051_tc1_n151) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u158 ( .A(
        oc8051_sfr1_oc8051_tc1_n192), .B(oc8051_sfr1_oc8051_tc1_n151), .S0(
        oc8051_sfr1_oc8051_tc1_n120), .Y(oc8051_sfr1_oc8051_tc1_n146) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u157 ( .A(
        oc8051_sfr1_oc8051_tc1_n233), .B(oc8051_sfr1_oc8051_tc1_n99), .Y(
        oc8051_sfr1_oc8051_tc1_n148) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u156 ( .A(oc8051_sfr1_tl1[3]), .B(
        oc8051_sfr1_tl1[2]), .C(oc8051_sfr1_tl1[1]), .D(oc8051_sfr1_tl1[0]), 
        .Y(oc8051_sfr1_oc8051_tc1_n149) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u155 ( .A(oc8051_sfr1_tl1[7]), .B(
        oc8051_sfr1_tl1[6]), .C(oc8051_sfr1_tl1[5]), .D(oc8051_sfr1_tl1[4]), 
        .Y(oc8051_sfr1_oc8051_tc1_n150) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u154 ( .A(
        oc8051_sfr1_oc8051_tc1_n149), .B(oc8051_sfr1_oc8051_tc1_n150), .Y(
        oc8051_sfr1_oc8051_tc1_n145) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u153 ( .A(oc8051_sfr1_tmod[5]), .B(
        oc8051_sfr1_oc8051_tc1_n119), .C(oc8051_sfr1_oc8051_tc1_n145), .Y(
        oc8051_sfr1_oc8051_tc1_n86) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u152 ( .A(oc8051_sfr1_oc8051_tc1_n86), 
        .Y(oc8051_sfr1_oc8051_tc1_n127) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u151 ( .A(
        oc8051_sfr1_oc8051_tc1_n148), .B(oc8051_sfr1_oc8051_tc1_n127), .S0(
        oc8051_sfr1_oc8051_tc1_n124), .Y(oc8051_sfr1_oc8051_tc1_n147) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u150 ( .A0(
        oc8051_sfr1_oc8051_tc1_n138), .A1(oc8051_sfr1_oc8051_tc1_n146), .B0(
        oc8051_sfr1_oc8051_tc1_n147), .Y(oc8051_sfr1_oc8051_tc1_n234) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u149 ( .A(oc8051_sfr1_oc8051_tc1_n92), .B(oc8051_sfr1_oc8051_tc1_n145), .Y(oc8051_sfr1_oc8051_tc1_n91) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u148 ( .A0(
        oc8051_sfr1_oc8051_tc1_n202), .A1(oc8051_sfr1_oc8051_tc1_n91), .B0(
        oc8051_sfr1_oc8051_tc1_n167), .B1(oc8051_sfr1_oc8051_tc1_n92), .Y(
        oc8051_sfr1_oc8051_tc1_n142) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u147 ( .A0(
        oc8051_sfr1_oc8051_tc1_n92), .A1(oc8051_sfr1_oc8051_tc1_n120), .B0(
        oc8051_sfr1_oc8051_tc1_n122), .C0(oc8051_sfr1_oc8051_tc1_n125), .Y(
        oc8051_sfr1_oc8051_tc1_n144) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u146 ( .A(
        oc8051_sfr1_oc8051_tc1_n119), .B(oc8051_sfr1_oc8051_tc1_n144), .Y(
        oc8051_sfr1_oc8051_tc1_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u145 ( .A(oc8051_sfr1_oc8051_tc1_n144), .Y(oc8051_sfr1_oc8051_tc1_n89) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u144 ( .A0(
        oc8051_sfr1_oc8051_tc1_n89), .A1(oc8051_sfr1_tl1[6]), .B0(
        oc8051_sfr1_oc8051_tc1_n90), .B1(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n143) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u143 ( .A0(
        oc8051_sfr1_oc8051_tc1_n142), .A1(oc8051_sfr1_oc8051_tc1_n85), .B0(
        oc8051_sfr1_oc8051_tc1_n86), .B1(oc8051_sfr1_oc8051_tc1_n113), .C0(
        oc8051_sfr1_oc8051_tc1_n143), .Y(oc8051_sfr1_oc8051_tc1_n235) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u142 ( .A0(
        oc8051_sfr1_oc8051_tc1_n201), .A1(oc8051_sfr1_oc8051_tc1_n91), .B0(
        oc8051_sfr1_oc8051_tc1_n166), .B1(oc8051_sfr1_oc8051_tc1_n92), .Y(
        oc8051_sfr1_oc8051_tc1_n139) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u141 ( .A0(
        oc8051_sfr1_oc8051_tc1_n89), .A1(oc8051_sfr1_tl1[5]), .B0(
        oc8051_sfr1_oc8051_tc1_n90), .B1(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc1_n141) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u140 ( .A0(
        oc8051_sfr1_oc8051_tc1_n139), .A1(oc8051_sfr1_oc8051_tc1_n85), .B0(
        oc8051_sfr1_oc8051_tc1_n86), .B1(oc8051_sfr1_oc8051_tc1_n140), .C0(
        oc8051_sfr1_oc8051_tc1_n141), .Y(oc8051_sfr1_oc8051_tc1_n236) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u139 ( .A(oc8051_sfr1_tl1[4]), .Y(
        oc8051_sfr1_oc8051_tc1_n136) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u138 ( .AN(
        oc8051_sfr1_oc8051_tc1_n91), .B(oc8051_sfr1_oc8051_tc1_n138), .Y(
        oc8051_sfr1_oc8051_tc1_n128) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u137 ( .A(oc8051_sfr1_oc8051_tc1_n92), .B(oc8051_sfr1_tmod[4]), .Y(oc8051_sfr1_oc8051_tc1_n121) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u136 ( .A(
        oc8051_sfr1_oc8051_tc1_n138), .B(oc8051_sfr1_oc8051_tc1_n121), .Y(
        oc8051_sfr1_oc8051_tc1_n129) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u135 ( .A0(oc8051_sfr1_th1[4]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n200), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n165), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n137) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u134 ( .A0(
        oc8051_sfr1_oc8051_tc1_n136), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n36), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n137), .Y(oc8051_sfr1_oc8051_tc1_n237) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u133 ( .A(oc8051_sfr1_tl1[3]), .Y(
        oc8051_sfr1_oc8051_tc1_n134) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u132 ( .A(wr_dat[3]), .Y(
        oc8051_sfr1_oc8051_tc1_n34) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u131 ( .A0(oc8051_sfr1_th1[3]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n199), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1640), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n135) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u130 ( .A0(
        oc8051_sfr1_oc8051_tc1_n134), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n34), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n135), .Y(oc8051_sfr1_oc8051_tc1_n238) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u129 ( .A(oc8051_sfr1_tl1[2]), .Y(
        oc8051_sfr1_oc8051_tc1_n132) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u128 ( .A(wr_dat[2]), .Y(
        oc8051_sfr1_oc8051_tc1_n32) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u127 ( .A0(oc8051_sfr1_th1[2]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n198), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1630), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n133) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u126 ( .A0(
        oc8051_sfr1_oc8051_tc1_n132), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n32), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n133), .Y(oc8051_sfr1_oc8051_tc1_n239) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u125 ( .A(oc8051_sfr1_tl1[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n130) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u124 ( .A0(oc8051_sfr1_th1[1]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n197), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1620), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n131) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u123 ( .A0(
        oc8051_sfr1_oc8051_tc1_n130), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n30), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n131), .Y(oc8051_sfr1_oc8051_tc1_n240) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u122 ( .A(oc8051_sfr1_tl1[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n123) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u121 ( .A0(oc8051_sfr1_th1[0]), 
        .A1(oc8051_sfr1_oc8051_tc1_n127), .B0(oc8051_sfr1_oc8051_tc1_n196), 
        .B1(oc8051_sfr1_oc8051_tc1_n128), .C0(oc8051_sfr1_oc8051_tc1_n1610), 
        .C1(oc8051_sfr1_oc8051_tc1_n129), .Y(oc8051_sfr1_oc8051_tc1_n126) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u120 ( .A0(
        oc8051_sfr1_oc8051_tc1_n123), .A1(oc8051_sfr1_oc8051_tc1_n124), .B0(
        oc8051_sfr1_oc8051_tc1_n26), .B1(oc8051_sfr1_oc8051_tc1_n125), .C0(
        oc8051_sfr1_oc8051_tc1_n126), .Y(oc8051_sfr1_oc8051_tc1_n241) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u119 ( .A0(
        oc8051_sfr1_oc8051_tc1_n121), .A1(oc8051_sfr1_oc8051_tc1_n122), .B0(
        oc8051_sfr1_oc8051_tc1_n114), .Y(oc8051_sfr1_oc8051_tc1_n112) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u118 ( .A(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n9) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u117 ( .A(
        oc8051_sfr1_oc8051_tc1_n112), .B(oc8051_sfr1_oc8051_tc1_n120), .C(
        oc8051_sfr1_oc8051_tc1_n119), .Y(oc8051_sfr1_oc8051_tc1_n93) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u116 ( .A(oc8051_sfr1_oc8051_tc1_n93), 
        .Y(oc8051_sfr1_oc8051_tc1_n116) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u115 ( .A(
        oc8051_sfr1_oc8051_tc1_n119), .B(oc8051_sfr1_oc8051_tc1_n112), .C(
        oc8051_sfr1_tmod[4]), .Y(oc8051_sfr1_oc8051_tc1_n95) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u114 ( .A(oc8051_sfr1_oc8051_tc1_n95), 
        .Y(oc8051_sfr1_oc8051_tc1_n117) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u113 ( .A0(
        oc8051_sfr1_oc8051_tc1_n173), .A1(oc8051_sfr1_oc8051_tc1_n116), .B0(
        oc8051_sfr1_oc8051_tc1_n191), .B1(oc8051_sfr1_oc8051_tc1_n117), .Y(
        oc8051_sfr1_oc8051_tc1_n118) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u112 ( .A0(
        oc8051_sfr1_oc8051_tc1_n87), .A1(oc8051_sfr1_oc8051_tc1_n112), .B0(
        oc8051_sfr1_oc8051_tc1_n9), .B1(oc8051_sfr1_oc8051_tc1_n114), .C0(
        oc8051_sfr1_oc8051_tc1_n118), .Y(oc8051_sfr1_oc8051_tc1_n242) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u111 ( .A(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc1_n40) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u110 ( .A0(
        oc8051_sfr1_oc8051_tc1_n172), .A1(oc8051_sfr1_oc8051_tc1_n116), .B0(
        oc8051_sfr1_oc8051_tc1_n190), .B1(oc8051_sfr1_oc8051_tc1_n117), .Y(
        oc8051_sfr1_oc8051_tc1_n115) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u109 ( .A0(
        oc8051_sfr1_oc8051_tc1_n112), .A1(oc8051_sfr1_oc8051_tc1_n113), .B0(
        oc8051_sfr1_oc8051_tc1_n40), .B1(oc8051_sfr1_oc8051_tc1_n114), .C0(
        oc8051_sfr1_oc8051_tc1_n115), .Y(oc8051_sfr1_oc8051_tc1_n243) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u108 ( .A(oc8051_sfr1_oc8051_tc1_n171), .Y(oc8051_sfr1_oc8051_tc1_n104) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u107 ( .A(oc8051_sfr1_oc8051_tc1_n112), .Y(oc8051_sfr1_oc8051_tc1_n98) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u106 ( .A0(oc8051_sfr1_th1[5]), 
        .A1(oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[5]), .Y(oc8051_sfr1_oc8051_tc1_n111) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u105 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n104), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n110), .C0(
        oc8051_sfr1_oc8051_tc1_n111), .Y(oc8051_sfr1_oc8051_tc1_n244) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u104 ( .A(oc8051_sfr1_oc8051_tc1_n170), .Y(oc8051_sfr1_oc8051_tc1_n101) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u103 ( .A(oc8051_sfr1_oc8051_tc1_n173), .Y(oc8051_sfr1_oc8051_tc1_n108) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u102 ( .A0(oc8051_sfr1_th1[4]), 
        .A1(oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[4]), .Y(oc8051_sfr1_oc8051_tc1_n109) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u101 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n101), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n108), .C0(
        oc8051_sfr1_oc8051_tc1_n109), .Y(oc8051_sfr1_oc8051_tc1_n245) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u100 ( .A(oc8051_sfr1_oc8051_tc1_n169), .Y(oc8051_sfr1_oc8051_tc1_n96) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u99 ( .A(oc8051_sfr1_oc8051_tc1_n172), 
        .Y(oc8051_sfr1_oc8051_tc1_n106) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u98 ( .A0(oc8051_sfr1_th1[3]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[3]), .Y(oc8051_sfr1_oc8051_tc1_n107) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u97 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n96), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n106), .C0(
        oc8051_sfr1_oc8051_tc1_n107), .Y(oc8051_sfr1_oc8051_tc1_n246) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u96 ( .A(oc8051_sfr1_oc8051_tc1_n168), 
        .Y(oc8051_sfr1_oc8051_tc1_n103) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u95 ( .A0(oc8051_sfr1_th1[2]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[2]), .Y(oc8051_sfr1_oc8051_tc1_n105) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u94 ( .A0(
        oc8051_sfr1_oc8051_tc1_n103), .A1(oc8051_sfr1_oc8051_tc1_n93), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n104), .C0(
        oc8051_sfr1_oc8051_tc1_n105), .Y(oc8051_sfr1_oc8051_tc1_n247) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u93 ( .A(oc8051_sfr1_oc8051_tc1_n167), 
        .Y(oc8051_sfr1_oc8051_tc1_n100) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u92 ( .A0(oc8051_sfr1_th1[1]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[1]), .Y(oc8051_sfr1_oc8051_tc1_n102) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u91 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n100), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n101), .C0(
        oc8051_sfr1_oc8051_tc1_n102), .Y(oc8051_sfr1_oc8051_tc1_n248) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u90 ( .A(oc8051_sfr1_oc8051_tc1_n166), 
        .Y(oc8051_sfr1_oc8051_tc1_n94) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u89 ( .A0(oc8051_sfr1_th1[0]), .A1(
        oc8051_sfr1_oc8051_tc1_n98), .B0(oc8051_sfr1_oc8051_tc1_n99), .B1(
        wr_dat[0]), .Y(oc8051_sfr1_oc8051_tc1_n97) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u88 ( .A0(
        oc8051_sfr1_oc8051_tc1_n93), .A1(oc8051_sfr1_oc8051_tc1_n94), .B0(
        oc8051_sfr1_oc8051_tc1_n95), .B1(oc8051_sfr1_oc8051_tc1_n96), .C0(
        oc8051_sfr1_oc8051_tc1_n97), .Y(oc8051_sfr1_oc8051_tc1_n249) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u87 ( .A0(
        oc8051_sfr1_oc8051_tc1_n203), .A1(oc8051_sfr1_oc8051_tc1_n91), .B0(
        oc8051_sfr1_oc8051_tc1_n168), .B1(oc8051_sfr1_oc8051_tc1_n92), .Y(
        oc8051_sfr1_oc8051_tc1_n84) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u86 ( .A0(
        oc8051_sfr1_oc8051_tc1_n89), .A1(oc8051_sfr1_tl1[7]), .B0(
        oc8051_sfr1_oc8051_tc1_n90), .B1(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n88) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u85 ( .A0(
        oc8051_sfr1_oc8051_tc1_n84), .A1(oc8051_sfr1_oc8051_tc1_n85), .B0(
        oc8051_sfr1_oc8051_tc1_n86), .B1(oc8051_sfr1_oc8051_tc1_n87), .C0(
        oc8051_sfr1_oc8051_tc1_n88), .Y(oc8051_sfr1_oc8051_tc1_n250) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u84 ( .A0(
        oc8051_sfr1_oc8051_tc1_n920), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n630), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n600), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n76) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u83 ( .A(oc8051_sfr1_oc8051_tc1_n82), .B(oc8051_sfr1_oc8051_tc1_n83), .Y(oc8051_sfr1_oc8051_tc1_n25) );
  OR3_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u82 ( .A(oc8051_sfr1_oc8051_tc1_n80), 
        .B(wr_addr[0]), .C(oc8051_sfr1_oc8051_tc1_n81), .Y(
        oc8051_sfr1_oc8051_tc1_n8) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u81 ( .A(oc8051_sfr1_oc8051_tc1_n25), .B(oc8051_sfr1_oc8051_tc1_n8), .Y(oc8051_sfr1_oc8051_tc1_n15) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u80 ( .A(oc8051_sfr1_oc8051_tc1_n79), 
        .B(oc8051_sfr1_tmod[0]), .Y(oc8051_sfr1_oc8051_tc1_n68) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u79 ( .A(oc8051_sfr1_oc8051_tc1_n15), 
        .Y(oc8051_sfr1_oc8051_tc1_n21) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u78 ( .A(oc8051_sfr1_tl0[3]), .B(
        oc8051_sfr1_tl0[2]), .C(oc8051_sfr1_tl0[1]), .D(oc8051_sfr1_tl0[0]), 
        .Y(oc8051_sfr1_oc8051_tc1_n77) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u77 ( .A(oc8051_sfr1_tl0[7]), .B(
        oc8051_sfr1_tl0[6]), .C(oc8051_sfr1_tl0[5]), .D(oc8051_sfr1_tl0[4]), 
        .Y(oc8051_sfr1_oc8051_tc1_n78) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u76 ( .A(oc8051_sfr1_oc8051_tc1_n77), 
        .B(oc8051_sfr1_oc8051_tc1_n78), .Y(oc8051_sfr1_oc8051_tc1_n71) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u75 ( .A(oc8051_sfr1_oc8051_tc1_n68), .B(oc8051_sfr1_oc8051_tc1_n21), .C(oc8051_sfr1_oc8051_tc1_n71), .Y(
        oc8051_sfr1_oc8051_tc1_n10) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u74 ( .A0(
        oc8051_sfr1_oc8051_tc1_n76), .A1(oc8051_sfr1_oc8051_tc1_n15), .B0(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n73) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u73 ( .A0(
        oc8051_sfr1_oc8051_tc1_n75), .A1(oc8051_sfr1_oc8051_tc1_n15), .B0(
        oc8051_sfr1_oc8051_tc1_n8), .Y(oc8051_sfr1_oc8051_tc1_n45) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u72 ( .AN(
        oc8051_sfr1_oc8051_tc1_n25), .B(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n74) );
  MXT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u71 ( .A(oc8051_sfr1_oc8051_tc1_n73), 
        .B(oc8051_sfr1_tf0), .S0(oc8051_sfr1_oc8051_tc1_n74), .Y(
        oc8051_sfr1_oc8051_tc1_n251) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u70 ( .A(oc8051_sfr1_oc8051_tc1_n27), 
        .Y(oc8051_sfr1_oc8051_tc1_n18) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u69 ( .A(oc8051_sfr1_oc8051_tc1_n15), 
        .B(oc8051_sfr1_oc8051_tc1_n18), .Y(oc8051_sfr1_oc8051_tc1_n4) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u68 ( .A(oc8051_sfr1_oc8051_tc1_n68), 
        .Y(oc8051_sfr1_oc8051_tc1_n19) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u67 ( .A(oc8051_sfr1_oc8051_tc1_n20), 
        .Y(oc8051_sfr1_oc8051_tc1_n72) );
  OA21A1OI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u66 ( .A0(
        oc8051_sfr1_oc8051_tc1_n19), .A1(oc8051_sfr1_oc8051_tc1_n71), .B0(
        oc8051_sfr1_oc8051_tc1_n72), .C0(oc8051_sfr1_oc8051_tc1_n15), .Y(
        oc8051_sfr1_oc8051_tc1_n6) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u65 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n40), .B0(oc8051_sfr1_oc8051_tc1_n217), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n70) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u64 ( .A0(
        oc8051_sfr1_oc8051_tc1_n530), .A1(oc8051_sfr1_oc8051_tc1_n4), .B0(
        oc8051_sfr1_oc8051_tc1_n900), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n70), .Y(oc8051_sfr1_oc8051_tc1_n65) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u63 ( .A0(
        oc8051_sfr1_oc8051_tc1_n68), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n69), .Y(oc8051_sfr1_oc8051_tc1_n67) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u62 ( .A0(
        oc8051_sfr1_oc8051_tc1_n66), .A1(oc8051_sfr1_oc8051_tc1_n67), .B0(
        oc8051_sfr1_oc8051_tc1_n15), .C0(oc8051_sfr1_oc8051_tc1_n8), .Y(
        oc8051_sfr1_oc8051_tc1_n3) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u61 ( .A(oc8051_sfr1_oc8051_tc1_n64), .B(oc8051_sfr1_oc8051_tc1_n65), .S0(oc8051_sfr1_oc8051_tc1_n3), .Y(
        oc8051_sfr1_oc8051_tc1_n252) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u60 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n38), .B0(oc8051_sfr1_oc8051_tc1_n218), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n63) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u59 ( .A0(
        oc8051_sfr1_oc8051_tc1_n520), .A1(oc8051_sfr1_oc8051_tc1_n4), .B0(
        oc8051_sfr1_oc8051_tc1_n890), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n63), .Y(oc8051_sfr1_oc8051_tc1_n62) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u58 ( .A(oc8051_sfr1_oc8051_tc1_n61), .B(oc8051_sfr1_oc8051_tc1_n62), .S0(oc8051_sfr1_oc8051_tc1_n3), .Y(
        oc8051_sfr1_oc8051_tc1_n253) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u57 ( .A(oc8051_sfr1_oc8051_tc1_n28), 
        .Y(oc8051_sfr1_oc8051_tc1_n17) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u56 ( .A0(
        oc8051_sfr1_oc8051_tc1_n17), .A1(oc8051_sfr1_oc8051_tc1_n18), .B0(
        oc8051_sfr1_oc8051_tc1_n15), .Y(oc8051_sfr1_oc8051_tc1_n46) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u55 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n36), .B0(oc8051_sfr1_oc8051_tc1_n219), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n60) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u54 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n510), .B0(
        oc8051_sfr1_oc8051_tc1_n880), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n60), .Y(oc8051_sfr1_oc8051_tc1_n59) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u53 ( .A(oc8051_sfr1_oc8051_tc1_n58), .B(oc8051_sfr1_oc8051_tc1_n59), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n254) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u52 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n34), .B0(oc8051_sfr1_oc8051_tc1_n220), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n57) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u51 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n500), .B0(
        oc8051_sfr1_oc8051_tc1_n870), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n57), .Y(oc8051_sfr1_oc8051_tc1_n56) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u50 ( .A(oc8051_sfr1_oc8051_tc1_n55), .B(oc8051_sfr1_oc8051_tc1_n56), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n255) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u49 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n32), .B0(oc8051_sfr1_oc8051_tc1_n221), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n54) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u48 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n490), .B0(
        oc8051_sfr1_oc8051_tc1_n860), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n54), .Y(oc8051_sfr1_oc8051_tc1_n53) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u47 ( .A(oc8051_sfr1_oc8051_tc1_n52), .B(oc8051_sfr1_oc8051_tc1_n53), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n256) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u46 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n30), .B0(oc8051_sfr1_oc8051_tc1_n222), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n51) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u45 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n480), .B0(
        oc8051_sfr1_oc8051_tc1_n850), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n51), .Y(oc8051_sfr1_oc8051_tc1_n50) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u44 ( .A(oc8051_sfr1_oc8051_tc1_n49), .B(oc8051_sfr1_oc8051_tc1_n50), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n257) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u43 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_0), .Y(oc8051_sfr1_oc8051_tc1_n47) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u42 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n26), .B0(oc8051_sfr1_oc8051_tc1_n223), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n48) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u41 ( .A0(
        oc8051_sfr1_oc8051_tc1_n46), .A1(oc8051_sfr1_oc8051_tc1_n47), .B0(
        oc8051_sfr1_oc8051_tc1_n840), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n48), .Y(oc8051_sfr1_oc8051_tc1_n44) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u40 ( .A(oc8051_sfr1_oc8051_tc1_n43), .B(oc8051_sfr1_oc8051_tc1_n44), .S0(oc8051_sfr1_oc8051_tc1_n45), .Y(
        oc8051_sfr1_oc8051_tc1_n258) );
  AO21A1AI2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u39 ( .A0(
        oc8051_sfr1_oc8051_tc1_n42), .A1(oc8051_sfr1_oc8051_tc1_n16), .B0(
        oc8051_sfr1_oc8051_tc1_n15), .C0(oc8051_sfr1_oc8051_tc1_n25), .Y(
        oc8051_sfr1_oc8051_tc1_n22) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u38 ( .A0(
        oc8051_sfr1_oc8051_tc1_n20), .A1(oc8051_sfr1_oc8051_tc1_n540), .B0(
        oc8051_sfr1_oc8051_tc1_n620), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n590), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n41) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u37 ( .A(oc8051_sfr1_oc8051_tc1_n21), .B(oc8051_sfr1_oc8051_tc1_n22), .Y(oc8051_sfr1_oc8051_tc1_n24) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u36 ( .A0(
        oc8051_sfr1_oc8051_tc1_n216), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n41), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n9), .C1(oc8051_sfr1_oc8051_tc1_n25), .Y(
        oc8051_sfr1_oc8051_tc1_n259) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u35 ( .A0(
        oc8051_sfr1_oc8051_tc1_n530), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n610), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n580), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n39) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u34 ( .A0(
        oc8051_sfr1_oc8051_tc1_n217), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n39), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n40), .Y(
        oc8051_sfr1_oc8051_tc1_n260) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u33 ( .A0(
        oc8051_sfr1_oc8051_tc1_n520), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n600), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n570), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n37) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u32 ( .A0(
        oc8051_sfr1_oc8051_tc1_n218), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n37), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n38), .Y(
        oc8051_sfr1_oc8051_tc1_n261) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u31 ( .A0(
        oc8051_sfr1_oc8051_tc1_n510), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n590), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n560), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n35) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u30 ( .A0(
        oc8051_sfr1_oc8051_tc1_n219), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n35), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n36), .Y(
        oc8051_sfr1_oc8051_tc1_n262) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u29 ( .A0(
        oc8051_sfr1_oc8051_tc1_n500), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n580), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n28), .C1(oc8051_sfr1_oc8051_tc1_n550), .Y(
        oc8051_sfr1_oc8051_tc1_n33) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u28 ( .A0(
        oc8051_sfr1_oc8051_tc1_n220), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n33), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n34), .Y(
        oc8051_sfr1_oc8051_tc1_n263) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u27 ( .A0(
        oc8051_sfr1_oc8051_tc1_n490), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n570), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n28), .C1(oc8051_sfr1_oc8051_tc1_n540), .Y(
        oc8051_sfr1_oc8051_tc1_n31) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u26 ( .A0(
        oc8051_sfr1_oc8051_tc1_n221), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n31), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n32), .Y(
        oc8051_sfr1_oc8051_tc1_n264) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u25 ( .A0(
        oc8051_sfr1_oc8051_tc1_n480), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n560), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n530), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n29) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u24 ( .A0(
        oc8051_sfr1_oc8051_tc1_n222), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n29), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n30), .Y(
        oc8051_sfr1_oc8051_tc1_n265) );
  AOI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u23 ( .A0(
        oc8051_sfr1_oc8051_tc1_n470), .A1(oc8051_sfr1_oc8051_tc1_n20), .B0(
        oc8051_sfr1_oc8051_tc1_n550), .B1(oc8051_sfr1_oc8051_tc1_n27), .C0(
        oc8051_sfr1_oc8051_tc1_n520), .C1(oc8051_sfr1_oc8051_tc1_n28), .Y(
        oc8051_sfr1_oc8051_tc1_n23) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u22 ( .A0(
        oc8051_sfr1_oc8051_tc1_n223), .A1(oc8051_sfr1_oc8051_tc1_n22), .B0(
        oc8051_sfr1_oc8051_tc1_n23), .B1(oc8051_sfr1_oc8051_tc1_n24), .C0(
        oc8051_sfr1_oc8051_tc1_n25), .C1(oc8051_sfr1_oc8051_tc1_n26), .Y(
        oc8051_sfr1_oc8051_tc1_n266) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u21 ( .A(oc8051_sfr1_oc8051_tc1_n20), .B(oc8051_sfr1_oc8051_tc1_n21), .C(oc8051_sfr1_oc8051_tc1_n550), .Y(
        oc8051_sfr1_oc8051_tc1_n11) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u20 ( .A(oc8051_sfr1_oc8051_tc1_n17), .B(oc8051_sfr1_oc8051_tc1_n18), .C(oc8051_sfr1_oc8051_tc1_n19), .Y(
        oc8051_sfr1_oc8051_tc1_n13) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u19 ( .A(oc8051_sfr1_oc8051_tc1_n16), 
        .Y(oc8051_sfr1_oc8051_tc1_n14) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u18 ( .A(oc8051_sfr1_oc8051_tc1_n13), 
        .B(oc8051_sfr1_oc8051_tc1_n14), .C(oc8051_sfr1_oc8051_tc1_n15), .Y(
        oc8051_sfr1_oc8051_tc1_n12) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u17 ( .A(oc8051_sfr1_oc8051_tc1_n11), .B(oc8051_sfr1_oc8051_tc1_n232), .S0(oc8051_sfr1_oc8051_tc1_n12), .Y(
        oc8051_sfr1_oc8051_tc1_n267) );
  OAI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u16 ( .A0(oc8051_sfr1_oc8051_tc1_n8), .A1(oc8051_sfr1_oc8051_tc1_n9), .B0(oc8051_sfr1_oc8051_tc1_n216), .B1(
        oc8051_sfr1_oc8051_tc1_n10), .Y(oc8051_sfr1_oc8051_tc1_n7) );
  AOI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u15 ( .A0(
        oc8051_sfr1_oc8051_tc1_n540), .A1(oc8051_sfr1_oc8051_tc1_n4), .B0(
        oc8051_sfr1_oc8051_tc1_n910), .B1(oc8051_sfr1_oc8051_tc1_n6), .C0(
        oc8051_sfr1_oc8051_tc1_n7), .Y(oc8051_sfr1_oc8051_tc1_n2) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u14 ( .A(oc8051_sfr1_oc8051_tc1_n1), 
        .B(oc8051_sfr1_oc8051_tc1_n2), .S0(oc8051_sfr1_oc8051_tc1_n3), .Y(
        oc8051_sfr1_oc8051_tc1_n268) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u13 ( .A(oc8051_sfr1_oc8051_tc1_n216), 
        .Y(oc8051_sfr1_th0[7]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u12 ( .A(oc8051_sfr1_oc8051_tc1_n217), 
        .Y(oc8051_sfr1_th0[6]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u11 ( .A(oc8051_sfr1_oc8051_tc1_n218), 
        .Y(oc8051_sfr1_th0[5]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u10 ( .A(oc8051_sfr1_oc8051_tc1_n219), 
        .Y(oc8051_sfr1_th0[4]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u9 ( .A(oc8051_sfr1_oc8051_tc1_n220), 
        .Y(oc8051_sfr1_th0[3]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u8 ( .A(oc8051_sfr1_oc8051_tc1_n221), 
        .Y(oc8051_sfr1_th0[2]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u7 ( .A(oc8051_sfr1_oc8051_tc1_n222), 
        .Y(oc8051_sfr1_th0[1]) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc1_u6 ( .A(oc8051_sfr1_oc8051_tc1_n223), 
        .Y(oc8051_sfr1_th0[0]) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc1_u5 ( .A(oc8051_sfr1_oc8051_tc1_n233), .B(oc8051_sfr1_oc8051_tc1_n232), .Y(oc8051_sfr1_tf1) );
  TIELO_X1M_A12TS oc8051_sfr1_oc8051_tc1_u4 ( .Y(oc8051_sfr1_oc8051_tc1_n5) );
  INV_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_u3 ( .A(wr_dat[1]), .Y(
        oc8051_sfr1_oc8051_tc1_n30) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n259), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n216) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n260), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n217) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n261), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n218) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n264), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n221) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n265), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n222) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n266), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n223) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n262), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n219) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_th0_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n263), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n220) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n241), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n228), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[4]) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_tf1_0_reg ( .D(
        oc8051_sfr1_oc8051_tc1_n267), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n232) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc1_tf1_1_reg ( .D(
        oc8051_sfr1_oc8051_tc1_n234), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc1_n233) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n238), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n237), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n240), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n239), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n258), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n236), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n235), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n255), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n268), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n254), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n253), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n257), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n256), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl0_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n252), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl0[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tl1_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n250), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl1[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc1_n245), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n246), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n247), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n248), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n249), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n229), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc1_n224), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc1_n225), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc1_n244), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc1_n226), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n230), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc1_n227), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n242), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_th1_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc1_n243), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th1[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tmod_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc1_n231), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tmod[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_tf0_reg ( .D(
        oc8051_sfr1_oc8051_tc1_n251), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tf0) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_t1_buff_reg ( .D(t1_i), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc1_t1_buff) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc1_t0_buff_reg ( .D(t0_i), .CK(wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc1_t0_buff) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1 ( .A(oc8051_sfr1_tl1[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n1610) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_13 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_13), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[13]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[14]), .S(oc8051_sfr1_oc8051_tc1_n174) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_14 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_14), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[14]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[15]), .S(oc8051_sfr1_oc8051_tc1_n190) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_15 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_15), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[15]), .CO(
        oc8051_sfr1_oc8051_tc1_n192), .S(oc8051_sfr1_oc8051_tc1_n191) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_5 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_5), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[6]), .S(oc8051_sfr1_oc8051_tc1_n166)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_6 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_6), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[7]), .S(oc8051_sfr1_oc8051_tc1_n167)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_7 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_7), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[8]), .S(oc8051_sfr1_oc8051_tc1_n168)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_8 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_8), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[8]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[9]), .S(oc8051_sfr1_oc8051_tc1_n169)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_9 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_9), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[9]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[10]), .S(oc8051_sfr1_oc8051_tc1_n170) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_10 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_10), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[10]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[11]), .S(oc8051_sfr1_oc8051_tc1_n171) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_11 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_11), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[11]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[12]), .S(oc8051_sfr1_oc8051_tc1_n172) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_12 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u8_z_12), .B(
        oc8051_sfr1_oc8051_tc1_r372_carry[12]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[13]), .S(oc8051_sfr1_oc8051_tc1_n173) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_1 ( .A(oc8051_sfr1_tl1[1]), 
        .B(oc8051_sfr1_tl1[0]), .CO(oc8051_sfr1_oc8051_tc1_r372_carry[2]), .S(
        oc8051_sfr1_oc8051_tc1_n1620) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_3 ( .A(oc8051_sfr1_tl1[3]), 
        .B(oc8051_sfr1_oc8051_tc1_r372_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[4]), .S(oc8051_sfr1_oc8051_tc1_n1640) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_2 ( .A(oc8051_sfr1_tl1[2]), 
        .B(oc8051_sfr1_oc8051_tc1_r372_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[3]), .S(oc8051_sfr1_oc8051_tc1_n1630) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r372_u1_1_4 ( .A(oc8051_sfr1_tl1[4]), 
        .B(oc8051_sfr1_oc8051_tc1_r372_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_r372_carry[5]), .S(oc8051_sfr1_oc8051_tc1_n165)
         );
  XOR2_X0P5M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u2 ( .A(
        oc8051_sfr1_oc8051_tc1_add_220_carry[7]), .B(oc8051_sfr1_tl1[7]), .Y(
        oc8051_sfr1_oc8051_tc1_n203) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1 ( .A(oc8051_sfr1_tl1[0]), 
        .Y(oc8051_sfr1_oc8051_tc1_n196) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_1 ( .A(oc8051_sfr1_tl1[1]), .B(oc8051_sfr1_tl1[0]), .CO(oc8051_sfr1_oc8051_tc1_add_220_carry[2]), .S(
        oc8051_sfr1_oc8051_tc1_n197) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_3 ( .A(oc8051_sfr1_tl1[3]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[4]), .S(
        oc8051_sfr1_oc8051_tc1_n199) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_2 ( .A(oc8051_sfr1_tl1[2]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[3]), .S(
        oc8051_sfr1_oc8051_tc1_n198) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_4 ( .A(oc8051_sfr1_tl1[4]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[5]), .S(
        oc8051_sfr1_oc8051_tc1_n200) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_5 ( .A(oc8051_sfr1_tl1[5]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[6]), .S(
        oc8051_sfr1_oc8051_tc1_n201) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_add_220_u1_1_6 ( .A(oc8051_sfr1_tl1[6]), .B(oc8051_sfr1_oc8051_tc1_add_220_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_add_220_carry[7]), .S(
        oc8051_sfr1_oc8051_tc1_n202) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1 ( .A(oc8051_sfr1_tl0[0]), .Y(
        oc8051_sfr1_oc8051_tc1_n840) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_1 ( .A(oc8051_sfr1_tl0[1]), 
        .B(oc8051_sfr1_tl0[0]), .CO(oc8051_sfr1_oc8051_tc1_r364_carry[2]), .S(
        oc8051_sfr1_oc8051_tc1_n850) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_2 ( .A(oc8051_sfr1_tl0[2]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[3]), .S(oc8051_sfr1_oc8051_tc1_n860)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_3 ( .A(oc8051_sfr1_tl0[3]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[4]), .S(oc8051_sfr1_oc8051_tc1_n870)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_4 ( .A(oc8051_sfr1_tl0[4]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[5]), .S(oc8051_sfr1_oc8051_tc1_n880)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_5 ( .A(oc8051_sfr1_tl0[5]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[6]), .S(oc8051_sfr1_oc8051_tc1_n890)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_6 ( .A(oc8051_sfr1_tl0[6]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_r364_carry[7]), .S(oc8051_sfr1_oc8051_tc1_n900)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r364_u1_1_7 ( .A(oc8051_sfr1_tl0[7]), 
        .B(oc8051_sfr1_oc8051_tc1_r364_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc1_n920), .S(oc8051_sfr1_oc8051_tc1_n910) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_0), .Y(oc8051_sfr1_oc8051_tc1_n470) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_1 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_1), .B(oc8051_sfr1_oc8051_tc1_u3_u1_z_0), .CO(oc8051_sfr1_oc8051_tc1_r360_carry[2]), .S(oc8051_sfr1_oc8051_tc1_n480)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_5 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_5), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[6]), .S(oc8051_sfr1_oc8051_tc1_n520)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_6 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_6), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[7]), .S(oc8051_sfr1_oc8051_tc1_n530)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_7 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_7), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[8]), .S(oc8051_sfr1_oc8051_tc1_n540)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_2 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_2), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[3]), .S(oc8051_sfr1_oc8051_tc1_n490)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_3 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_3), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[4]), .S(oc8051_sfr1_oc8051_tc1_n500)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_4 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_4), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[5]), .S(oc8051_sfr1_oc8051_tc1_n510)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_9 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_9), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[9]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[10]), .S(oc8051_sfr1_oc8051_tc1_n560) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_10 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_10), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[10]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[11]), .S(oc8051_sfr1_oc8051_tc1_n570) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_11 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_11), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[11]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[12]), .S(oc8051_sfr1_oc8051_tc1_n580) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_12 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_12), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[12]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[13]), .S(oc8051_sfr1_oc8051_tc1_n590) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_8 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_8), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[8]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[9]), .S(oc8051_sfr1_oc8051_tc1_n550)
         );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_14 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_14), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[14]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[15]), .S(oc8051_sfr1_oc8051_tc1_n610) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_13 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_13), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[13]), .CO(
        oc8051_sfr1_oc8051_tc1_r360_carry[14]), .S(oc8051_sfr1_oc8051_tc1_n600) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc1_r360_u1_1_15 ( .A(
        oc8051_sfr1_oc8051_tc1_u3_u1_z_15), .B(
        oc8051_sfr1_oc8051_tc1_r360_carry[15]), .CO(
        oc8051_sfr1_oc8051_tc1_n630), .S(oc8051_sfr1_oc8051_tc1_n620) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u186 ( .AN(
        oc8051_sfr1_oc8051_tc21_t2ex_r), .B(t2ex_i), .Y(
        oc8051_sfr1_oc8051_tc21_n217) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u185 ( .AN(
        oc8051_sfr1_oc8051_tc21_t2_r), .B(t2_i), .Y(
        oc8051_sfr1_oc8051_tc21_n220) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u184 ( .A(oc8051_sfr1_t2con_3_), 
        .B(oc8051_sfr1_oc8051_tc21_neg_trans), .Y(oc8051_sfr1_oc8051_tc21_n115) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u183 ( .A(oc8051_sfr1_oc8051_tc21_n7), .Y(oc8051_sfr1_tclk) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u182 ( .A(oc8051_sfr1_oc8051_tc21_n8), .Y(oc8051_sfr1_rclk) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u181 ( .A(oc8051_sfr1_tclk), .B(
        oc8051_sfr1_rclk), .Y(oc8051_sfr1_oc8051_tc21_n116) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u180 ( .AN(
        oc8051_sfr1_oc8051_tc21_n116), .B(oc8051_sfr1_t2con_0_), .Y(
        oc8051_sfr1_oc8051_tc21_n11) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u179 ( .A(
        oc8051_sfr1_oc8051_tc21_n11), .Y(oc8051_sfr1_oc8051_tc21_n135) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u178 ( .AN(wr_addr[2]), .B(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_tc21_n34) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u177 ( .A(n_5_net_), .Y(
        oc8051_sfr1_oc8051_tc21_n139) );
  NOR3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u176 ( .A(
        oc8051_sfr1_oc8051_tc21_n139), .B(wr_addr[5]), .C(wr_addr[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n138) );
  AND4_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u175 ( .A(wr_addr[6]), .B(
        wr_addr[3]), .C(wr_addr[7]), .D(oc8051_sfr1_oc8051_tc21_n138), .Y(
        oc8051_sfr1_oc8051_tc21_n127) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u174 ( .AN(
        oc8051_sfr1_oc8051_tc21_n127), .B(oc8051_sfr1_wr_bit_r), .Y(
        oc8051_sfr1_oc8051_tc21_n114) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u173 ( .A(
        oc8051_sfr1_oc8051_tc21_n34), .B(oc8051_sfr1_oc8051_tc21_n114), .C(
        wr_addr[0]), .Y(oc8051_sfr1_oc8051_tc21_n83) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u172 ( .AN(
        oc8051_sfr1_oc8051_tc21_n114), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n113) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u171 ( .A(
        oc8051_sfr1_oc8051_tc21_n113), .B(oc8051_sfr1_oc8051_tc21_n34), .Y(
        oc8051_sfr1_oc8051_tc21_n77) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u170 ( .A(
        oc8051_sfr1_oc8051_tc21_n83), .B(oc8051_sfr1_oc8051_tc21_n77), .Y(
        oc8051_sfr1_oc8051_tc21_n2) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u169 ( .A(oc8051_sfr1_pres_ow), 
        .B(oc8051_sfr1_oc8051_tc21_tc2_event), .S0(oc8051_sfr1_t2con_1_), .Y(
        oc8051_sfr1_oc8051_tc21_n137) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u168 ( .AN(oc8051_sfr1_t2con_2_), 
        .B(oc8051_sfr1_oc8051_tc21_n137), .Y(oc8051_sfr1_oc8051_tc21_n136) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u167 ( .A0(
        oc8051_sfr1_oc8051_tc21_n115), .A1(oc8051_sfr1_oc8051_tc21_n135), .B0(
        oc8051_sfr1_oc8051_tc21_n2), .C0(oc8051_sfr1_oc8051_tc21_n136), .Y(
        oc8051_sfr1_oc8051_tc21_n79) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u166 ( .A(
        oc8051_sfr1_oc8051_tc21_n79), .B(oc8051_sfr1_oc8051_tc21_n116), .Y(
        oc8051_sfr1_oc8051_tc21_n129) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u165 ( .A(oc8051_sfr1_brate2), .B(
        oc8051_sfr1_oc8051_tc21_n850), .S0(oc8051_sfr1_oc8051_tc21_n129), .Y(
        oc8051_sfr1_oc8051_tc21_n128) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u164 ( .A(oc8051_sfr1_tl2[3]), .B(
        oc8051_sfr1_tl2[2]), .C(oc8051_sfr1_tl2[1]), .D(oc8051_sfr1_tl2[0]), 
        .Y(oc8051_sfr1_oc8051_tc21_n131) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u163 ( .A(oc8051_sfr1_tl2[7]), .B(
        oc8051_sfr1_tl2[6]), .C(oc8051_sfr1_tl2[5]), .D(oc8051_sfr1_tl2[4]), 
        .Y(oc8051_sfr1_oc8051_tc21_n132) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u162 ( .A(oc8051_sfr1_th2[3]), .B(
        oc8051_sfr1_th2[2]), .C(oc8051_sfr1_th2[1]), .D(oc8051_sfr1_th2[0]), 
        .Y(oc8051_sfr1_oc8051_tc21_n133) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u161 ( .A(oc8051_sfr1_th2[7]), .B(
        oc8051_sfr1_th2[6]), .C(oc8051_sfr1_th2[5]), .D(oc8051_sfr1_th2[4]), 
        .Y(oc8051_sfr1_oc8051_tc21_n134) );
  OR4_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u160 ( .A(
        oc8051_sfr1_oc8051_tc21_n131), .B(oc8051_sfr1_oc8051_tc21_n132), .C(
        oc8051_sfr1_oc8051_tc21_n133), .D(oc8051_sfr1_oc8051_tc21_n134), .Y(
        oc8051_sfr1_oc8051_tc21_n130) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u159 ( .A(
        oc8051_sfr1_oc8051_tc21_n130), .Y(oc8051_sfr1_oc8051_tc21_n100) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u158 ( .A(
        oc8051_sfr1_oc8051_tc21_n129), .B(oc8051_sfr1_oc8051_tc21_n100), .Y(
        oc8051_sfr1_oc8051_tc21_n101) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u157 ( .A(
        oc8051_sfr1_oc8051_tc21_n128), .B(oc8051_sfr1_oc8051_tc21_n101), .Y(
        oc8051_sfr1_oc8051_tc21_n150) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u156 ( .A(wr_addr[2]), .B(
        wr_addr[1]), .Y(oc8051_sfr1_oc8051_tc21_n19) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u155 ( .A(
        oc8051_sfr1_oc8051_tc21_n19), .B(oc8051_sfr1_oc8051_tc21_n113), .Y(
        oc8051_sfr1_oc8051_tc21_n17) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u154 ( .A(
        oc8051_sfr1_oc8051_tc21_n17), .Y(oc8051_sfr1_oc8051_tc21_n122) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u153 ( .A(oc8051_sfr1_wr_bit_r), 
        .B(oc8051_sfr1_oc8051_tc21_n127), .Y(oc8051_sfr1_oc8051_tc21_n121) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u152 ( .A(
        oc8051_sfr1_oc8051_tc21_n121), .Y(oc8051_sfr1_oc8051_tc21_n120) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u151 ( .A(descy), .B(
        oc8051_sfr1_oc8051_tc21_n120), .Y(oc8051_sfr1_oc8051_tc21_n14) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u150 ( .A0(
        oc8051_sfr1_oc8051_tc21_n122), .A1(oc8051_sfr1_oc8051_tc21_n120), .B0(
        oc8051_sfr1_oc8051_tc21_n14), .Y(oc8051_sfr1_oc8051_tc21_n123) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u149 ( .A0(wr_dat[7]), .A1(
        oc8051_sfr1_oc8051_tc21_n122), .B0(oc8051_sfr1_oc8051_tc21_n123), .Y(
        oc8051_sfr1_oc8051_tc21_n124) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u148 ( .AN(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_tc21_n121), .Y(oc8051_sfr1_oc8051_tc21_n23) );
  AOI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u147 ( .A0(
        oc8051_sfr1_oc8051_tc21_tf2_set), .A1(oc8051_sfr1_oc8051_tc21_n121), 
        .B0(oc8051_sfr1_oc8051_tc21_n122), .C0(oc8051_sfr1_oc8051_tc21_n126), 
        .Y(oc8051_sfr1_oc8051_tc21_n125) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u146 ( .A(
        oc8051_sfr1_oc8051_tc21_n124), .B(oc8051_sfr1_oc8051_tc21_n6), .S0(
        oc8051_sfr1_oc8051_tc21_n125), .Y(oc8051_sfr1_oc8051_tc21_n151) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u145 ( .A0(wr_dat[6]), .A1(
        oc8051_sfr1_oc8051_tc21_n122), .B0(oc8051_sfr1_oc8051_tc21_n123), .Y(
        oc8051_sfr1_oc8051_tc21_n117) );
  NOR2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u144 ( .A(
        oc8051_sfr1_oc8051_tc21_n121), .B(wr_addr[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n18) );
  OAI31_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u143 ( .A0(
        oc8051_sfr1_oc8051_tc21_n115), .A1(oc8051_sfr1_oc8051_tc21_tf2_set), 
        .A2(oc8051_sfr1_oc8051_tc21_n120), .B0(oc8051_sfr1_oc8051_tc21_n17), 
        .Y(oc8051_sfr1_oc8051_tc21_n119) );
  AOI31_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u142 ( .A0(
        oc8051_sfr1_oc8051_tc21_n18), .A1(wr_addr[2]), .A2(wr_addr[1]), .B0(
        oc8051_sfr1_oc8051_tc21_n119), .Y(oc8051_sfr1_oc8051_tc21_n118) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u141 ( .A(
        oc8051_sfr1_oc8051_tc21_n117), .B(oc8051_sfr1_oc8051_tc21_n5), .S0(
        oc8051_sfr1_oc8051_tc21_n118), .Y(oc8051_sfr1_oc8051_tc21_n152) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u140 ( .A(oc8051_sfr1_th2[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n97) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u139 ( .A(oc8051_sfr1_t2con_0_), 
        .B(oc8051_sfr1_oc8051_tc21_n116), .Y(oc8051_sfr1_oc8051_tc21_n99) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u138 ( .A(
        oc8051_sfr1_oc8051_tc21_n99), .Y(oc8051_sfr1_oc8051_tc21_n10) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u137 ( .A(
        oc8051_sfr1_oc8051_tc21_n115), .Y(oc8051_sfr1_oc8051_tc21_n102) );
  NOR2B_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u136 ( .AN(wr_addr[1]), .B(
        wr_addr[2]), .Y(oc8051_sfr1_oc8051_tc21_n27) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u135 ( .A(wr_addr[0]), .B(
        oc8051_sfr1_oc8051_tc21_n114), .C(oc8051_sfr1_oc8051_tc21_n27), .Y(
        oc8051_sfr1_oc8051_tc21_n105) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u134 ( .A(
        oc8051_sfr1_oc8051_tc21_n27), .B(oc8051_sfr1_oc8051_tc21_n113), .Y(
        oc8051_sfr1_oc8051_tc21_n43) );
  NAND4_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u133 ( .A(
        oc8051_sfr1_oc8051_tc21_n10), .B(oc8051_sfr1_oc8051_tc21_n102), .C(
        oc8051_sfr1_oc8051_tc21_n105), .D(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n39) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u132 ( .A(oc8051_sfr1_rcap2h[7]), 
        .Y(oc8051_sfr1_oc8051_tc21_n112) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u131 ( .A(
        oc8051_sfr1_oc8051_tc21_n105), .B(oc8051_sfr1_oc8051_tc21_n39), .Y(
        oc8051_sfr1_oc8051_tc21_n104) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u130 ( .A(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n64) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u129 ( .A0(
        oc8051_sfr1_oc8051_tc21_n97), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n112), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n64), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n153) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u128 ( .A(oc8051_sfr1_th2[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n95) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u127 ( .A(oc8051_sfr1_rcap2h[6]), 
        .Y(oc8051_sfr1_oc8051_tc21_n111) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u126 ( .A(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n61) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u125 ( .A0(
        oc8051_sfr1_oc8051_tc21_n95), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n111), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n61), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n154) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u124 ( .A(oc8051_sfr1_th2[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n93) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u123 ( .A(oc8051_sfr1_rcap2h[5]), 
        .Y(oc8051_sfr1_oc8051_tc21_n110) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u122 ( .A(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n58) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u121 ( .A0(
        oc8051_sfr1_oc8051_tc21_n93), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n110), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n58), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n155) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u120 ( .A(oc8051_sfr1_th2[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n91) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u119 ( .A(oc8051_sfr1_rcap2h[4]), 
        .Y(oc8051_sfr1_oc8051_tc21_n109) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u118 ( .A(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n55) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u117 ( .A0(
        oc8051_sfr1_oc8051_tc21_n91), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n109), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n55), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n156) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u116 ( .A(oc8051_sfr1_th2[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n89) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u115 ( .A(oc8051_sfr1_rcap2h[3]), 
        .Y(oc8051_sfr1_oc8051_tc21_n108) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u114 ( .A(wr_dat[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n52) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u113 ( .A0(
        oc8051_sfr1_oc8051_tc21_n89), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n108), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n52), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n157) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u112 ( .A(oc8051_sfr1_th2[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n87) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u111 ( .A(oc8051_sfr1_rcap2h[2]), 
        .Y(oc8051_sfr1_oc8051_tc21_n107) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u110 ( .A(wr_dat[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n49) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u109 ( .A0(
        oc8051_sfr1_oc8051_tc21_n87), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n107), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n49), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n158) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u108 ( .A(oc8051_sfr1_th2[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n85) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u107 ( .A(oc8051_sfr1_rcap2h[1]), 
        .Y(oc8051_sfr1_oc8051_tc21_n106) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u106 ( .A0(
        oc8051_sfr1_oc8051_tc21_n85), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n106), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n46), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n159) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u105 ( .A(oc8051_sfr1_th2[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n81) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u104 ( .A(oc8051_sfr1_rcap2h[0]), 
        .Y(oc8051_sfr1_oc8051_tc21_n103) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u103 ( .A(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n42) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u102 ( .A0(
        oc8051_sfr1_oc8051_tc21_n81), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n103), .B1(oc8051_sfr1_oc8051_tc21_n104), .C0(
        oc8051_sfr1_oc8051_tc21_n42), .C1(oc8051_sfr1_oc8051_tc21_n105), .Y(
        oc8051_sfr1_oc8051_tc21_n160) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u101 ( .A(
        oc8051_sfr1_oc8051_tc21_n11), .B(oc8051_sfr1_oc8051_tc21_n102), .C(
        oc8051_sfr1_oc8051_tc21_n2), .Y(oc8051_sfr1_oc8051_tc21_n80) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u100 ( .A(
        oc8051_sfr1_oc8051_tc21_n79), .B(oc8051_sfr1_oc8051_tc21_n83), .C(
        oc8051_sfr1_oc8051_tc21_n80), .Y(oc8051_sfr1_oc8051_tc21_n82) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u99 ( .A(oc8051_sfr1_oc8051_tc21_n79), .Y(oc8051_sfr1_oc8051_tc21_n12) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u98 ( .A(
        oc8051_sfr1_oc8051_tc21_n100), .B(oc8051_sfr1_oc8051_tc21_n11), .C(
        oc8051_sfr1_oc8051_tc21_n12), .Y(oc8051_sfr1_oc8051_tc21_n9) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u97 ( .A(
        oc8051_sfr1_oc8051_tc21_n101), .B(oc8051_sfr1_oc8051_tc21_n9), .C(
        oc8051_sfr1_oc8051_tc21_n80), .Y(oc8051_sfr1_oc8051_tc21_n78) );
  AOI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u96 ( .A0(
        oc8051_sfr1_oc8051_tc21_n99), .A1(oc8051_sfr1_oc8051_tc21_n100), .B0(
        oc8051_sfr1_oc8051_tc21_n79), .Y(oc8051_sfr1_oc8051_tc21_n68) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u95 ( .A0(oc8051_sfr1_rcap2h[7]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n840), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n98) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u94 ( .A0(
        oc8051_sfr1_oc8051_tc21_n97), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n64), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n98), .Y(oc8051_sfr1_oc8051_tc21_n161) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u93 ( .A0(oc8051_sfr1_rcap2h[6]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n830), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n96) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u92 ( .A0(
        oc8051_sfr1_oc8051_tc21_n95), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n61), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n96), .Y(oc8051_sfr1_oc8051_tc21_n162) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u91 ( .A0(oc8051_sfr1_rcap2h[5]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n820), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n94) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u90 ( .A0(
        oc8051_sfr1_oc8051_tc21_n93), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n58), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n94), .Y(oc8051_sfr1_oc8051_tc21_n163) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u89 ( .A0(oc8051_sfr1_rcap2h[4]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n810), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n92) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u88 ( .A0(
        oc8051_sfr1_oc8051_tc21_n91), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n55), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n92), .Y(oc8051_sfr1_oc8051_tc21_n164) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u87 ( .A0(oc8051_sfr1_rcap2h[3]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n800), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n90) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u86 ( .A0(
        oc8051_sfr1_oc8051_tc21_n89), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n52), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n90), .Y(oc8051_sfr1_oc8051_tc21_n165) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u85 ( .A0(oc8051_sfr1_rcap2h[2]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n790), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n88) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u84 ( .A0(
        oc8051_sfr1_oc8051_tc21_n87), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n49), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n88), .Y(oc8051_sfr1_oc8051_tc21_n166) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u83 ( .A0(oc8051_sfr1_rcap2h[1]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n780), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n86) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u82 ( .A0(
        oc8051_sfr1_oc8051_tc21_n85), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n46), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n86), .Y(oc8051_sfr1_oc8051_tc21_n167) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u81 ( .A0(oc8051_sfr1_rcap2h[0]), 
        .A1(oc8051_sfr1_oc8051_tc21_n78), .B0(oc8051_sfr1_oc8051_tc21_n770), 
        .B1(oc8051_sfr1_oc8051_tc21_n68), .Y(oc8051_sfr1_oc8051_tc21_n84) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u80 ( .A0(
        oc8051_sfr1_oc8051_tc21_n81), .A1(oc8051_sfr1_oc8051_tc21_n82), .B0(
        oc8051_sfr1_oc8051_tc21_n42), .B1(oc8051_sfr1_oc8051_tc21_n83), .C0(
        oc8051_sfr1_oc8051_tc21_n84), .Y(oc8051_sfr1_oc8051_tc21_n168) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u79 ( .A(oc8051_sfr1_tl2[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n62) );
  NAND3_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u78 ( .A(
        oc8051_sfr1_oc8051_tc21_n79), .B(oc8051_sfr1_oc8051_tc21_n77), .C(
        oc8051_sfr1_oc8051_tc21_n80), .Y(oc8051_sfr1_oc8051_tc21_n65) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u77 ( .A(oc8051_sfr1_oc8051_tc21_n78), .Y(oc8051_sfr1_oc8051_tc21_n66) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u76 ( .A(oc8051_sfr1_rcap2l[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n63) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u75 ( .A(oc8051_sfr1_oc8051_tc21_n77), .Y(oc8051_sfr1_oc8051_tc21_n69) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u74 ( .A0(
        oc8051_sfr1_oc8051_tc21_n760), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[7]), .Y(
        oc8051_sfr1_oc8051_tc21_n76) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u73 ( .A0(
        oc8051_sfr1_oc8051_tc21_n62), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n63), .C0(
        oc8051_sfr1_oc8051_tc21_n76), .Y(oc8051_sfr1_oc8051_tc21_n169) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u72 ( .A(oc8051_sfr1_tl2[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n59) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u71 ( .A(oc8051_sfr1_rcap2l[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n60) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u70 ( .A0(
        oc8051_sfr1_oc8051_tc21_n750), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[6]), .Y(
        oc8051_sfr1_oc8051_tc21_n75) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u69 ( .A0(
        oc8051_sfr1_oc8051_tc21_n59), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n60), .C0(
        oc8051_sfr1_oc8051_tc21_n75), .Y(oc8051_sfr1_oc8051_tc21_n170) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u68 ( .A(oc8051_sfr1_tl2[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n56) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u67 ( .A(oc8051_sfr1_rcap2l[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n57) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u66 ( .A0(
        oc8051_sfr1_oc8051_tc21_n740), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[5]), .Y(
        oc8051_sfr1_oc8051_tc21_n74) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u65 ( .A0(
        oc8051_sfr1_oc8051_tc21_n56), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n57), .C0(
        oc8051_sfr1_oc8051_tc21_n74), .Y(oc8051_sfr1_oc8051_tc21_n171) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u64 ( .A(oc8051_sfr1_tl2[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n53) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u63 ( .A(oc8051_sfr1_rcap2l[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n54) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u62 ( .A0(
        oc8051_sfr1_oc8051_tc21_n730), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[4]), .Y(
        oc8051_sfr1_oc8051_tc21_n73) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u61 ( .A0(
        oc8051_sfr1_oc8051_tc21_n53), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n54), .C0(
        oc8051_sfr1_oc8051_tc21_n73), .Y(oc8051_sfr1_oc8051_tc21_n172) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u60 ( .A(oc8051_sfr1_tl2[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n50) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u59 ( .A(oc8051_sfr1_rcap2l[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n51) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u58 ( .A0(
        oc8051_sfr1_oc8051_tc21_n720), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[3]), .Y(
        oc8051_sfr1_oc8051_tc21_n72) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u57 ( .A0(
        oc8051_sfr1_oc8051_tc21_n50), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n51), .C0(
        oc8051_sfr1_oc8051_tc21_n72), .Y(oc8051_sfr1_oc8051_tc21_n173) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u56 ( .A(oc8051_sfr1_tl2[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n47) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u55 ( .A(oc8051_sfr1_rcap2l[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n48) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u54 ( .A0(
        oc8051_sfr1_oc8051_tc21_n710), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[2]), .Y(
        oc8051_sfr1_oc8051_tc21_n71) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u53 ( .A0(
        oc8051_sfr1_oc8051_tc21_n47), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n48), .C0(
        oc8051_sfr1_oc8051_tc21_n71), .Y(oc8051_sfr1_oc8051_tc21_n174) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u52 ( .A(oc8051_sfr1_tl2[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n44) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u51 ( .A(oc8051_sfr1_rcap2l[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n45) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u50 ( .A0(
        oc8051_sfr1_oc8051_tc21_n700), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n70) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u49 ( .A0(
        oc8051_sfr1_oc8051_tc21_n44), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n45), .C0(
        oc8051_sfr1_oc8051_tc21_n70), .Y(oc8051_sfr1_oc8051_tc21_n175) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u48 ( .A(oc8051_sfr1_tl2[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n38) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u47 ( .A(oc8051_sfr1_rcap2l[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n41) );
  AOI22_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u46 ( .A0(
        oc8051_sfr1_oc8051_tc21_n690), .A1(oc8051_sfr1_oc8051_tc21_n68), .B0(
        oc8051_sfr1_oc8051_tc21_n69), .B1(wr_dat[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n67) );
  OAI221_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u45 ( .A0(
        oc8051_sfr1_oc8051_tc21_n38), .A1(oc8051_sfr1_oc8051_tc21_n65), .B0(
        oc8051_sfr1_oc8051_tc21_n66), .B1(oc8051_sfr1_oc8051_tc21_n41), .C0(
        oc8051_sfr1_oc8051_tc21_n67), .Y(oc8051_sfr1_oc8051_tc21_n176) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u44 ( .A(
        oc8051_sfr1_oc8051_tc21_n43), .B(oc8051_sfr1_oc8051_tc21_n39), .Y(
        oc8051_sfr1_oc8051_tc21_n40) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u43 ( .A0(
        oc8051_sfr1_oc8051_tc21_n62), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n63), .C0(
        oc8051_sfr1_oc8051_tc21_n43), .C1(oc8051_sfr1_oc8051_tc21_n64), .Y(
        oc8051_sfr1_oc8051_tc21_n177) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u42 ( .A0(
        oc8051_sfr1_oc8051_tc21_n59), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n60), .C0(
        oc8051_sfr1_oc8051_tc21_n43), .C1(oc8051_sfr1_oc8051_tc21_n61), .Y(
        oc8051_sfr1_oc8051_tc21_n178) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u41 ( .A0(
        oc8051_sfr1_oc8051_tc21_n56), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n57), .C0(
        oc8051_sfr1_oc8051_tc21_n58), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n179) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u40 ( .A0(
        oc8051_sfr1_oc8051_tc21_n53), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n54), .C0(
        oc8051_sfr1_oc8051_tc21_n55), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n180) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u39 ( .A0(
        oc8051_sfr1_oc8051_tc21_n50), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n51), .C0(
        oc8051_sfr1_oc8051_tc21_n52), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n181) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u38 ( .A0(
        oc8051_sfr1_oc8051_tc21_n47), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n48), .C0(
        oc8051_sfr1_oc8051_tc21_n49), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n182) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u37 ( .A0(
        oc8051_sfr1_oc8051_tc21_n44), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n45), .C0(
        oc8051_sfr1_oc8051_tc21_n46), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n183) );
  OAI222_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u36 ( .A0(
        oc8051_sfr1_oc8051_tc21_n38), .A1(oc8051_sfr1_oc8051_tc21_n39), .B0(
        oc8051_sfr1_oc8051_tc21_n40), .B1(oc8051_sfr1_oc8051_tc21_n41), .C0(
        oc8051_sfr1_oc8051_tc21_n42), .C1(oc8051_sfr1_oc8051_tc21_n43), .Y(
        oc8051_sfr1_oc8051_tc21_n184) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u35 ( .A(
        oc8051_sfr1_oc8051_tc21_n23), .B(oc8051_sfr1_oc8051_tc21_n34), .Y(
        oc8051_sfr1_oc8051_tc21_n35) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u34 ( .A(
        oc8051_sfr1_oc8051_tc21_n35), .B(oc8051_sfr1_rclk), .Y(
        oc8051_sfr1_oc8051_tc21_n37) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u33 ( .A(wr_dat[5]), .B(
        oc8051_sfr1_oc8051_tc21_n37), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n36) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u32 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n35), .B0(
        oc8051_sfr1_oc8051_tc21_n36), .Y(oc8051_sfr1_oc8051_tc21_n185) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u31 ( .A(
        oc8051_sfr1_oc8051_tc21_n18), .B(oc8051_sfr1_oc8051_tc21_n34), .Y(
        oc8051_sfr1_oc8051_tc21_n31) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u30 ( .A(
        oc8051_sfr1_oc8051_tc21_n31), .B(oc8051_sfr1_tclk), .Y(
        oc8051_sfr1_oc8051_tc21_n33) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u29 ( .A(wr_dat[4]), .B(
        oc8051_sfr1_oc8051_tc21_n33), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n32) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u28 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n31), .B0(
        oc8051_sfr1_oc8051_tc21_n32), .Y(oc8051_sfr1_oc8051_tc21_n186) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u27 ( .A(
        oc8051_sfr1_oc8051_tc21_n27), .B(oc8051_sfr1_oc8051_tc21_n23), .Y(
        oc8051_sfr1_oc8051_tc21_n28) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u26 ( .A(
        oc8051_sfr1_oc8051_tc21_n28), .B(oc8051_sfr1_t2con_3_), .Y(
        oc8051_sfr1_oc8051_tc21_n30) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u25 ( .A(wr_dat[3]), .B(
        oc8051_sfr1_oc8051_tc21_n30), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n29) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u24 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n28), .B0(
        oc8051_sfr1_oc8051_tc21_n29), .Y(oc8051_sfr1_oc8051_tc21_n187) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u23 ( .A(
        oc8051_sfr1_oc8051_tc21_n27), .B(oc8051_sfr1_oc8051_tc21_n18), .Y(
        oc8051_sfr1_oc8051_tc21_n24) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u22 ( .A(
        oc8051_sfr1_oc8051_tc21_n24), .B(oc8051_sfr1_t2con_2_), .Y(
        oc8051_sfr1_oc8051_tc21_n26) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u21 ( .A(wr_dat[2]), .B(
        oc8051_sfr1_oc8051_tc21_n26), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n25) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u20 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n24), .B0(
        oc8051_sfr1_oc8051_tc21_n25), .Y(oc8051_sfr1_oc8051_tc21_n188) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u19 ( .A(
        oc8051_sfr1_oc8051_tc21_n23), .B(oc8051_sfr1_oc8051_tc21_n19), .Y(
        oc8051_sfr1_oc8051_tc21_n20) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u18 ( .A(
        oc8051_sfr1_oc8051_tc21_n20), .B(oc8051_sfr1_t2con_1_), .Y(
        oc8051_sfr1_oc8051_tc21_n22) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u17 ( .A(wr_dat[1]), .B(
        oc8051_sfr1_oc8051_tc21_n22), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n21) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u16 ( .A0(
        oc8051_sfr1_oc8051_tc21_n14), .A1(oc8051_sfr1_oc8051_tc21_n20), .B0(
        oc8051_sfr1_oc8051_tc21_n21), .Y(oc8051_sfr1_oc8051_tc21_n189) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u15 ( .A(
        oc8051_sfr1_oc8051_tc21_n18), .B(oc8051_sfr1_oc8051_tc21_n19), .Y(
        oc8051_sfr1_oc8051_tc21_n13) );
  AND2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u14 ( .A(
        oc8051_sfr1_oc8051_tc21_n13), .B(oc8051_sfr1_t2con_0_), .Y(
        oc8051_sfr1_oc8051_tc21_n16) );
  MXIT2_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u13 ( .A(wr_dat[0]), .B(
        oc8051_sfr1_oc8051_tc21_n16), .S0(oc8051_sfr1_oc8051_tc21_n17), .Y(
        oc8051_sfr1_oc8051_tc21_n15) );
  OAI21_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u12 ( .A0(
        oc8051_sfr1_oc8051_tc21_n13), .A1(oc8051_sfr1_oc8051_tc21_n14), .B0(
        oc8051_sfr1_oc8051_tc21_n15), .Y(oc8051_sfr1_oc8051_tc21_n190) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u11 ( .A(
        oc8051_sfr1_oc8051_tc21_tf2_set), .Y(oc8051_sfr1_oc8051_tc21_n3) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u10 ( .A0(
        oc8051_sfr1_oc8051_tc21_n10), .A1(oc8051_sfr1_oc8051_tc21_n11), .B0(
        oc8051_sfr1_oc8051_tc21_n12), .C0(oc8051_sfr1_oc8051_tc21_n850), .Y(
        oc8051_sfr1_oc8051_tc21_n4) );
  OAI211_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u9 ( .A0(
        oc8051_sfr1_oc8051_tc21_n2), .A1(oc8051_sfr1_oc8051_tc21_n3), .B0(
        oc8051_sfr1_oc8051_tc21_n4), .C0(oc8051_sfr1_oc8051_tc21_n9), .Y(
        oc8051_sfr1_oc8051_tc21_n191) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u8 ( .A(oc8051_sfr1_oc8051_tc21_n5), 
        .Y(oc8051_sfr1_t2con_6_) );
  INV_X0P5B_A12TS oc8051_sfr1_oc8051_tc21_u7 ( .A(oc8051_sfr1_oc8051_tc21_n6), 
        .Y(oc8051_sfr1_t2con_7_) );
  NAND2_X0P5A_A12TS oc8051_sfr1_oc8051_tc21_u6 ( .A(oc8051_sfr1_oc8051_tc21_n5), .B(oc8051_sfr1_oc8051_tc21_n6), .Y(oc8051_sfr1_tc2_int) );
  TIELO_X1M_A12TS oc8051_sfr1_oc8051_tc21_u5 ( .Y(oc8051_sfr1_oc8051_tc21_n1)
         );
  AND3_X0P7M_A12TS oc8051_sfr1_oc8051_tc21_u4 ( .A(wr_addr[1]), .B(wr_addr[2]), 
        .C(oc8051_sfr1_oc8051_tc21_n23), .Y(oc8051_sfr1_oc8051_tc21_n126) );
  INV_X0P5M_A12TS oc8051_sfr1_oc8051_tc21_u3 ( .A(wr_dat[1]), .Y(
        oc8051_sfr1_oc8051_tc21_n46) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n152), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n5) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n151), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n6) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n186), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n7) );
  DFFRPQN_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n185), .CK(wb_clk_i), .R(wb_rst_i), .QN(
        oc8051_sfr1_oc8051_tc21_n8) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n176), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n169), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n173), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n161), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n165), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n172), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n164), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n168), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n171), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n175), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n170), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tl2_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n174), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_tl2[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n163), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n167), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n162), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_th2_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n166), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_th2[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n190), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_0_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n189), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_1_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n187), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_3_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2con_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n188), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_t2con_2_) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tf2_set_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n191), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_tc21_tf2_set) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n153), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n154), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n155), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n156), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n157), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n158), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n159), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2h_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n160), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2h[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_brate2_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n150), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_brate2) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_1_ ( .D(
        oc8051_sfr1_oc8051_tc21_n183), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[1]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_7_ ( .D(
        oc8051_sfr1_oc8051_tc21_n177), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[7]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_6_ ( .D(
        oc8051_sfr1_oc8051_tc21_n178), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[6]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_5_ ( .D(
        oc8051_sfr1_oc8051_tc21_n179), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[5]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_4_ ( .D(
        oc8051_sfr1_oc8051_tc21_n180), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[4]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_3_ ( .D(
        oc8051_sfr1_oc8051_tc21_n181), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[3]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_2_ ( .D(
        oc8051_sfr1_oc8051_tc21_n182), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[2]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_rcap2l_reg_0_ ( .D(
        oc8051_sfr1_oc8051_tc21_n184), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_rcap2l[0]) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_tc2_event_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n220), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_tc21_tc2_event) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_neg_trans_reg ( .D(
        oc8051_sfr1_oc8051_tc21_n217), .CK(wb_clk_i), .R(wb_rst_i), .Q(
        oc8051_sfr1_oc8051_tc21_neg_trans) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2_r_reg ( .D(t2_i), .CK(wb_clk_i), 
        .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc21_t2_r) );
  DFFRPQ_X1M_A12TS oc8051_sfr1_oc8051_tc21_t2ex_r_reg ( .D(t2ex_i), .CK(
        wb_clk_i), .R(wb_rst_i), .Q(oc8051_sfr1_oc8051_tc21_t2ex_r) );
  INV_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1 ( .A(oc8051_sfr1_tl2[0]), .Y(
        oc8051_sfr1_oc8051_tc21_n690) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_1 ( .A(oc8051_sfr1_tl2[1]), 
        .B(oc8051_sfr1_tl2[0]), .CO(oc8051_sfr1_oc8051_tc21_r320_carry[2]), 
        .S(oc8051_sfr1_oc8051_tc21_n700) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_2 ( .A(oc8051_sfr1_tl2[2]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[2]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[3]), .S(
        oc8051_sfr1_oc8051_tc21_n710) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_3 ( .A(oc8051_sfr1_tl2[3]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[3]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[4]), .S(
        oc8051_sfr1_oc8051_tc21_n720) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_4 ( .A(oc8051_sfr1_tl2[4]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[4]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[5]), .S(
        oc8051_sfr1_oc8051_tc21_n730) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_5 ( .A(oc8051_sfr1_tl2[5]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[5]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[6]), .S(
        oc8051_sfr1_oc8051_tc21_n740) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_6 ( .A(oc8051_sfr1_tl2[6]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[6]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[7]), .S(
        oc8051_sfr1_oc8051_tc21_n750) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_7 ( .A(oc8051_sfr1_tl2[7]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[7]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[8]), .S(
        oc8051_sfr1_oc8051_tc21_n760) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_8 ( .A(oc8051_sfr1_th2[0]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[8]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[9]), .S(
        oc8051_sfr1_oc8051_tc21_n770) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_9 ( .A(oc8051_sfr1_th2[1]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[9]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[10]), .S(
        oc8051_sfr1_oc8051_tc21_n780) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_10 ( .A(oc8051_sfr1_th2[2]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[10]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[11]), .S(
        oc8051_sfr1_oc8051_tc21_n790) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_11 ( .A(oc8051_sfr1_th2[3]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[11]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[12]), .S(
        oc8051_sfr1_oc8051_tc21_n800) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_12 ( .A(oc8051_sfr1_th2[4]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[12]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[13]), .S(
        oc8051_sfr1_oc8051_tc21_n810) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_13 ( .A(oc8051_sfr1_th2[5]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[13]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[14]), .S(
        oc8051_sfr1_oc8051_tc21_n820) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_14 ( .A(oc8051_sfr1_th2[6]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[14]), .CO(
        oc8051_sfr1_oc8051_tc21_r320_carry[15]), .S(
        oc8051_sfr1_oc8051_tc21_n830) );
  ADDH_X1M_A12TS oc8051_sfr1_oc8051_tc21_r320_u1_1_15 ( .A(oc8051_sfr1_th2[7]), 
        .B(oc8051_sfr1_oc8051_tc21_r320_carry[15]), .CO(
        oc8051_sfr1_oc8051_tc21_n850), .S(oc8051_sfr1_oc8051_tc21_n840) );
endmodule

