

module oc8051_top ( wb_rst_i, wb_clk_i, wbi_adr_o, wbi_dat_i, wbi_stb_o, 
                    wbi_ack_i, wbi_cyc_o, wbi_err_i, wbd_dat_i, wbd_dat_o, 
                    wbd_adr_o, wbd_we_o, wbd_ack_i, wbd_stb_o, wbd_cyc_o, 
                    wbd_err_i, int0_i, int1_i, p0_i, p0_o, p1_i, p1_o, p2_i, 
                    p2_o, p3_i, p3_o, rxd_i, txd_o, t0_i, t1_i, t2_i, t2ex_i, 
                    ea_in ) ;

    input wb_rst_i ;
    input wb_clk_i ;
    output [15:0]wbi_adr_o ;
    input [31:0]wbi_dat_i ;
    output wbi_stb_o ;
    input wbi_ack_i ;
    output wbi_cyc_o ;
    input wbi_err_i ;
    input [7:0]wbd_dat_i ;
    output [7:0]wbd_dat_o ;
    output [15:0]wbd_adr_o ;
    output wbd_we_o ;
    input wbd_ack_i ;
    output wbd_stb_o ;
    output wbd_cyc_o ;
    input wbd_err_i ;
    input int0_i ;
    input int1_i ;
    input [7:0]p0_i ;
    output [7:0]p0_o ;
    input [7:0]p1_i ;
    output [7:0]p1_o ;
    input [7:0]p2_i ;
    output [7:0]p2_o ;
    input [7:0]p3_i ;
    output [7:0]p3_o ;
    input rxd_i ;
    output txd_o ;
    input t0_i ;
    input t1_i ;
    input t2_i ;
    input t2ex_i ;
    input ea_in ;

    wire sub_result_7, sub_result_6, sub_result_5, sub_result_4, sub_result_3, 
         sub_result_2, sub_result_1, sub_result_0, wait_data, bit_out, bit_data, 
         bit_addr, op1_cur_2, op1_cur_1, op1_cur_0, comp_wait, wr_ind, cy, srcAc, 
         eq, comp_sel_1, comp_sel_0, op3_n_7, op3_n_6, op3_n_5, op3_n_4, op3_n_3, 
         op3_n_2, op3_n_1, op3_n_0, op2_n_7, op2_n_6, op2_n_5, op2_n_4, op2_n_3, 
         op2_n_2, op2_n_1, op2_n_0, op1_n_7, op1_n_6, op1_n_5, op1_n_4, op1_n_3, 
         op1_n_2, op1_n_1, op1_n_0, pc_wr_sel_2, pc_wr_sel_1, pc_wr_sel_0, pc_wr, 
         rd, wr, alu_cy, desOv, desAc, desCy, des2_7, des2_6, des2_5, des2_4, 
         des2_3, des2_2, des2_1, des2_0, des1_7, des1_6, des1_5, des1_4, des1_3, 
         des1_2, des1_1, des1_0, des_acc_7, des_acc_6, des_acc_5, des_acc_4, 
         des_acc_3, des_acc_2, des_acc_1, des_acc_0, src3_7, src3_6, src3_5, 
         src3_4, src3_3, src3_2, src3_1, src3_0, src2_7, src2_6, src2_5, src2_4, 
         src2_3, src2_2, src2_1, src2_0, src1_7, src1_6, src1_5, src1_4, src1_3, 
         src1_2, src1_1, src1_0, psw_set_1, psw_set_0, alu_op_3, alu_op_2, 
         alu_op_1, alu_op_0, mem_act_2, mem_act_1, mem_act_0, mem_wait, 
         int_src_7, int_src_5, int_src_4, int_src_3, int_src_1, int_ack, intr, 
         reti, rmw, bank_sel_1, bank_sel_0, cy_sel_1, cy_sel_0, sfr_bit, 
         rd_addr_7, rd_addr_6, rd_addr_5, rd_addr_4, rd_addr_3, rd_addr_2, 
         rd_addr_1, rd_addr_0, wr_addr_7, wr_addr_6, wr_addr_5, wr_addr_4, 
         wr_addr_3, wr_addr_2, wr_addr_1, wr_addr_0, sfr_out_7, sfr_out_6, 
         sfr_out_5, sfr_out_4, sfr_out_3, sfr_out_2, sfr_out_1, sfr_out_0, 
         ram_out_7, ram_out_6, ram_out_5, ram_out_4, ram_out_3, ram_out_2, 
         ram_out_1, ram_out_0, ram_data_7, ram_data_6, ram_data_5, ram_data_4, 
         ram_data_3, ram_data_2, ram_data_1, ram_data_0, src_sel1_2, src_sel1_1, 
         src_sel1_0, ram_wr_sel_2, ram_wr_sel_1, ram_wr_sel_0, ram_rd_sel_2, 
         ram_rd_sel_1, ram_rd_sel_0, src_sel2_1, src_sel2_0, wr_sfr_1, wr_sfr_0, 
         src_sel3, pc_15, pc_14, pc_13, pc_12, pc_11, pc_10, pc_9, pc_8, pc_7, 
         pc_6, pc_5, pc_4, pc_3, pc_2, pc_1, pc_0, sp_w_7, sp_w_6, sp_w_5, 
         sp_w_4, sp_w_3, sp_w_2, sp_w_1, sp_w_0, sp_7, sp_6, sp_5, sp_4, sp_3, 
         sp_2, sp_1, sp_0, acc_7, acc_6, acc_5, acc_4, acc_3, acc_2, acc_1, 
         acc_0, ri_7, ri_6, ri_5, ri_4, ri_3, ri_2, ri_1, ri_0, dptr_lo_7, 
         dptr_lo_6, dptr_lo_5, dptr_lo_4, dptr_lo_3, dptr_lo_2, dptr_lo_1, 
         dptr_lo_0, dptr_hi_7, dptr_hi_6, dptr_hi_5, dptr_hi_4, dptr_hi_3, 
         dptr_hi_2, dptr_hi_1, dptr_hi_0, wr_dup_1054, pc_wr_dup_1371, we, 
         ea_int, nx747, nx749, state_0, nx4, state_1, nx10, nx24, nx48, nx64, 
         nx78, nx82, nx84, op_2, nx98, nx102, nx110, op_3, nx124, nx126, op_1, 
         op_0, nx148, nx150, op_4, nx160, op_5, nx170, nx174, op_6, nx184, op_7, 
         nx194, nx196, nx198, nx200, nx206, nx216, nx224, nx234, nx242, nx250, 
         nx254, nx262, nx264, nx266, nx272, nx274, nx276, nx282, nx288, nx290, 
         nx304, nx306, nx308, nx318, nx328, nx330, nx332, nx346, nx352, nx364, 
         nx368, nx376, nx380, nx396, nx398, nx400, nx406, nx420, nx424, nx430, 
         nx434, nx442, nx450, nx460, nx462, nx472, nx484, nx488, nx492, nx494, 
         nx506, nx508, nx516, nx530, nx532, nx544, nx554, nx564, nx570, nx582, 
         nx588, nx608, nx656, nx658, nx674, nx734, wr_dup_832, nx756, nx760, 
         nx780, nx784, nx792, nx794, nx796, nx804, nx806, nx810, nx820, nx834, 
         nx844, nx850, nx860, nx870, nx878, ram_wr_sel_0__dup_833, nx904, nx914, 
         nx930, nx946, nx948, nx952, nx968, nx1002, nx1006, nx1012, nx1020, 
         nx1046, ram_wr_sel_1__dup_834, nx1066, nx1068, nx1076, nx1080, nx1084, 
         nx1128, nx1136, ram_wr_sel_2__dup_835, wr_sfr_0__dup_836, nx1168, 
         nx1178, nx1188, nx1196, nx1214, nx1228, nx1240, nx1242, nx1252, nx1254, 
         nx1256, nx1272, nx1282, wr_sfr_1__dup_837, nx1292, nx1302, nx1312, 
         nx1324, alu_op_0__dup_838, nx1356, nx1372, nx1388, nx1396, nx1408, 
         alu_op_1__dup_839, nx1444, nx1454, nx1466, nx1472, nx1484, 
         alu_op_2__dup_840, nx1510, nx1526, nx1540, nx1556, alu_op_3__dup_841, 
         nx1568, nx1596, nx1620, nx1660, nx1672, nx1684, nx1712, nx1730, nx1742, 
         nx1748, nx1762, nx1766, nx1780, nx1802, nx1816, nx1820, nx1842, nx1850, 
         nx1872, nx1898, nx1920, nx1932, nx1952, nx1972, nx2002, nx2010, nx2036, 
         nx2042, nx2046, nx2054, nx2084, nx2098, nx2120, nx2148, nx2172, nx2188, 
         nx2192, nx2204, nx2250, nx2272, nx2292, nx2304, nx2322, nx2336, nx2342, 
         nx2360, nx2388, nx2394, nx2414, nx2426, ram_rd_sel_r_0, nx2452, nx2462, 
         nx2484, nx2500, ram_rd_sel_r_1, nx2532, ram_rd_sel_r_2, nx3887, nx3897, 
         NOT_nx10, nx3987, nx4007, nx4017, nx4037, nx4047, nx4057, nx4077, 
         nx4097, nx4117, nx4127, nx4137, nx4147, nx4157, nx4177, nx4188, nx4193, 
         nx4198, nx4202, nx4204, nx4207, nx4210, nx4212, nx4214, nx4216, nx4221, 
         nx4226, nx4230, nx4240, nx4246, nx4255, nx4257, nx4259, nx4267, nx4271, 
         nx4273, nx4275, nx4278, nx4281, nx4283, nx4285, nx4288, nx4294, nx4297, 
         nx4299, nx4302, nx4306, nx4308, nx4310, nx4317, nx4322, nx4325, nx4332, 
         nx4334, nx4338, nx4340, nx4344, nx4346, nx4348, nx4350, nx4354, nx4356, 
         nx4361, nx4364, nx4372, nx4377, nx4382, nx4390, nx4395, nx4398, nx4400, 
         nx4402, nx4404, nx4415, nx4420, nx4422, nx4424, nx4429, nx4432, nx4434, 
         nx4436, nx4439, nx4444, nx4446, nx4448, nx4451, nx4456, nx4460, nx4466, 
         nx4468, nx4471, nx4476, nx4478, nx4482, nx4486, nx4488, nx4490, nx4492, 
         nx4495, nx4498, nx4503, nx4507, nx4511, nx4514, nx4516, nx4519, nx4524, 
         nx4526, nx4533, nx4536, nx4538, nx4544, nx4546, nx4550, nx4553, nx4556, 
         nx4560, nx4563, nx4567, nx4569, nx4571, nx4574, nx4576, nx4578, nx4582, 
         nx4588, nx4590, nx4592, nx4597, nx4600, nx4602, nx4604, nx4606, nx4608, 
         nx4610, nx4614, nx4617, nx4621, nx4626, nx4628, nx4630, nx4633, nx4637, 
         nx4642, nx4649, nx4653, nx4657, nx4662, nx4664, nx4667, nx4670, nx4673, 
         nx4675, nx4683, nx4685, nx4688, nx4692, nx4694, nx4696, nx4699, nx4704, 
         nx4707, nx4710, nx4712, nx4714, nx4721, nx4723, nx4726, nx4737, nx4741, 
         nx4743, nx4745, nx4749, nx4755, nx4761, nx4766, nx4771, nx4773, nx4777, 
         nx4779, nx4785, nx4791, nx4794, nx4798, nx4800, nx4802, nx4805, nx4807, 
         nx4812, nx4817, nx4819, nx4823, nx4825, nx4827, nx4830, nx4832, nx4834, 
         nx4838, nx4844, nx4847, nx4849, nx4853, nx4858, nx4865, nx4869, nx4872, 
         nx4875, nx4883, nx4887, nx4889, nx4896, nx4899, nx4901, nx4905, nx4907, 
         nx4910, nx4914, nx4916, nx4918, nx4921, nx4924, nx4933, nx4935, nx4937, 
         nx4941, nx4944, nx4947, nx4956, nx4959, nx4961, nx4969, nx4973, nx4977, 
         nx4981, nx4983, nx4987, nx4989, nx4994, nx4998, nx5001, nx5003, nx5006, 
         nx5009, nx5012, nx5016, nx5018, nx5023, nx5027, nx5029, nx5033, divOv, 
         divsrc2_7, divsrc2_6, divsrc2_5, divsrc2_4, divsrc2_3, divsrc2_2, 
         divsrc2_1, divsrc2_0, divsrc1_7, divsrc1_6, divsrc1_5, divsrc1_4, 
         divsrc1_3, divsrc1_2, divsrc1_1, divsrc1_0, mulOv, mulsrc2_7, mulsrc2_6, 
         mulsrc2_5, mulsrc2_4, mulsrc2_3, mulsrc2_2, mulsrc2_1, mulsrc2_0, 
         mulsrc1_7, mulsrc1_6, mulsrc1_5, mulsrc1_4, mulsrc1_3, mulsrc1_2, 
         mulsrc1_1, mulsrc1_0, enable_mul, enable_div, nx2, nx6, nx969, nx12, 
         nx18, nx22, nx40, nx44, nx50, nx56, nx60, nx970, nx76, nx80, nx94, 
         nx971, nx972, nx114, nx128, nx136, nx162, nx168, nx182, nx188, nx973, 
         nx974, nx975, nx222, nx240, nx244, nx252, nx258, nx976, nx278, nx977, 
         nx298, nx978, nx326, nx979, nx980, nx338, nx350, nx981, nx358, nx982, 
         nx370, nx983, nx984, nx410, nx414, nx440, nx985, nx454, nx458, nx986, 
         nx502, nx987, nx514, nx520, nx536, nx550, nx988, nx989, nx580, nx610, 
         nx622, nx642, nx648, nx990, nx662, nx664, nx680, nx684, nx694, nx710, 
         nx714, nx744, nx750, nx991, nx762, nx768, nx776, nx992, nx786, nx993, 
         nx814, nx836, nx868, nx994, nx876, nx882, nx888, nx900, nx910, nx916, 
         nx936, nx995, nx996, nx997, nx1028, nx1032, nx1048, nx1052, nx1104, 
         nx1118, nx1140, nx1152, nx1172, nx1176, nx1184, nx1208, nx1212, nx1224, 
         nx998, nx1258, nx1270, nx1300, nx1304, nx1316, nx1346, nx1350, nx1362, 
         nx1386, nx1398, nx1402, nx1414, nx999, nx1448, nx1490, nx1494, nx1520, 
         nx1534, nx1546, nx1000, nx1598, nx1614, nx1618, nx1630, nx1658, nx1495, 
         nx1501, nx1505, nx1509, nx1511, nx1513, nx1519, nx1521, nx1523, nx1533, 
         nx1537, nx1539, nx1541, nx1543, nx1547, nx1557, nx1559, nx1561, nx1563, 
         nx1565, nx1569, nx1579, nx1581, nx1583, nx1585, nx1591, nx1593, nx1595, 
         nx1603, nx1605, nx1607, nx1611, nx1615, nx1623, nx1625, nx1627, nx1629, 
         nx1633, nx1637, nx1639, nx1641, nx1643, nx1645, nx1651, nx1653, nx1657, 
         nx1661, nx1663, nx1668, nx1671, nx1674, nx1676, nx1679, nx1681, nx1685, 
         nx1687, nx1689, nx1693, nx1696, nx1698, nx1700, nx1706, nx1711, nx1714, 
         nx1718, nx1722, nx1724, nx1727, nx1001, nx1733, nx1736, nx1739, nx1743, 
         nx1746, nx1750, nx1754, nx1757, nx1760, nx1763, nx1765, nx1768, nx1770, 
         nx1773, nx1776, nx1778, nx1003, nx1782, nx1787, nx1790, nx1793, nx1795, 
         nx1798, nx1800, nx1803, nx1808, nx1811, nx1815, nx1819, nx1824, nx1826, 
         nx1828, nx1831, nx1835, nx1837, nx1839, nx1004, nx1847, nx1849, nx1854, 
         nx1859, nx1862, nx1866, nx1868, nx1870, nx1873, nx1877, nx1880, nx1882, 
         nx1887, nx1890, nx1894, nx1896, nx1005, nx1901, nx1903, nx1906, nx1911, 
         nx1914, nx1917, nx1007, nx1922, nx1924, nx1926, nx1931, nx1933, nx1935, 
         nx1938, nx1940, nx1943, nx1945, nx1947, nx1950, nx1958, nx1963, nx1968, 
         nx1970, nx1974, nx1976, nx1978, nx1981, nx1983, nx1986, nx1988, nx1991, 
         nx1994, nx1997, nx2000, nx1008, nx2004, nx2006, nx2013, nx2016, nx2019, 
         nx2021, nx2023, nx2026, nx2028, nx2031, nx2033, nx2035, nx2038, nx2040, 
         nx2043, nx2045, nx2048, nx2051, nx1009, nx2059, nx2061, nx2063, nx2066, 
         nx2068, nx2071, nx2074, nx2077, nx2079, nx2081, nx2083, nx2086, nx2089, 
         nx2092, nx2097, nx2099, nx2101, nx2103, nx2108, nx2111, nx2114, nx2119, 
         nx2121, nx2123, nx2125, nx2130, nx2133, nx2137, nx2140, nx2142, nx2144, 
         nx2146, nx2151, nx2154, nx2157, nx2162, nx2164, nx2166, nx2168, nx2173, 
         nx2176, nx2179, nx2184, nx2186, nx1010, nx2190, nx2195, nx2198, nx2202, 
         nx2207, nx2209, rd_data_m_7, rd_data_m_6, rd_data_m_5, rd_data_m_4, 
         rd_data_m_3, rd_data_m_2, rd_data_m_1, rd_data_m_0, wr_addr_m_5, 
         wr_addr_m_3, wr_addr_m_2, wr_addr_m_1, wr_addr_m_0, rd_addr_m_5, 
         rd_addr_m_3, rd_addr_m_2, rd_addr_m_1, rd_addr_m_0, wr_data_m_7, 
         wr_data_m_6, wr_data_m_5, wr_data_m_4, wr_data_m_3, wr_data_m_2, 
         wr_data_m_1, wr_data_m_0, NOT_rd_en, rd_addr_m_6, rd_addr_m_4, 
         wr_addr_m_6, wr_addr_m_4, bit_addr_r, nx20, bit_select_0, rd_en_r, nx88, 
         nx106, nx1055, nx142, nx144, nx1056, nx154, wr_data_r_6, bit_select_2, 
         bit_select_1, nx1057, nx192, wr_data_r_4, nx226, wr_data_r_2, nx1058, 
         wr_data_r_0, nx302, wr_data_r_7, wr_data_r_5, wr_data_r_3, wr_data_r_1, 
         nx339, nx341, nx351, nx353, nx363, nx365, nx367, nx371, nx373, nx375, 
         nx379, nx383, nx387, nx391, nx395, nx397, nx401, nx403, nx409, nx423, 
         nx427, nx447, nx451, nx453, nx455, nx1059, nx467, nx471, nx475, nx481, 
         nx487, nx491, nx1060, nx498, nx1061, nx1062, nx509, nx513, nx531, nx533, 
         nx535, nx537, nx539, nx541, nx543, nx545, nx547, nx1144, nx1145, 
         op2_r_0, nx1146, op2_r_1, op2_r_2, op2_r_3, op2_r_4, op2_r_5, op2_r_6, 
         op2_r_7, op3_r_0, nx134, op1_r_0, nx1147, nx1148, nx1149, nx176, nx1150, 
         nx1151, op3_r_1, op1_r_1, op3_r_2, op1_r_2, op3_r_3, op1_r_3, op3_r_4, 
         op1_r_4, op3_r_5, op1_r_5, op3_r_6, op1_r_6, op3_r_7, op1_r_7, nx526, 
         nx1153, nx1154, nx1155, nx1156, nx551, nx555, nx559, nx563, nx567, 
         nx1157, nx572, nx575, nx578, nx585, nx587, nx589, nx594, nx596, nx598, 
         nx603, nx605, nx607, nx612, nx614, nx616, nx621, nx623, nx625, nx630, 
         nx632, nx634, nx639, nx641, nx643, nx8, nx14, nx1175, nx28, nx1177, 
         nx46, nx54, nx1179, nx74, nx111, nx1180, nx119, nx125, nx43, buff_3__0, 
         wr_bit_r, nx1234, nx1235, nx66, buff_2__0, nx86, buff_1__0, nx1236, 
         buff_7__0, nx118, nx130, buff_0__0, nx152, buff_6__0, nx1237, buff_5__0, 
         nx190, buff_4__0, nx212, buff_3__1, buff_2__1, buff_1__1, buff_7__1, 
         buff_0__1, buff_6__1, buff_5__1, buff_4__1, buff_3__2, buff_2__2, 
         buff_1__2, buff_7__2, buff_0__2, buff_6__2, buff_5__2, buff_4__2, 
         buff_3__3, buff_2__3, buff_1__3, buff_7__3, buff_0__3, buff_6__3, 
         buff_5__3, buff_4__3, buff_3__4, buff_2__4, buff_1__4, buff_7__4, 
         buff_0__4, buff_6__4, buff_5__4, buff_4__4, buff_3__5, buff_2__5, 
         buff_1__5, buff_7__5, buff_0__5, buff_6__5, buff_5__5, buff_4__5, 
         buff_3__6, buff_2__6, buff_1__6, buff_7__6, buff_0__6, buff_6__6, 
         buff_5__6, buff_4__6, buff_3__7, buff_2__7, buff_1__7, buff_7__7, 
         buff_0__7, buff_6__7, buff_5__7, buff_4__7, NOT_nx14, NOT_nx74, 
         NOT_nx94, NOT_nx122, NOT_nx140, NOT_nx164, NOT_nx182, NOT_nx202, nx1992, 
         nx1995, nx1238, nx2001, nx2003, nx2005, nx1239, nx2015, nx2017, nx2020, 
         nx2024, nx1241, nx2032, nx1243, nx1244, nx1245, nx1246, nx2069, nx2073, 
         nx1247, nx1248, nx1249, nx2090, nx2094, nx2100, nx1250, nx2107, nx1251, 
         nx2117, nx1253, nx2124, nx2128, nx2134, nx1255, nx2141, nx2145, nx1257, 
         nx1259, nx2158, nx1260, nx1261, nx2171, nx2175, nx1262, rd_ind, nx1465, 
         nx1467, nx1468, op2_buff_0, idat_old_16, nx1469, nx26, pc_wr_r2, 
         pc_wr_r, nx36, op_pos_2, nx5672, nx1470, op_pos_0, ddat_ir_7, dack_ir, 
         idat_old_15, idat_cur_15, op_pos_1, ddat_ir_3, idat_old_11, idat_cur_11, 
         nx5675, idat_cur_3, nx120, int_ack_t, nx1471, nx1473, nx138, nx1474, 
         idat_old_3, nx164, nx1475, idat_old_19, idat_cur_19, idat_old_27, 
         idat_cur_27, nx1476, nx1477, cdone, istb_t, imem_wait, nx260, cdata_3, 
         nx270, ddat_ir_1, idat_cur_9, idat_old_17, idat_cur_17, idat_old_25, 
         idat_cur_25, idat_old_9, idat_old_1, idat_cur_1, nx378, nx388, nx392, 
         nx1478, cdata_1, nx416, ddat_ir_5, idat_old_13, idat_cur_13, idat_cur_5, 
         nx1479, nx466, idat_old_5, idat_old_21, idat_cur_21, idat_old_29, 
         idat_cur_29, nx518, nx1480, cdata_5, ddat_ir_0, idat_old_8, idat_cur_8, 
         idat_cur_0, nx576, nx1481, idat_old_0, idat_old_24, idat_cur_24, nx618, 
         cdata_0, nx1482, ddat_ir_4, idat_cur_12, idat_old_20, idat_cur_20, 
         idat_old_28, idat_cur_28, idat_old_12, idat_old_4, idat_cur_4, nx1483, 
         nx754, nx1485, cdata_4, nx778, ddat_ir_6, idat_old_14, idat_cur_14, 
         idat_cur_6, nx822, nx828, idat_old_6, idat_old_22, idat_cur_22, 
         idat_old_30, idat_cur_30, nx880, cdata_6, ddat_ir_2, idat_old_10, 
         idat_cur_10, idat_cur_2, nx1486, nx1487, idat_old_2, idat_old_18, 
         idat_cur_18, idat_old_26, idat_cur_26, nx1488, nx1489, cdata_2, nx1491, 
         nx1038, nx1042, nx5677, nx1492, nx1070, idat_cur_7, nx1108, nx1114, 
         idat_old_7, idat_old_23, idat_cur_23, idat_old_31, idat_cur_31, nx1166, 
         nx1493, cdata_7, nx1496, nx1497, nx1498, nx1499, nx1276, nx1500, nx1306, 
         nx1318, nx1340, nx1352, nx1354, idat_cur_16, nx1502, nx1404, nx1503, 
         nx1420, nx1428, NOT_rd, nx1504, nx1456, op2_buff_2, nx1506, op2_buff_3, 
         nx1538, imm2_r_0, op3_buff_0, int_vec_buff_0, nx1580, nx1507, nx1602, 
         ri_r_0, nx1616, nx1624, imm_r_0, nx1638, rn_r_0, nx1654, imm2_r_1, 
         op3_buff_1, int_vec_buff_1, nx1682, ri_r_1, imm_r_1, op2_buff_1, nx1734, 
         rn_r_1, imm2_r_2, op3_buff_2, int_vec_buff_2, nx1784, ri_r_2, imm_r_2, 
         rn_r_2, imm2_r_3, op3_buff_3, int_vec_buff_3, nx1852, ri_r_3, imm_r_3, 
         rn_r_3, nx1900, imm2_r_4, op3_buff_4, int_vec_buff_4, nx1508, ri_r_4, 
         imm_r_4, op2_buff_4, nx1512, rn_r_4, ri_r_5, imm_r_5, op2_buff_5, 
         nx1514, nx2056, imm2_r_5, op3_buff_5, int_vec_buff_5, nx2088, ri_r_6, 
         imm_r_6, op2_buff_6, nx1515, imm2_r_6, op3_buff_6, int_vec_buff_6, 
         nx1516, imm_r_7, op2_buff_7, nx2232, ri_r_7, imm2_r_7, op3_buff_7, 
         int_vec_buff_7, nx2282, nx2324, nx2332, nx1517, nx2356, nx1518, 
         pc_buf_0, nx2430, nx2438, nx2446, nx2454, nx2464, nx2478, nx2488, 
         nx2504, nx2512, pc_buf_1, nx2558, NOT_nx2554, nx2562, nx2572, nx2588, 
         nx2604, nx2612, pc_buf_2, nx2638, nx2648, nx2658, nx2662, nx2674, 
         pc_buf_3, nx2686, nx2696, nx2710, nx2722, nx2730, nx2746, nx2754, 
         nx2770, pc_buf_4, nx2818, nx2826, nx2838, nx2850, nx2858, pc_buf_5, 
         nx2874, nx2884, nx2892, nx2898, nx2904, nx2916, nx2932, nx2938, nx2954, 
         pc_buf_6, nx3002, nx3010, nx3016, nx3022, nx3034, nx3042, pc_buf_7, 
         nx3058, nx3068, nx3076, nx3082, nx3088, nx3100, nx3116, nx3122, nx3138, 
         pc_buf_8, nx3146, nx3156, nx3158, nx3168, NOT_nx2552, nx3184, nx3206, 
         NOT_nx2430, nx3222, nx3228, nx3234, nx3246, nx3254, pc_buf_9, nx3266, 
         nx3274, nx3296, nx3302, nx3308, nx3324, nx3338, nx3344, nx3360, 
         pc_buf_10, nx3368, nx3376, nx3410, nx3426, nx3432, nx3438, nx3450, 
         nx3458, pc_buf_11, nx3472, nx3476, nx3484, nx3486, nx3496, nx3502, 
         nx3508, nx3528, nx3542, nx3548, nx3564, pc_buf_12, nx3574, nx3582, 
         nx3610, nx3624, nx3630, nx3636, nx3648, nx3656, pc_buf_13, nx3670, 
         nx3678, nx3688, nx3694, nx3700, nx3720, nx3734, nx3740, nx3756, 
         pc_buf_14, nx3802, nx3816, nx3822, nx3828, nx3840, nx3848, pc_buf_15, 
         nx3872, nx3882, nx3886, nx3894, nx3908, int_ack_buff, nx3924, nx3944, 
         nx3968, NOT_dack_i, nx3976, nx4036, nx4048, nx4060, nx4072, nx4084, 
         nx4096, nx4108, nx4120, iadr_t_0, iadr_t_1, iadr_t_2, iadr_t_3, 
         iadr_t_4, iadr_t_5, iadr_t_6, iadr_t_7, iadr_t_8, iadr_t_9, iadr_t_10, 
         iadr_t_11, iadr_t_12, iadr_t_13, iadr_t_14, iadr_t_15, rd_addr_r, 
         NOT_nx5673, nx5694, nx5724, nx5744, nx5754, nx5774, nx5794, nx5814, 
         nx5824, nx5834, nx5854, nx5864, nx5884, nx5914, nx5934, nx5954, nx5974, 
         nx5994, nx6014, nx6034, nx6054, nx6074, nx6094, nx6114, nx6134, nx6144, 
         nx6164, nx6194, nx6214, nx6234, nx6254, nx6274, nx6294, nx6314, nx6334, 
         nx6354, nx6374, nx6394, nx6414, nx6424, nx6434, nx6454, nx6474, nx6494, 
         nx6504, nx6514, nx6524, NOT_intr, NOT_nx2426, nx6794, nx6814, nx6824, 
         nx6874, nx6884, nx6914, nx6924, nx6954, nx6994, nx7034, nx7074, nx7094, 
         nx7104, nx7114, nx7124, nx7134, nx7144, nx7154, nx7164, nx7174, nx7264, 
         nx7274, nx7284, nx7294, nx7304, nx7314, nx7324, nx7334, NOT_nx226, 
         nx7505, nx7512, nx7515, nx7519, nx7521, nx7526, nx7533, nx7537, nx7539, 
         nx7541, nx7545, nx7553, nx7555, nx7559, nx7566, nx7568, nx7570, nx7572, 
         nx7575, nx7581, nx7586, nx7588, nx7591, nx7593, nx7595, nx7600, nx7603, 
         nx7607, nx7610, nx7613, nx7617, nx7621, nx7623, nx7625, nx7628, nx7633, 
         nx7635, nx7638, nx7643, nx7645, nx7650, nx7652, nx7654, nx7656, nx7661, 
         nx7663, nx7665, nx7668, nx7670, nx7674, nx7679, nx7683, nx7685, nx7687, 
         nx7699, nx7704, nx7708, nx7710, nx7714, nx7719, nx7721, nx7726, nx7728, 
         nx7730, nx7735, nx7742, nx7744, nx7747, nx7749, nx7751, nx7761, nx7763, 
         nx7766, nx7770, nx7774, nx7776, nx7778, nx7780, nx7785, nx7788, nx7793, 
         nx7795, nx7800, nx7802, nx7804, nx7808, nx7812, nx7814, nx7818, nx7823, 
         nx7825, nx7830, nx7832, nx7834, nx7839, nx7846, nx7848, nx7851, nx7853, 
         nx7856, nx7860, nx7862, nx7864, nx7867, nx7872, nx7874, nx7877, nx7882, 
         nx7884, nx7889, nx7891, nx7893, nx7898, nx7901, nx7903, nx7905, nx7908, 
         nx7912, nx7914, nx7916, nx7919, nx7924, nx7926, nx7929, nx7934, nx7936, 
         nx7941, nx7943, nx7945, nx7950, nx7953, nx7955, nx7958, nx7965, nx7975, 
         nx7981, nx7984, nx7989, nx7991, nx7996, nx7998, nx8000, nx8005, nx8010, 
         nx8012, nx8014, nx8017, nx8019, nx8022, nx8025, nx8028, nx8031, nx8035, 
         nx8037, nx8040, nx8043, nx8046, nx8049, nx8056, nx8059, nx8062, nx8067, 
         nx8069, nx8071, nx8073, nx8075, nx8079, nx8081, nx8083, nx8086, nx8091, 
         nx8093, nx8098, nx8100, nx8102, nx8106, nx8108, nx8119, nx8123, nx8127, 
         nx8131, nx8135, nx8139, nx8143, nx8147, nx8155, nx8161, nx8167, nx8173, 
         nx8179, nx8183, nx8185, nx8189, nx8191, nx8197, nx8201, nx8205, nx8209, 
         nx8213, nx8217, nx8221, nx8225, nx8229, nx8235, nx8239, nx8246, nx8253, 
         nx8256, nx8260, nx8264, nx8268, nx8270, nx8273, nx8277, nx8283, nx8285, 
         nx8288, nx8292, nx8298, nx8300, nx8303, nx8307, nx8311, nx8315, nx8317, 
         nx8320, nx8324, nx8330, nx8332, nx8335, nx8339, nx8345, nx8347, nx8350, 
         nx8354, nx8360, nx8362, nx8365, nx8369, nx8371, nx8374, nx8378, nx8381, 
         nx8385, nx8387, nx8389, nx8392, nx8396, nx8398, nx8400, nx8403, nx8407, 
         nx8409, nx8411, nx8414, nx8418, nx8420, nx8422, nx8425, nx8429, nx8431, 
         nx8433, nx8436, nx8440, nx8442, nx8444, nx8447, nx8451, nx8453, nx8455, 
         nx8458, nx8462, nx8466, nx8468, nx8472, nx8474, nx8478, nx8481, nx8483, 
         nx8489, nx8494, nx8498, nx8502, nx8504, nx8506, nx8508, nx8512, nx8515, 
         nx8517, nx8519, nx8521, nx8523, nx8525, nx8528, nx8533, nx8537, nx8541, 
         nx8544, nx8546, nx8549, nx8551, nx8560, nx8562, nx8564, nx8567, nx8570, 
         nx8574, nx8578, nx8581, nx8583, nx8585, nx8592, nx8595, nx8599, nx8601, 
         nx8604, nx8606, nx8610, nx8613, nx8620, nx8622, nx8624, nx8626, nx8628, 
         nx8634, nx8637, nx8641, nx8643, nx8645, nx8648, nx8652, nx8655, nx8659, 
         nx8661, nx8664, nx8666, nx8669, nx8672, nx8676, nx8678, nx8681, nx8684, 
         nx8686, nx8689, nx8691, nx8695, nx8698, nx8700, nx8703, nx8705, nx8710, 
         nx8717, nx8720, nx8724, nx8726, nx8728, nx8731, nx8735, nx8738, nx8742, 
         nx8745, nx8747, nx8749, nx8752, nx8756, nx8758, nx8761, nx8764, nx8766, 
         nx8769, nx8771, nx8775, nx8778, nx8780, nx8783, nx8787, nx8794, nx8797, 
         nx8801, nx8803, nx8806, nx8811, nx8813, nx8815, nx8819, nx8822, nx8826, 
         nx8830, nx8832, nx8835, nx8839, nx8842, nx8854, nx8856, nx8860, nx8863, 
         nx8865, nx8868, nx8871, nx8873, nx8875, nx8879, nx8886, nx8889, nx8893, 
         nx8895, nx8897, nx8901, nx8904, nx8908, nx8912, nx8914, nx8917, nx8919, 
         nx8921, nx8923, nx8926, nx8930, nx8932, nx8935, nx8937, nx8941, nx8943, 
         nx8946, nx8948, nx8951, nx8954, nx8956, nx8959, nx8966, nx8973, nx8976, 
         nx8980, nx8982, nx8986, nx8989, nx8993, nx8997, nx9000, nx9003, nx9005, 
         nx9007, nx9009, nx9012, nx9016, nx9018, nx9021, nx9025, nx9027, nx9030, 
         nx9032, nx9035, nx9038, nx9040, nx9043, nx9047, nx9054, nx9057, nx9061, 
         nx9063, nx9067, nx9070, nx9076, nx9078, nx9081, nx9083, nx9085, nx9087, 
         nx9090, nx9094, nx9099, nx9102, nx9104, nx9106, nx9109, nx9112, nx9116, 
         nx9120, nx9124, nx9127, nx9129, nx9141, nx9147, nx9149, nx9154, nx9159, 
         nx9163, nx9168, nx9172, nx9177, nx9181, nx9186, nx9190, nx9193, nx9199, 
         nx9202, nx9205, nx9207, nx9210, nx9215, nx9218, nx9221, nx9225, nx9228, 
         nx9234, nx9237, nx9239, nx9244, nx9246, nx9248, nx9250, nx9252, nx9255, 
         nx9257, nx9260, nx9262, nx9265, nx9269, nx9272, nx9275, nx9277, nx9279, 
         nx9282, nx9284, nx9295, nx9297, pres_ow, ip_7, ip_6, ip_5, ip_4, ip_3, 
         ip_2, ip_1, ip_0, tcon_7, tcon_5, tcon_3, tcon_2, tcon_1, tcon_0, ie_7, 
         ie_6, ie_5, ie_4, ie_3, ie_2, ie_1, ie_0, sbuf_7, sbuf_6, sbuf_5, 
         sbuf_4, sbuf_3, sbuf_2, sbuf_1, sbuf_0, pcon_7, pcon_6, pcon_5, pcon_4, 
         pcon_3, pcon_2, pcon_1, pcon_0, scon_7, scon_6, scon_5, scon_4, scon_3, 
         scon_2, scon_1, scon_0, th1_7, th1_6, th1_5, th1_4, th1_3, th1_2, th1_1, 
         th1_0, tl1_7, tl1_6, tl1_5, tl1_4, tl1_3, tl1_2, tl1_1, tl1_0, th0_7, 
         th0_6, th0_5, th0_4, th0_3, th0_2, th0_1, th0_0, tl0_7, tl0_6, tl0_5, 
         tl0_4, tl0_3, tl0_2, tl0_1, tl0_0, tmod_7, tmod_6, tmod_5, tmod_4, 
         tmod_3, tmod_2, tmod_1, tmod_0, rcap2h_7, rcap2h_6, rcap2h_5, rcap2h_4, 
         rcap2h_3, rcap2h_2, rcap2h_1, rcap2h_0, rcap2l_7, rcap2l_6, rcap2l_5, 
         rcap2l_4, rcap2l_3, rcap2l_2, rcap2l_1, rcap2l_0, th2_7, th2_6, th2_5, 
         th2_4, th2_3, th2_2, th2_1, th2_0, tl2_7, tl2_6, tl2_5, tl2_4, tl2_3, 
         tl2_2, tl2_1, tl2_0, t2con_7, t2con_6, t2con_3, t2con_2, t2con_1, 
         t2con_0, psw_5, psw_4, psw_3, psw_2, psw_1, b_reg_7, b_reg_6, b_reg_5, 
         b_reg_4, b_reg_3, b_reg_2, b_reg_1, b_reg_0, tc2_int, brate2, tclk, 
         rclk, tr1, tr0, tf1, tf0, uart_int, p, wr_bit_r_dup_1790, p3_data_7, 
         p3_data_6, p3_data_5, p3_data_4, p3_data_3, p3_data_2, p3_data_1, 
         p3_data_0, p2_data_7, p2_data_6, p2_data_5, p2_data_4, p2_data_3, 
         p2_data_2, p2_data_1, p2_data_0, p1_data_7, p1_data_6, p1_data_5, 
         p1_data_4, p1_data_3, p1_data_2, p1_data_1, p1_data_0, p0_data_7, 
         p0_data_6, p0_data_5, p0_data_4, p0_data_3, p0_data_2, p0_data_1, 
         p0_data_0, prescaler_1, prescaler_0, nx2080, nx1791, nx1792, 
         prescaler_3, prescaler_2, nx2082, nx34, nx1794, nx1796, nx1797, nx1799, 
         nx96, nx1801, nx1804, nx1805, nx158, nx1806, nx1807, nx204, nx1809, 
         nx230, nx236, nx1810, nx1812, nx1813, nx284, nx1814, nx300, nx1817, 
         nx372, nx408, nx1818, nx470, nx1821, nx1822, nx528, nx560, nx1823, 
         nx1825, nx624, nx1827, nx682, nx688, nx696, nx704, nx742, nx1829, nx758, 
         NOT_NOT__68049, nx1830, nx1832, nx1833, nx1834, nx1836, nx1838, nx830, 
         nx1840, nx1841, nx848, nx1843, nx1844, nx1845, nx1846, nx894, nx1848, 
         nx1851, nx918, nx920, nx924, nx932, nx942, nx1853, nx960, nx964, nx1855, 
         nx1856, nx1857, nx1858, nx1860, nx1861, nx1863, nx1016, nx1030, nx1034, 
         nx1864, nx1865, nx1090, nx1116, nx1170, nx1200, nx1226, nx1280, nx1310, 
         nx1336, nx1390, nx1867, nx1446, nx1869, nx1530, nx1871, nx1610, nx1640, 
         nx1666, nx1720, nx1874, nx1875, nx1876, nx1878, nx1879, nx1881, nx1883, 
         nx1884, nx2183, nx2187, nx2189, nx2193, nx1885, nx2201, nx2203, nx1886, 
         nx2210, nx2212, nx2214, nx2217, nx2220, nx2222, nx2227, nx2231, nx2234, 
         nx2236, nx2238, nx2243, nx2245, nx2247, nx2249, nx2251, nx2254, nx2256, 
         nx2259, nx2261, nx2263, nx2265, nx2268, nx2270, nx2274, nx2276, nx2279, 
         nx1888, nx2284, nx2286, nx2289, nx2293, nx2296, nx2300, nx2303, nx2306, 
         nx2310, nx2312, nx2315, nx2317, nx2320, nx1889, nx2325, nx2328, nx2330, 
         nx2333, nx1891, nx2338, nx2340, nx2343, nx2345, nx2347, nx2350, nx2352, 
         nx2354, nx2357, nx2359, nx2361, nx2363, nx2366, nx2368, nx2370, nx2373, 
         nx2375, nx2378, nx2380, nx2383, nx2385, nx2387, nx2389, nx2391, nx1892, 
         nx2396, nx2398, nx2401, nx2403, nx2405, nx2407, nx2409, nx2412, nx1893, 
         nx2416, nx2418, nx2420, nx2422, nx2425, nx2427, nx2429, nx2431, nx2434, 
         nx2436, nx1895, nx2441, nx2443, nx2445, nx2447, nx2450, nx1897, nx2455, 
         nx2458, nx2460, nx1899, nx2465, nx2467, nx2471, nx1902, nx2481, nx1904, 
         nx2486, nx1905, nx2490, nx2495, nx2499, nx2502, nx2505, nx2508, nx1907, 
         nx2515, nx2521, nx2526, nx1908, nx2536, nx2542, nx2544, nx2546, nx2548, 
         nx2550, nx2552, nx2554, nx2557, nx2559, nx2561, nx2564, nx2566, nx2568, 
         nx1909, nx2574, nx2576, nx2578, nx1910, nx2582, nx2584, nx2587, nx2589, 
         nx2591, nx2594, nx2596, nx2598, nx2602, nx1912, nx2606, nx2608, nx2610, 
         nx1913, nx2614, nx2617, nx2619, nx2621, nx2624, nx2626, nx2628, nx2632, 
         nx2634, nx2636, nx1915, nx2640, nx2642, nx2644, nx2647, nx2649, nx2651, 
         nx2654, nx2656, nx1916, nx1918, nx2664, nx2666, nx2668, nx2670, nx2672, 
         nx1919, nx2677, nx2679, nx2681, nx2684, nx1921, nx2688, nx2692, nx2694, 
         nx1923, nx2698, nx2700, nx2702, nx2704, nx2707, nx2709, nx2711, nx2714, 
         nx2716, nx2718, nx1925, nx2724, nx2726, nx2728, nx1927, nx2732, nx2734, 
         nx2737, nx2739, nx2741, nx2744, nx1928, nx2748, cycle_1, cycle_0, 
         NOT_cycle_0, nx386, nx2085, tmp_mul_11, tmp_mul_9, tmp_mul_6, tmp_mul_3, 
         tmp_mul_0, nx42, nx72, nx2087, nx2091, tmp_mul_1, nx2093, nx146, nx2095, 
         tmp_mul_2, nx178, nx2096, nx202, nx210, tmp_mul_4, nx2102, nx2104, 
         nx2105, nx2106, tmp_mul_5, nx2109, tmp_mul_7, tmp_mul_8, nx2110, nx2112, 
         tmp_mul_10, nx374, nx2113, tmp_mul_12, nx2115, tmp_mul_13, NOT_enable, 
         nx415, nx433, nx435, nx437, nx2116, nx2118, nx444, nx449, nx452, nx2122, 
         nx459, nx463, nx468, nx2126, nx474, nx480, nx2127, nx2129, nx489, 
         nx2131, nx495, nx2132, nx500, nx2135, nx504, nx2136, nx510, nx2138, 
         nx515, nx517, nx519, nx524, nx527, nx2139, nx2143, nx2147, nx2149, 
         nx2150, nx2152, nx546, nx2153, nx552, nx2155, nx556, nx558, nx561, 
         nx565, nx2156, nx2159, nx2160, nx579, nx581, nx583, nx2161, nx593, 
         nx2163, nx601, nx2165, nx2167, nx609, nx611, nx613, cycle_1__dup_2348, 
         cycle_0__dup_2349, nx2351, nx730, nx2353, nx104, nx2355, nx2358, 
         tmp_rem_7, nx2362, tmp_rem_6, nx2364, nx2365, tmp_rem_5, nx2367, nx2369, 
         tmp_rem_4, nx2371, tmp_rem_3, nx214, tmp_rem_2, tmp_rem_1, nx238, 
         tmp_rem_0, nx739, nx2372, nx743, nx746, nx334, nx342, nx2374, nx354, 
         nx2376, nx2377, nx2379, nx2381, nx426, nx428, nx2382, nx446, nx464, 
         nx2384, nx482, nx2386, nx2390, nx2392, nx2393, nx2395, nx2397, nx2399, 
         nx2400, nx2402, nx2404, nx590, nx759, nx769, nx2406, nx2408, nx801, 
         nx2410, nx808, nx812, nx2411, nx819, nx821, nx823, nx826, nx829, nx832, 
         nx835, nx841, nx843, nx849, nx851, nx853, nx855, nx861, nx865, nx2413, 
         nx871, nx873, nx879, nx2415, nx884, nx887, nx890, nx893, nx895, nx897, 
         nx901, nx2417, nx907, nx2419, nx913, nx915, nx919, nx923, nx926, nx929, 
         nx931, nx937, nx940, nx2421, nx945, nx2423, nx950, nx953, nx957, nx2424, 
         nx963, nx966, nx2428, nx2432, nx2433, nx2435, nx2437, nx2439, nx2440, 
         nx2442, nx2444, nx1025, nx3204, nx3205, nx3207, nx3208, nx3209, nx3210, 
         nx3211, nx3212, modgen_ram_ix167_a_0__dup_2653, nx3213, nx62, 
         modgen_ram_ix167_a_1__dup_2652, nx3214, modgen_ram_ix167_a_2__dup_2651, 
         nx3215, nx132, modgen_ram_ix167_a_3__dup_2650, nx140, nx166, 
         modgen_ram_ix167_a_4__dup_2649, nx172, modgen_ram_ix167_a_5__dup_2648, 
         nx3216, modgen_ram_ix167_a_6__dup_2647, nx3217, 
         modgen_ram_ix167_a_7__dup_2646, nx3218, nx3219, 
         modgen_ram_ix167_a_8__dup_2645, nx3220, modgen_ram_ix167_a_9__dup_2644, 
         nx292, modgen_ram_ix167_a_10__dup_2643, nx316, nx3221, 
         modgen_ram_ix167_a_11__dup_2642, nx336, nx362, 
         modgen_ram_ix167_a_12__dup_2641, nx3223, 
         modgen_ram_ix167_a_13__dup_2640, nx390, modgen_ram_ix167_a_14__dup_2639, 
         nx3224, modgen_ram_ix167_a_15__dup_2638, nx3225, nx456, nx3226, 
         modgen_ram_ix167_a_16__dup_2637, nx3227, 
         modgen_ram_ix167_a_17__dup_2636, modgen_ram_ix167_a_18__dup_2635, 
         modgen_ram_ix167_a_19__dup_2634, nx3229, 
         modgen_ram_ix167_a_20__dup_2633, modgen_ram_ix167_a_21__dup_2632, 
         modgen_ram_ix167_a_22__dup_2631, modgen_ram_ix167_a_23__dup_2630, nx638, 
         modgen_ram_ix167_a_24__dup_2629, modgen_ram_ix167_a_25__dup_2628, 
         modgen_ram_ix167_a_26__dup_2627, modgen_ram_ix167_a_27__dup_2626, nx726, 
         modgen_ram_ix167_a_28__dup_2625, modgen_ram_ix167_a_29__dup_2624, 
         modgen_ram_ix167_a_30__dup_2623, modgen_ram_ix167_a_31__dup_2622, 
         nx3230, nx818, modgen_ram_ix167_a_32__dup_2621, nx3231, 
         modgen_ram_ix167_a_33__dup_2620, modgen_ram_ix167_a_34__dup_2619, 
         nx3232, modgen_ram_ix167_a_35__dup_2618, nx3233, 
         modgen_ram_ix167_a_36__dup_2617, modgen_ram_ix167_a_37__dup_2616, 
         modgen_ram_ix167_a_38__dup_2615, modgen_ram_ix167_a_39__dup_2614, 
         nx3235, modgen_ram_ix167_a_40__dup_2613, 
         modgen_ram_ix167_a_41__dup_2612, modgen_ram_ix167_a_42__dup_2611, 
         nx3236, modgen_ram_ix167_a_43__dup_2610, nx1088, 
         modgen_ram_ix167_a_44__dup_2609, modgen_ram_ix167_a_45__dup_2608, 
         modgen_ram_ix167_a_46__dup_2607, modgen_ram_ix167_a_47__dup_2606, 
         nx3237, nx3238, modgen_ram_ix167_a_48__dup_2605, nx3239, 
         modgen_ram_ix167_a_49__dup_2604, modgen_ram_ix167_a_50__dup_2603, 
         modgen_ram_ix167_a_51__dup_2602, nx1268, 
         modgen_ram_ix167_a_52__dup_2601, modgen_ram_ix167_a_53__dup_2600, 
         modgen_ram_ix167_a_54__dup_2599, modgen_ram_ix167_a_55__dup_2598, 
         nx3240, modgen_ram_ix167_a_56__dup_2597, 
         modgen_ram_ix167_a_57__dup_2596, modgen_ram_ix167_a_58__dup_2595, 
         modgen_ram_ix167_a_59__dup_2594, nx1440, 
         modgen_ram_ix167_a_60__dup_2593, modgen_ram_ix167_a_61__dup_2592, 
         modgen_ram_ix167_a_62__dup_2591, modgen_ram_ix167_a_63__dup_2590, 
         nx1524, nx1532, nx1544, modgen_ram_ix167_a_64__dup_2589, nx1550, 
         modgen_ram_ix167_a_65__dup_2588, modgen_ram_ix167_a_66__dup_2587, 
         nx1608, modgen_ram_ix167_a_67__dup_2586, nx1634, 
         modgen_ram_ix167_a_68__dup_2585, modgen_ram_ix167_a_69__dup_2584, 
         modgen_ram_ix167_a_70__dup_2583, modgen_ram_ix167_a_71__dup_2582, 
         nx3241, modgen_ram_ix167_a_72__dup_2581, 
         modgen_ram_ix167_a_73__dup_2580, modgen_ram_ix167_a_74__dup_2579, 
         nx3242, modgen_ram_ix167_a_75__dup_2578, nx3243, 
         modgen_ram_ix167_a_76__dup_2577, modgen_ram_ix167_a_77__dup_2576, 
         modgen_ram_ix167_a_78__dup_2575, modgen_ram_ix167_a_79__dup_2574, 
         nx3244, nx3245, modgen_ram_ix167_a_80__dup_2573, nx3247, 
         modgen_ram_ix167_a_81__dup_2572, modgen_ram_ix167_a_82__dup_2571, 
         modgen_ram_ix167_a_83__dup_2570, nx1980, 
         modgen_ram_ix167_a_84__dup_2569, modgen_ram_ix167_a_85__dup_2568, 
         modgen_ram_ix167_a_86__dup_2567, modgen_ram_ix167_a_87__dup_2566, 
         nx2064, modgen_ram_ix167_a_88__dup_2565, 
         modgen_ram_ix167_a_89__dup_2564, modgen_ram_ix167_a_90__dup_2563, 
         modgen_ram_ix167_a_91__dup_2562, nx3248, 
         modgen_ram_ix167_a_92__dup_2561, modgen_ram_ix167_a_93__dup_2560, 
         modgen_ram_ix167_a_94__dup_2559, modgen_ram_ix167_a_95__dup_2558, 
         nx3249, nx2244, modgen_ram_ix167_a_96__dup_2557, nx3250, 
         modgen_ram_ix167_a_97__dup_2556, modgen_ram_ix167_a_98__dup_2555, 
         nx3251, modgen_ram_ix167_a_99__dup_2554, nx3252, 
         modgen_ram_ix167_a_100__dup_2553, modgen_ram_ix167_a_101__dup_2552, 
         modgen_ram_ix167_a_102__dup_2551, modgen_ram_ix167_a_103__dup_2550, 
         nx3253, modgen_ram_ix167_a_104__dup_2549, 
         modgen_ram_ix167_a_105__dup_2548, modgen_ram_ix167_a_106__dup_2547, 
         nx3255, modgen_ram_ix167_a_107__dup_2546, nx2510, 
         modgen_ram_ix167_a_108__dup_2545, modgen_ram_ix167_a_109__dup_2544, 
         modgen_ram_ix167_a_110__dup_2543, modgen_ram_ix167_a_111__dup_2542, 
         nx2590, nx3256, modgen_ram_ix167_a_112__dup_2541, nx3257, 
         modgen_ram_ix167_a_113__dup_2540, modgen_ram_ix167_a_114__dup_2539, 
         modgen_ram_ix167_a_115__dup_2538, nx3258, 
         modgen_ram_ix167_a_116__dup_2537, modgen_ram_ix167_a_117__dup_2536, 
         modgen_ram_ix167_a_118__dup_2535, modgen_ram_ix167_a_119__dup_2534, 
         nx2768, modgen_ram_ix167_a_120__dup_2533, 
         modgen_ram_ix167_a_121__dup_2532, modgen_ram_ix167_a_122__dup_2531, 
         modgen_ram_ix167_a_123__dup_2530, nx2856, 
         modgen_ram_ix167_a_124__dup_2529, modgen_ram_ix167_a_125__dup_2528, 
         modgen_ram_ix167_a_126__dup_2527, modgen_ram_ix167_a_127__dup_2526, 
         nx2940, nx2948, nx2956, nx2964, modgen_ram_ix167_a_128__dup_2525, 
         nx2970, modgen_ram_ix167_a_129__dup_2524, 
         modgen_ram_ix167_a_130__dup_2523, nx3028, 
         modgen_ram_ix167_a_131__dup_2522, nx3054, 
         modgen_ram_ix167_a_132__dup_2521, modgen_ram_ix167_a_133__dup_2520, 
         modgen_ram_ix167_a_134__dup_2519, modgen_ram_ix167_a_135__dup_2518, 
         nx3134, modgen_ram_ix167_a_136__dup_2517, 
         modgen_ram_ix167_a_137__dup_2516, modgen_ram_ix167_a_138__dup_2515, 
         nx3200, modgen_ram_ix167_a_139__dup_2514, nx3259, 
         modgen_ram_ix167_a_140__dup_2513, modgen_ram_ix167_a_141__dup_2512, 
         modgen_ram_ix167_a_142__dup_2511, modgen_ram_ix167_a_143__dup_2510, 
         nx3306, nx3318, modgen_ram_ix167_a_144__dup_2509, nx3320, 
         modgen_ram_ix167_a_145__dup_2508, modgen_ram_ix167_a_146__dup_2507, 
         modgen_ram_ix167_a_147__dup_2506, nx3400, 
         modgen_ram_ix167_a_148__dup_2505, modgen_ram_ix167_a_149__dup_2504, 
         modgen_ram_ix167_a_150__dup_2503, modgen_ram_ix167_a_151__dup_2502, 
         nx3260, modgen_ram_ix167_a_152__dup_2501, 
         modgen_ram_ix167_a_153__dup_2500, modgen_ram_ix167_a_154__dup_2499, 
         modgen_ram_ix167_a_155__dup_2498, nx3572, 
         modgen_ram_ix167_a_156__dup_2497, modgen_ram_ix167_a_157__dup_2496, 
         modgen_ram_ix167_a_158__dup_2495, modgen_ram_ix167_a_159__dup_2494, 
         nx3261, nx3664, modgen_ram_ix167_a_160__dup_2493, nx3674, 
         modgen_ram_ix167_a_161__dup_2492, modgen_ram_ix167_a_162__dup_2491, 
         nx3732, modgen_ram_ix167_a_163__dup_2490, nx3758, 
         modgen_ram_ix167_a_164__dup_2489, modgen_ram_ix167_a_165__dup_2488, 
         modgen_ram_ix167_a_166__dup_2487, modgen_ram_ix167_a_167__dup_2486, 
         nx3838, modgen_ram_ix167_a_168__dup_2485, 
         modgen_ram_ix167_a_169__dup_2484, modgen_ram_ix167_a_170__dup_2483, 
         nx3904, modgen_ram_ix167_a_171__dup_2482, nx3930, 
         modgen_ram_ix167_a_172__dup_2481, modgen_ram_ix167_a_173__dup_2480, 
         modgen_ram_ix167_a_174__dup_2479, modgen_ram_ix167_a_175__dup_2478, 
         nx4010, nx4022, modgen_ram_ix167_a_176__dup_2477, nx4024, 
         modgen_ram_ix167_a_177__dup_2476, modgen_ram_ix167_a_178__dup_2475, 
         modgen_ram_ix167_a_179__dup_2474, nx4104, 
         modgen_ram_ix167_a_180__dup_2473, modgen_ram_ix167_a_181__dup_2472, 
         modgen_ram_ix167_a_182__dup_2471, modgen_ram_ix167_a_183__dup_2470, 
         nx3262, modgen_ram_ix167_a_184__dup_2469, 
         modgen_ram_ix167_a_185__dup_2468, modgen_ram_ix167_a_186__dup_2467, 
         modgen_ram_ix167_a_187__dup_2466, nx4276, 
         modgen_ram_ix167_a_188__dup_2465, modgen_ram_ix167_a_189__dup_2464, 
         modgen_ram_ix167_a_190__dup_2463, modgen_ram_ix167_a_191__dup_2462, 
         nx4360, nx4368, nx4380, modgen_ram_ix167_a_192__dup_2461, nx3263, 
         modgen_ram_ix167_a_193__dup_2460, modgen_ram_ix167_a_194__dup_2459, 
         nx3264, modgen_ram_ix167_a_195__dup_2458, nx4472, 
         modgen_ram_ix167_a_196__dup_2457, modgen_ram_ix167_a_197__dup_2456, 
         modgen_ram_ix167_a_198__dup_2455, modgen_ram_ix167_a_199__dup_2454, 
         nx4552, modgen_ram_ix167_a_200__dup_2453, 
         modgen_ram_ix167_a_201__dup_2452, modgen_ram_ix167_a_202__dup_2451, 
         nx4618, modgen_ram_ix167_a_203__dup_2450, nx4644, 
         modgen_ram_ix167_a_204__dup_2449, modgen_ram_ix167_a_205__dup_2448, 
         modgen_ram_ix167_a_206__dup_2447, modgen_ram_ix167_a_207__dup_2446, 
         nx4724, nx4736, modgen_ram_ix167_a_208__dup_2445, nx4738, 
         modgen_ram_ix167_a_209__dup_2444, modgen_ram_ix167_a_210__dup_2443, 
         modgen_ram_ix167_a_211__dup_2442, nx4818, 
         modgen_ram_ix167_a_212__dup_2441, modgen_ram_ix167_a_213__dup_2440, 
         modgen_ram_ix167_a_214__dup_2439, modgen_ram_ix167_a_215__dup_2438, 
         nx4902, modgen_ram_ix167_a_216__dup_2437, 
         modgen_ram_ix167_a_217__dup_2436, modgen_ram_ix167_a_218__dup_2435, 
         modgen_ram_ix167_a_219__dup_2434, nx4990, 
         modgen_ram_ix167_a_220__dup_2433, modgen_ram_ix167_a_221__dup_2432, 
         modgen_ram_ix167_a_222__dup_2431, modgen_ram_ix167_a_223__dup_2430, 
         nx5074, nx5082, modgen_ram_ix167_a_224__dup_2429, nx5092, 
         modgen_ram_ix167_a_225__dup_2428, modgen_ram_ix167_a_226__dup_2427, 
         nx5150, modgen_ram_ix167_a_227__dup_2426, nx5176, 
         modgen_ram_ix167_a_228__dup_2425, modgen_ram_ix167_a_229__dup_2424, 
         modgen_ram_ix167_a_230__dup_2423, modgen_ram_ix167_a_231__dup_2422, 
         nx5256, modgen_ram_ix167_a_232__dup_2421, 
         modgen_ram_ix167_a_233__dup_2420, modgen_ram_ix167_a_234__dup_2419, 
         nx5322, modgen_ram_ix167_a_235__dup_2418, nx5348, 
         modgen_ram_ix167_a_236__dup_2417, modgen_ram_ix167_a_237__dup_2416, 
         modgen_ram_ix167_a_238__dup_2415, modgen_ram_ix167_a_239__dup_2414, 
         nx5428, nx5440, modgen_ram_ix167_a_240__dup_2413, nx5442, 
         modgen_ram_ix167_a_241__dup_2412, modgen_ram_ix167_a_242__dup_2411, 
         modgen_ram_ix167_a_243__dup_2410, nx5522, 
         modgen_ram_ix167_a_244__dup_2409, modgen_ram_ix167_a_245__dup_2408, 
         modgen_ram_ix167_a_246__dup_2407, modgen_ram_ix167_a_247__dup_2406, 
         nx5606, modgen_ram_ix167_a_248__dup_2405, 
         modgen_ram_ix167_a_249__dup_2404, modgen_ram_ix167_a_250__dup_2403, 
         modgen_ram_ix167_a_251__dup_2402, nx3265, 
         modgen_ram_ix167_a_252__dup_2401, modgen_ram_ix167_a_253__dup_2400, 
         modgen_ram_ix167_a_254__dup_2399, modgen_ram_ix167_a_255__dup_2398, 
         nx5778, nx5786, nx5796, nx5810, modgen_ram_ix167_a_0__dup_2389, 
         modgen_ram_ix167_a_1__dup_2388, modgen_ram_ix167_a_2__dup_2387, nx5848, 
         modgen_ram_ix167_a_3__dup_2386, nx5866, modgen_ram_ix167_a_4__dup_2385, 
         modgen_ram_ix167_a_5__dup_2384, modgen_ram_ix167_a_6__dup_2383, 
         modgen_ram_ix167_a_7__dup_2382, nx3267, modgen_ram_ix167_a_8__dup_2381, 
         modgen_ram_ix167_a_9__dup_2380, modgen_ram_ix167_a_10__dup_2379, nx5956, 
         modgen_ram_ix167_a_11__dup_2378, nx3268, 
         modgen_ram_ix167_a_12__dup_2377, modgen_ram_ix167_a_13__dup_2376, 
         modgen_ram_ix167_a_14__dup_2375, modgen_ram_ix167_a_15__dup_2374, 
         nx6022, nx3269, modgen_ram_ix167_a_16__dup_2373, 
         modgen_ram_ix167_a_17__dup_2372, modgen_ram_ix167_a_18__dup_2371, 
         modgen_ram_ix167_a_19__dup_2370, nx6082, 
         modgen_ram_ix167_a_20__dup_2369, modgen_ram_ix167_a_21__dup_2368, 
         modgen_ram_ix167_a_22__dup_2367, modgen_ram_ix167_a_23__dup_2366, 
         nx3270, modgen_ram_ix167_a_24__dup_2365, 
         modgen_ram_ix167_a_25__dup_2364, modgen_ram_ix167_a_26__dup_2363, 
         modgen_ram_ix167_a_27__dup_2362, nx6190, 
         modgen_ram_ix167_a_28__dup_2361, modgen_ram_ix167_a_29__dup_2360, 
         modgen_ram_ix167_a_30__dup_2359, modgen_ram_ix167_a_31__dup_2358, 
         nx6242, nx6250, modgen_ram_ix167_a_32__dup_2357, 
         modgen_ram_ix167_a_33__dup_2356, modgen_ram_ix167_a_34__dup_2355, 
         nx6292, modgen_ram_ix167_a_35__dup_2354, nx6310, 
         modgen_ram_ix167_a_36__dup_2353, modgen_ram_ix167_a_37__dup_2352, 
         modgen_ram_ix167_a_38__dup_2351, modgen_ram_ix167_a_39__dup_2350, 
         nx6358, modgen_ram_ix167_a_40__dup_2349, 
         modgen_ram_ix167_a_41__dup_2348, modgen_ram_ix167_a_42__dup_2347, 
         nx6400, modgen_ram_ix167_a_43__dup_2346, nx6418, 
         modgen_ram_ix167_a_44__dup_2345, modgen_ram_ix167_a_45__dup_2344, 
         modgen_ram_ix167_a_46__dup_2343, modgen_ram_ix167_a_47__dup_2342, 
         nx6466, nx6478, modgen_ram_ix167_a_48__dup_2341, 
         modgen_ram_ix167_a_49__dup_2340, modgen_ram_ix167_a_50__dup_2339, 
         modgen_ram_ix167_a_51__dup_2338, nx6526, 
         modgen_ram_ix167_a_52__dup_2337, modgen_ram_ix167_a_53__dup_2336, 
         modgen_ram_ix167_a_54__dup_2335, modgen_ram_ix167_a_55__dup_2334, 
         nx6578, modgen_ram_ix167_a_56__dup_2333, 
         modgen_ram_ix167_a_57__dup_2332, modgen_ram_ix167_a_58__dup_2331, 
         modgen_ram_ix167_a_59__dup_2330, nx6634, 
         modgen_ram_ix167_a_60__dup_2329, modgen_ram_ix167_a_61__dup_2328, 
         modgen_ram_ix167_a_62__dup_2327, modgen_ram_ix167_a_63__dup_2326, 
         nx6686, nx6694, nx6706, modgen_ram_ix167_a_64__dup_2325, 
         modgen_ram_ix167_a_65__dup_2324, modgen_ram_ix167_a_66__dup_2323, 
         nx6740, modgen_ram_ix167_a_67__dup_2322, nx6758, 
         modgen_ram_ix167_a_68__dup_2321, modgen_ram_ix167_a_69__dup_2320, 
         modgen_ram_ix167_a_70__dup_2319, modgen_ram_ix167_a_71__dup_2318, 
         nx6806, modgen_ram_ix167_a_72__dup_2317, 
         modgen_ram_ix167_a_73__dup_2316, modgen_ram_ix167_a_74__dup_2315, 
         nx6848, modgen_ram_ix167_a_75__dup_2314, nx6866, 
         modgen_ram_ix167_a_76__dup_2313, modgen_ram_ix167_a_77__dup_2312, 
         modgen_ram_ix167_a_78__dup_2311, modgen_ram_ix167_a_79__dup_2310, 
         nx3271, nx6926, modgen_ram_ix167_a_80__dup_2309, 
         modgen_ram_ix167_a_81__dup_2308, modgen_ram_ix167_a_82__dup_2307, 
         modgen_ram_ix167_a_83__dup_2306, nx6974, 
         modgen_ram_ix167_a_84__dup_2305, modgen_ram_ix167_a_85__dup_2304, 
         modgen_ram_ix167_a_86__dup_2303, modgen_ram_ix167_a_87__dup_2302, 
         nx7026, modgen_ram_ix167_a_88__dup_2301, 
         modgen_ram_ix167_a_89__dup_2300, modgen_ram_ix167_a_90__dup_2299, 
         modgen_ram_ix167_a_91__dup_2298, nx7082, 
         modgen_ram_ix167_a_92__dup_2297, modgen_ram_ix167_a_93__dup_2296, 
         modgen_ram_ix167_a_94__dup_2295, modgen_ram_ix167_a_95__dup_2294, 
         nx3272, nx7142, modgen_ram_ix167_a_96__dup_2293, 
         modgen_ram_ix167_a_97__dup_2292, modgen_ram_ix167_a_98__dup_2291, 
         nx7184, modgen_ram_ix167_a_99__dup_2290, nx7202, 
         modgen_ram_ix167_a_100__dup_2289, modgen_ram_ix167_a_101__dup_2288, 
         modgen_ram_ix167_a_102__dup_2287, modgen_ram_ix167_a_103__dup_2286, 
         nx7250, modgen_ram_ix167_a_104__dup_2285, 
         modgen_ram_ix167_a_105__dup_2284, modgen_ram_ix167_a_106__dup_2283, 
         nx7292, modgen_ram_ix167_a_107__dup_2282, nx7310, 
         modgen_ram_ix167_a_108__dup_2281, modgen_ram_ix167_a_109__dup_2280, 
         modgen_ram_ix167_a_110__dup_2279, modgen_ram_ix167_a_111__dup_2278, 
         nx7358, nx7370, modgen_ram_ix167_a_112__dup_2277, 
         modgen_ram_ix167_a_113__dup_2276, modgen_ram_ix167_a_114__dup_2275, 
         modgen_ram_ix167_a_115__dup_2274, nx7418, 
         modgen_ram_ix167_a_116__dup_2273, modgen_ram_ix167_a_117__dup_2272, 
         modgen_ram_ix167_a_118__dup_2271, modgen_ram_ix167_a_119__dup_2270, 
         nx7470, modgen_ram_ix167_a_120__dup_2269, 
         modgen_ram_ix167_a_121__dup_2268, modgen_ram_ix167_a_122__dup_2267, 
         modgen_ram_ix167_a_123__dup_2266, nx3273, 
         modgen_ram_ix167_a_124__dup_2265, modgen_ram_ix167_a_125__dup_2264, 
         modgen_ram_ix167_a_126__dup_2263, modgen_ram_ix167_a_127__dup_2262, 
         nx7578, nx3275, nx7594, nx7602, modgen_ram_ix167_a_128__dup_2261, 
         modgen_ram_ix167_a_129__dup_2260, modgen_ram_ix167_a_130__dup_2259, 
         nx7636, modgen_ram_ix167_a_131__dup_2258, nx3276, 
         modgen_ram_ix167_a_132__dup_2257, modgen_ram_ix167_a_133__dup_2256, 
         modgen_ram_ix167_a_134__dup_2255, modgen_ram_ix167_a_135__dup_2254, 
         nx7702, modgen_ram_ix167_a_136__dup_2253, 
         modgen_ram_ix167_a_137__dup_2252, modgen_ram_ix167_a_138__dup_2251, 
         nx3277, modgen_ram_ix167_a_139__dup_2250, nx7762, 
         modgen_ram_ix167_a_140__dup_2249, modgen_ram_ix167_a_141__dup_2248, 
         modgen_ram_ix167_a_142__dup_2247, modgen_ram_ix167_a_143__dup_2246, 
         nx7810, nx7822, modgen_ram_ix167_a_144__dup_2245, 
         modgen_ram_ix167_a_145__dup_2244, modgen_ram_ix167_a_146__dup_2243, 
         modgen_ram_ix167_a_147__dup_2242, nx7870, 
         modgen_ram_ix167_a_148__dup_2241, modgen_ram_ix167_a_149__dup_2240, 
         modgen_ram_ix167_a_150__dup_2239, modgen_ram_ix167_a_151__dup_2238, 
         nx7922, modgen_ram_ix167_a_152__dup_2237, 
         modgen_ram_ix167_a_153__dup_2236, modgen_ram_ix167_a_154__dup_2235, 
         modgen_ram_ix167_a_155__dup_2234, nx7978, 
         modgen_ram_ix167_a_156__dup_2233, modgen_ram_ix167_a_157__dup_2232, 
         modgen_ram_ix167_a_158__dup_2231, modgen_ram_ix167_a_159__dup_2230, 
         nx8030, nx8038, modgen_ram_ix167_a_160__dup_2229, 
         modgen_ram_ix167_a_161__dup_2228, modgen_ram_ix167_a_162__dup_2227, 
         nx8080, modgen_ram_ix167_a_163__dup_2226, nx3278, 
         modgen_ram_ix167_a_164__dup_2225, modgen_ram_ix167_a_165__dup_2224, 
         modgen_ram_ix167_a_166__dup_2223, modgen_ram_ix167_a_167__dup_2222, 
         nx8146, modgen_ram_ix167_a_168__dup_2221, 
         modgen_ram_ix167_a_169__dup_2220, modgen_ram_ix167_a_170__dup_2219, 
         nx8188, modgen_ram_ix167_a_171__dup_2218, nx8206, 
         modgen_ram_ix167_a_172__dup_2217, modgen_ram_ix167_a_173__dup_2216, 
         modgen_ram_ix167_a_174__dup_2215, modgen_ram_ix167_a_175__dup_2214, 
         nx8254, nx8266, modgen_ram_ix167_a_176__dup_2213, 
         modgen_ram_ix167_a_177__dup_2212, modgen_ram_ix167_a_178__dup_2211, 
         modgen_ram_ix167_a_179__dup_2210, nx8314, 
         modgen_ram_ix167_a_180__dup_2209, modgen_ram_ix167_a_181__dup_2208, 
         modgen_ram_ix167_a_182__dup_2207, modgen_ram_ix167_a_183__dup_2206, 
         nx8366, modgen_ram_ix167_a_184__dup_2205, 
         modgen_ram_ix167_a_185__dup_2204, modgen_ram_ix167_a_186__dup_2203, 
         modgen_ram_ix167_a_187__dup_2202, nx3279, 
         modgen_ram_ix167_a_188__dup_2201, modgen_ram_ix167_a_189__dup_2200, 
         modgen_ram_ix167_a_190__dup_2199, modgen_ram_ix167_a_191__dup_2198, 
         nx3280, nx8482, nx3281, modgen_ram_ix167_a_192__dup_2197, 
         modgen_ram_ix167_a_193__dup_2196, modgen_ram_ix167_a_194__dup_2195, 
         nx3282, modgen_ram_ix167_a_195__dup_2194, nx3283, 
         modgen_ram_ix167_a_196__dup_2193, modgen_ram_ix167_a_197__dup_2192, 
         modgen_ram_ix167_a_198__dup_2191, modgen_ram_ix167_a_199__dup_2190, 
         nx8594, modgen_ram_ix167_a_200__dup_2189, 
         modgen_ram_ix167_a_201__dup_2188, modgen_ram_ix167_a_202__dup_2187, 
         nx8636, modgen_ram_ix167_a_203__dup_2186, nx8654, 
         modgen_ram_ix167_a_204__dup_2185, modgen_ram_ix167_a_205__dup_2184, 
         modgen_ram_ix167_a_206__dup_2183, modgen_ram_ix167_a_207__dup_2182, 
         nx8702, nx8714, modgen_ram_ix167_a_208__dup_2181, 
         modgen_ram_ix167_a_209__dup_2180, modgen_ram_ix167_a_210__dup_2179, 
         modgen_ram_ix167_a_211__dup_2178, nx8762, 
         modgen_ram_ix167_a_212__dup_2177, modgen_ram_ix167_a_213__dup_2176, 
         modgen_ram_ix167_a_214__dup_2175, modgen_ram_ix167_a_215__dup_2174, 
         nx8814, modgen_ram_ix167_a_216__dup_2173, 
         modgen_ram_ix167_a_217__dup_2172, modgen_ram_ix167_a_218__dup_2171, 
         modgen_ram_ix167_a_219__dup_2170, nx8870, 
         modgen_ram_ix167_a_220__dup_2169, modgen_ram_ix167_a_221__dup_2168, 
         modgen_ram_ix167_a_222__dup_2167, modgen_ram_ix167_a_223__dup_2166, 
         nx8922, nx3284, modgen_ram_ix167_a_224__dup_2165, 
         modgen_ram_ix167_a_225__dup_2164, modgen_ram_ix167_a_226__dup_2163, 
         nx8972, modgen_ram_ix167_a_227__dup_2162, nx8990, 
         modgen_ram_ix167_a_228__dup_2161, modgen_ram_ix167_a_229__dup_2160, 
         modgen_ram_ix167_a_230__dup_2159, modgen_ram_ix167_a_231__dup_2158, 
         nx3285, modgen_ram_ix167_a_232__dup_2157, 
         modgen_ram_ix167_a_233__dup_2156, modgen_ram_ix167_a_234__dup_2155, 
         nx9080, modgen_ram_ix167_a_235__dup_2154, nx9098, 
         modgen_ram_ix167_a_236__dup_2153, modgen_ram_ix167_a_237__dup_2152, 
         modgen_ram_ix167_a_238__dup_2151, modgen_ram_ix167_a_239__dup_2150, 
         nx9146, nx9158, modgen_ram_ix167_a_240__dup_2149, 
         modgen_ram_ix167_a_241__dup_2148, modgen_ram_ix167_a_242__dup_2147, 
         modgen_ram_ix167_a_243__dup_2146, nx9206, 
         modgen_ram_ix167_a_244__dup_2145, modgen_ram_ix167_a_245__dup_2144, 
         modgen_ram_ix167_a_246__dup_2143, modgen_ram_ix167_a_247__dup_2142, 
         nx9258, modgen_ram_ix167_a_248__dup_2141, 
         modgen_ram_ix167_a_249__dup_2140, modgen_ram_ix167_a_250__dup_2139, 
         modgen_ram_ix167_a_251__dup_2138, nx9314, 
         modgen_ram_ix167_a_252__dup_2137, modgen_ram_ix167_a_253__dup_2136, 
         modgen_ram_ix167_a_254__dup_2135, modgen_ram_ix167_a_255__dup_2134, 
         nx9366, nx9374, nx9384, nx9398, modgen_ram_ix167_a_0__dup_2125, 
         modgen_ram_ix167_a_1__dup_2124, modgen_ram_ix167_a_2__dup_2123, nx9436, 
         modgen_ram_ix167_a_3__dup_2122, nx9454, modgen_ram_ix167_a_4__dup_2121, 
         modgen_ram_ix167_a_5__dup_2120, modgen_ram_ix167_a_6__dup_2119, 
         modgen_ram_ix167_a_7__dup_2118, nx9502, modgen_ram_ix167_a_8__dup_2117, 
         modgen_ram_ix167_a_9__dup_2116, modgen_ram_ix167_a_10__dup_2115, nx9544, 
         modgen_ram_ix167_a_11__dup_2114, nx9562, 
         modgen_ram_ix167_a_12__dup_2113, modgen_ram_ix167_a_13__dup_2112, 
         modgen_ram_ix167_a_14__dup_2111, modgen_ram_ix167_a_15__dup_2110, 
         nx9610, nx9622, modgen_ram_ix167_a_16__dup_2109, 
         modgen_ram_ix167_a_17__dup_2108, modgen_ram_ix167_a_18__dup_2107, 
         modgen_ram_ix167_a_19__dup_2106, nx9670, 
         modgen_ram_ix167_a_20__dup_2105, modgen_ram_ix167_a_21__dup_2104, 
         modgen_ram_ix167_a_22__dup_2103, modgen_ram_ix167_a_23__dup_2102, 
         nx9722, modgen_ram_ix167_a_24__dup_2101, 
         modgen_ram_ix167_a_25__dup_2100, modgen_ram_ix167_a_26__dup_2099, 
         modgen_ram_ix167_a_27__dup_2098, nx9778, 
         modgen_ram_ix167_a_28__dup_2097, modgen_ram_ix167_a_29__dup_2096, 
         modgen_ram_ix167_a_30__dup_2095, modgen_ram_ix167_a_31__dup_2094, 
         nx9830, nx9838, modgen_ram_ix167_a_32__dup_2093, 
         modgen_ram_ix167_a_33__dup_2092, modgen_ram_ix167_a_34__dup_2091, 
         nx9880, modgen_ram_ix167_a_35__dup_2090, nx9898, 
         modgen_ram_ix167_a_36__dup_2089, modgen_ram_ix167_a_37__dup_2088, 
         modgen_ram_ix167_a_38__dup_2087, modgen_ram_ix167_a_39__dup_2086, 
         nx9946, modgen_ram_ix167_a_40__dup_2085, 
         modgen_ram_ix167_a_41__dup_2084, modgen_ram_ix167_a_42__dup_2083, 
         nx9988, modgen_ram_ix167_a_43__dup_2082, nx10006, 
         modgen_ram_ix167_a_44__dup_2081, modgen_ram_ix167_a_45__dup_2080, 
         modgen_ram_ix167_a_46__dup_2079, modgen_ram_ix167_a_47__dup_2078, 
         nx10054, nx10066, modgen_ram_ix167_a_48__dup_2077, 
         modgen_ram_ix167_a_49__dup_2076, modgen_ram_ix167_a_50__dup_2075, 
         modgen_ram_ix167_a_51__dup_2074, nx10114, 
         modgen_ram_ix167_a_52__dup_2073, modgen_ram_ix167_a_53__dup_2072, 
         modgen_ram_ix167_a_54__dup_2071, modgen_ram_ix167_a_55__dup_2070, 
         nx10166, modgen_ram_ix167_a_56__dup_2069, 
         modgen_ram_ix167_a_57__dup_2068, modgen_ram_ix167_a_58__dup_2067, 
         modgen_ram_ix167_a_59__dup_2066, nx10222, 
         modgen_ram_ix167_a_60__dup_2065, modgen_ram_ix167_a_61__dup_2064, 
         modgen_ram_ix167_a_62__dup_2063, modgen_ram_ix167_a_63__dup_2062, 
         nx10274, nx10282, nx10294, modgen_ram_ix167_a_64__dup_2061, 
         modgen_ram_ix167_a_65__dup_2060, modgen_ram_ix167_a_66__dup_2059, 
         nx10328, modgen_ram_ix167_a_67__dup_2058, nx10346, 
         modgen_ram_ix167_a_68__dup_2057, modgen_ram_ix167_a_69__dup_2056, 
         modgen_ram_ix167_a_70__dup_2055, modgen_ram_ix167_a_71__dup_2054, 
         nx10394, modgen_ram_ix167_a_72__dup_2053, 
         modgen_ram_ix167_a_73__dup_2052, modgen_ram_ix167_a_74__dup_2051, 
         nx10436, modgen_ram_ix167_a_75__dup_2050, nx10454, 
         modgen_ram_ix167_a_76__dup_2049, modgen_ram_ix167_a_77__dup_2048, 
         modgen_ram_ix167_a_78__dup_2047, modgen_ram_ix167_a_79__dup_2046, 
         nx10502, nx10514, modgen_ram_ix167_a_80__dup_2045, 
         modgen_ram_ix167_a_81__dup_2044, modgen_ram_ix167_a_82__dup_2043, 
         modgen_ram_ix167_a_83__dup_2042, nx10562, 
         modgen_ram_ix167_a_84__dup_2041, modgen_ram_ix167_a_85__dup_2040, 
         modgen_ram_ix167_a_86__dup_2039, modgen_ram_ix167_a_87__dup_2038, 
         nx10614, modgen_ram_ix167_a_88__dup_2037, 
         modgen_ram_ix167_a_89__dup_2036, modgen_ram_ix167_a_90__dup_2035, 
         modgen_ram_ix167_a_91__dup_2034, nx10670, 
         modgen_ram_ix167_a_92__dup_2033, modgen_ram_ix167_a_93__dup_2032, 
         modgen_ram_ix167_a_94__dup_2031, modgen_ram_ix167_a_95__dup_2030, 
         nx10722, nx10730, modgen_ram_ix167_a_96__dup_2029, 
         modgen_ram_ix167_a_97__dup_2028, modgen_ram_ix167_a_98__dup_2027, 
         nx10772, modgen_ram_ix167_a_99__dup_2026, nx10790, 
         modgen_ram_ix167_a_100__dup_2025, modgen_ram_ix167_a_101__dup_2024, 
         modgen_ram_ix167_a_102__dup_2023, modgen_ram_ix167_a_103__dup_2022, 
         nx10838, modgen_ram_ix167_a_104__dup_2021, 
         modgen_ram_ix167_a_105__dup_2020, modgen_ram_ix167_a_106__dup_2019, 
         nx10880, modgen_ram_ix167_a_107__dup_2018, nx10898, 
         modgen_ram_ix167_a_108__dup_2017, modgen_ram_ix167_a_109__dup_2016, 
         modgen_ram_ix167_a_110__dup_2015, modgen_ram_ix167_a_111__dup_2014, 
         nx10946, nx10958, modgen_ram_ix167_a_112__dup_2013, 
         modgen_ram_ix167_a_113__dup_2012, modgen_ram_ix167_a_114__dup_2011, 
         modgen_ram_ix167_a_115__dup_2010, nx11006, 
         modgen_ram_ix167_a_116__dup_2009, modgen_ram_ix167_a_117__dup_2008, 
         modgen_ram_ix167_a_118__dup_2007, modgen_ram_ix167_a_119__dup_2006, 
         nx11058, modgen_ram_ix167_a_120__dup_2005, 
         modgen_ram_ix167_a_121__dup_2004, modgen_ram_ix167_a_122__dup_2003, 
         modgen_ram_ix167_a_123__dup_2002, nx11114, 
         modgen_ram_ix167_a_124__dup_2001, modgen_ram_ix167_a_125__dup_2000, 
         modgen_ram_ix167_a_126__dup_1999, modgen_ram_ix167_a_127__dup_1998, 
         nx11166, nx11174, nx11182, nx11190, modgen_ram_ix167_a_128__dup_1997, 
         modgen_ram_ix167_a_129__dup_1996, modgen_ram_ix167_a_130__dup_1995, 
         nx11224, modgen_ram_ix167_a_131__dup_1994, nx11242, 
         modgen_ram_ix167_a_132__dup_1993, modgen_ram_ix167_a_133__dup_1992, 
         modgen_ram_ix167_a_134__dup_1991, modgen_ram_ix167_a_135__dup_1990, 
         nx11290, modgen_ram_ix167_a_136__dup_1989, 
         modgen_ram_ix167_a_137__dup_1988, modgen_ram_ix167_a_138__dup_1987, 
         nx11332, modgen_ram_ix167_a_139__dup_1986, nx11350, 
         modgen_ram_ix167_a_140__dup_1985, modgen_ram_ix167_a_141__dup_1984, 
         modgen_ram_ix167_a_142__dup_1983, modgen_ram_ix167_a_143__dup_1982, 
         nx11398, nx11410, modgen_ram_ix167_a_144__dup_1981, 
         modgen_ram_ix167_a_145__dup_1980, modgen_ram_ix167_a_146__dup_1979, 
         modgen_ram_ix167_a_147__dup_1978, nx11458, 
         modgen_ram_ix167_a_148__dup_1977, modgen_ram_ix167_a_149__dup_1976, 
         modgen_ram_ix167_a_150__dup_1975, modgen_ram_ix167_a_151__dup_1974, 
         nx11510, modgen_ram_ix167_a_152__dup_1973, 
         modgen_ram_ix167_a_153__dup_1972, modgen_ram_ix167_a_154__dup_1971, 
         modgen_ram_ix167_a_155__dup_1970, nx11566, 
         modgen_ram_ix167_a_156__dup_1969, modgen_ram_ix167_a_157__dup_1968, 
         modgen_ram_ix167_a_158__dup_1967, modgen_ram_ix167_a_159__dup_1966, 
         nx11618, nx11626, modgen_ram_ix167_a_160__dup_1965, 
         modgen_ram_ix167_a_161__dup_1964, modgen_ram_ix167_a_162__dup_1963, 
         nx11668, modgen_ram_ix167_a_163__dup_1962, nx11686, 
         modgen_ram_ix167_a_164__dup_1961, modgen_ram_ix167_a_165__dup_1960, 
         modgen_ram_ix167_a_166__dup_1959, modgen_ram_ix167_a_167__dup_1958, 
         nx11734, modgen_ram_ix167_a_168__dup_1957, 
         modgen_ram_ix167_a_169__dup_1956, modgen_ram_ix167_a_170__dup_1955, 
         nx11776, modgen_ram_ix167_a_171__dup_1954, nx11794, 
         modgen_ram_ix167_a_172__dup_1953, modgen_ram_ix167_a_173__dup_1952, 
         modgen_ram_ix167_a_174__dup_1951, modgen_ram_ix167_a_175__dup_1950, 
         nx11842, nx11854, modgen_ram_ix167_a_176__dup_1949, 
         modgen_ram_ix167_a_177__dup_1948, modgen_ram_ix167_a_178__dup_1947, 
         modgen_ram_ix167_a_179__dup_1946, nx11902, 
         modgen_ram_ix167_a_180__dup_1945, modgen_ram_ix167_a_181__dup_1944, 
         modgen_ram_ix167_a_182__dup_1943, modgen_ram_ix167_a_183__dup_1942, 
         nx11954, modgen_ram_ix167_a_184__dup_1941, 
         modgen_ram_ix167_a_185__dup_1940, modgen_ram_ix167_a_186__dup_1939, 
         modgen_ram_ix167_a_187__dup_1938, nx12010, 
         modgen_ram_ix167_a_188__dup_1937, modgen_ram_ix167_a_189__dup_1936, 
         modgen_ram_ix167_a_190__dup_1935, modgen_ram_ix167_a_191__dup_1934, 
         nx12062, nx12070, nx12082, modgen_ram_ix167_a_192__dup_1933, 
         modgen_ram_ix167_a_193__dup_1932, modgen_ram_ix167_a_194__dup_1931, 
         nx12116, modgen_ram_ix167_a_195__dup_1930, nx12134, 
         modgen_ram_ix167_a_196__dup_1929, modgen_ram_ix167_a_197__dup_1928, 
         modgen_ram_ix167_a_198__dup_1927, modgen_ram_ix167_a_199__dup_1926, 
         nx12182, modgen_ram_ix167_a_200__dup_1925, 
         modgen_ram_ix167_a_201__dup_1924, modgen_ram_ix167_a_202__dup_1923, 
         nx12224, modgen_ram_ix167_a_203__dup_1922, nx12242, 
         modgen_ram_ix167_a_204__dup_1921, modgen_ram_ix167_a_205__dup_1920, 
         modgen_ram_ix167_a_206__dup_1919, modgen_ram_ix167_a_207__dup_1918, 
         nx12290, nx12302, modgen_ram_ix167_a_208__dup_1917, 
         modgen_ram_ix167_a_209__dup_1916, modgen_ram_ix167_a_210__dup_1915, 
         modgen_ram_ix167_a_211__dup_1914, nx12350, 
         modgen_ram_ix167_a_212__dup_1913, modgen_ram_ix167_a_213__dup_1912, 
         modgen_ram_ix167_a_214__dup_1911, modgen_ram_ix167_a_215__dup_1910, 
         nx12402, modgen_ram_ix167_a_216__dup_1909, 
         modgen_ram_ix167_a_217__dup_1908, modgen_ram_ix167_a_218__dup_1907, 
         modgen_ram_ix167_a_219__dup_1906, nx12458, 
         modgen_ram_ix167_a_220__dup_1905, modgen_ram_ix167_a_221__dup_1904, 
         modgen_ram_ix167_a_222__dup_1903, modgen_ram_ix167_a_223__dup_1902, 
         nx12510, nx12518, modgen_ram_ix167_a_224__dup_1901, 
         modgen_ram_ix167_a_225__dup_1900, modgen_ram_ix167_a_226__dup_1899, 
         nx12560, modgen_ram_ix167_a_227__dup_1898, nx12578, 
         modgen_ram_ix167_a_228__dup_1897, modgen_ram_ix167_a_229__dup_1896, 
         modgen_ram_ix167_a_230__dup_1895, modgen_ram_ix167_a_231__dup_1894, 
         nx12626, modgen_ram_ix167_a_232__dup_1893, 
         modgen_ram_ix167_a_233__dup_1892, modgen_ram_ix167_a_234__dup_1891, 
         nx12668, modgen_ram_ix167_a_235__dup_1890, nx12686, 
         modgen_ram_ix167_a_236__dup_1889, modgen_ram_ix167_a_237__dup_1888, 
         modgen_ram_ix167_a_238__dup_1887, modgen_ram_ix167_a_239__dup_1886, 
         nx12734, nx12746, modgen_ram_ix167_a_240__dup_1885, 
         modgen_ram_ix167_a_241__dup_1884, modgen_ram_ix167_a_242__dup_1883, 
         modgen_ram_ix167_a_243__dup_1882, nx12794, 
         modgen_ram_ix167_a_244__dup_1881, modgen_ram_ix167_a_245__dup_1880, 
         modgen_ram_ix167_a_246__dup_1879, modgen_ram_ix167_a_247__dup_1878, 
         nx12846, modgen_ram_ix167_a_248__dup_1877, 
         modgen_ram_ix167_a_249__dup_1876, modgen_ram_ix167_a_250__dup_1875, 
         modgen_ram_ix167_a_251__dup_1874, nx12902, 
         modgen_ram_ix167_a_252__dup_1873, modgen_ram_ix167_a_253__dup_1872, 
         modgen_ram_ix167_a_254__dup_1871, modgen_ram_ix167_a_255__dup_1870, 
         nx12954, nx12962, nx12972, nx12986, modgen_ram_ix167_a_0__dup_1861, 
         modgen_ram_ix167_a_1__dup_1860, modgen_ram_ix167_a_2__dup_1859, nx13024, 
         modgen_ram_ix167_a_3__dup_1858, nx13042, modgen_ram_ix167_a_4__dup_1857, 
         modgen_ram_ix167_a_5__dup_1856, modgen_ram_ix167_a_6__dup_1855, 
         modgen_ram_ix167_a_7__dup_1854, nx13090, modgen_ram_ix167_a_8__dup_1853, 
         modgen_ram_ix167_a_9__dup_1852, modgen_ram_ix167_a_10__dup_1851, 
         nx13132, modgen_ram_ix167_a_11__dup_1850, nx13150, 
         modgen_ram_ix167_a_12__dup_1849, modgen_ram_ix167_a_13__dup_1848, 
         modgen_ram_ix167_a_14__dup_1847, modgen_ram_ix167_a_15__dup_1846, 
         nx13198, nx13210, modgen_ram_ix167_a_16__dup_1845, 
         modgen_ram_ix167_a_17__dup_1844, modgen_ram_ix167_a_18__dup_1843, 
         modgen_ram_ix167_a_19__dup_1842, nx13258, 
         modgen_ram_ix167_a_20__dup_1841, modgen_ram_ix167_a_21__dup_1840, 
         modgen_ram_ix167_a_22__dup_1839, modgen_ram_ix167_a_23__dup_1838, 
         nx13310, modgen_ram_ix167_a_24__dup_1837, 
         modgen_ram_ix167_a_25__dup_1836, modgen_ram_ix167_a_26__dup_1835, 
         modgen_ram_ix167_a_27__dup_1834, nx13366, 
         modgen_ram_ix167_a_28__dup_1833, modgen_ram_ix167_a_29__dup_1832, 
         modgen_ram_ix167_a_30__dup_1831, modgen_ram_ix167_a_31__dup_1830, 
         nx13418, nx13426, modgen_ram_ix167_a_32__dup_1829, 
         modgen_ram_ix167_a_33__dup_1828, modgen_ram_ix167_a_34__dup_1827, 
         nx13468, modgen_ram_ix167_a_35__dup_1826, nx13486, 
         modgen_ram_ix167_a_36__dup_1825, modgen_ram_ix167_a_37__dup_1824, 
         modgen_ram_ix167_a_38__dup_1823, modgen_ram_ix167_a_39__dup_1822, 
         nx13534, modgen_ram_ix167_a_40__dup_1821, 
         modgen_ram_ix167_a_41__dup_1820, modgen_ram_ix167_a_42__dup_1819, 
         nx13576, modgen_ram_ix167_a_43__dup_1818, nx13594, 
         modgen_ram_ix167_a_44__dup_1817, modgen_ram_ix167_a_45__dup_1816, 
         modgen_ram_ix167_a_46__dup_1815, modgen_ram_ix167_a_47__dup_1814, 
         nx13642, nx13654, modgen_ram_ix167_a_48__dup_1813, 
         modgen_ram_ix167_a_49__dup_1812, modgen_ram_ix167_a_50__dup_1811, 
         modgen_ram_ix167_a_51__dup_1810, nx13702, 
         modgen_ram_ix167_a_52__dup_1809, modgen_ram_ix167_a_53__dup_1808, 
         modgen_ram_ix167_a_54__dup_1807, modgen_ram_ix167_a_55__dup_1806, 
         nx13754, modgen_ram_ix167_a_56__dup_1805, 
         modgen_ram_ix167_a_57__dup_1804, modgen_ram_ix167_a_58__dup_1803, 
         modgen_ram_ix167_a_59__dup_1802, nx13810, 
         modgen_ram_ix167_a_60__dup_1801, modgen_ram_ix167_a_61__dup_1800, 
         modgen_ram_ix167_a_62__dup_1799, modgen_ram_ix167_a_63__dup_1798, 
         nx13862, nx13870, nx13882, modgen_ram_ix167_a_64__dup_1797, 
         modgen_ram_ix167_a_65__dup_1796, modgen_ram_ix167_a_66__dup_1795, 
         nx13916, modgen_ram_ix167_a_67__dup_1794, nx13934, 
         modgen_ram_ix167_a_68__dup_1793, modgen_ram_ix167_a_69__dup_1792, 
         modgen_ram_ix167_a_70__dup_1791, modgen_ram_ix167_a_71__dup_1790, 
         nx13982, modgen_ram_ix167_a_72__dup_1789, 
         modgen_ram_ix167_a_73__dup_1788, modgen_ram_ix167_a_74__dup_1787, 
         nx14024, modgen_ram_ix167_a_75__dup_1786, nx14042, 
         modgen_ram_ix167_a_76__dup_1785, modgen_ram_ix167_a_77__dup_1784, 
         modgen_ram_ix167_a_78__dup_1783, modgen_ram_ix167_a_79__dup_1782, 
         nx14090, nx14102, modgen_ram_ix167_a_80__dup_1781, 
         modgen_ram_ix167_a_81__dup_1780, modgen_ram_ix167_a_82__dup_1779, 
         modgen_ram_ix167_a_83__dup_1778, nx14150, 
         modgen_ram_ix167_a_84__dup_1777, modgen_ram_ix167_a_85__dup_1776, 
         modgen_ram_ix167_a_86__dup_1775, modgen_ram_ix167_a_87__dup_1774, 
         nx14202, modgen_ram_ix167_a_88__dup_1773, 
         modgen_ram_ix167_a_89__dup_1772, modgen_ram_ix167_a_90__dup_1771, 
         modgen_ram_ix167_a_91__dup_1770, nx14258, 
         modgen_ram_ix167_a_92__dup_1769, modgen_ram_ix167_a_93__dup_1768, 
         modgen_ram_ix167_a_94__dup_1767, modgen_ram_ix167_a_95__dup_1766, 
         nx14310, nx14318, modgen_ram_ix167_a_96__dup_1765, 
         modgen_ram_ix167_a_97__dup_1764, modgen_ram_ix167_a_98__dup_1763, 
         nx14360, modgen_ram_ix167_a_99__dup_1762, nx14378, 
         modgen_ram_ix167_a_100__dup_1761, modgen_ram_ix167_a_101__dup_1760, 
         modgen_ram_ix167_a_102__dup_1759, modgen_ram_ix167_a_103__dup_1758, 
         nx14426, modgen_ram_ix167_a_104__dup_1757, 
         modgen_ram_ix167_a_105__dup_1756, modgen_ram_ix167_a_106__dup_1755, 
         nx14468, modgen_ram_ix167_a_107__dup_1754, nx14486, 
         modgen_ram_ix167_a_108__dup_1753, modgen_ram_ix167_a_109__dup_1752, 
         modgen_ram_ix167_a_110__dup_1751, modgen_ram_ix167_a_111__dup_1750, 
         nx14534, nx14546, modgen_ram_ix167_a_112__dup_1749, 
         modgen_ram_ix167_a_113__dup_1748, modgen_ram_ix167_a_114__dup_1747, 
         modgen_ram_ix167_a_115__dup_1746, nx14594, 
         modgen_ram_ix167_a_116__dup_1745, modgen_ram_ix167_a_117__dup_1744, 
         modgen_ram_ix167_a_118__dup_1743, modgen_ram_ix167_a_119__dup_1742, 
         nx14646, modgen_ram_ix167_a_120__dup_1741, 
         modgen_ram_ix167_a_121__dup_1740, modgen_ram_ix167_a_122__dup_1739, 
         modgen_ram_ix167_a_123__dup_1738, nx14702, 
         modgen_ram_ix167_a_124__dup_1737, modgen_ram_ix167_a_125__dup_1736, 
         modgen_ram_ix167_a_126__dup_1735, modgen_ram_ix167_a_127__dup_1734, 
         nx14754, nx14762, nx14770, nx14778, modgen_ram_ix167_a_128__dup_1733, 
         modgen_ram_ix167_a_129__dup_1732, modgen_ram_ix167_a_130__dup_1731, 
         nx14812, modgen_ram_ix167_a_131__dup_1730, nx14830, 
         modgen_ram_ix167_a_132__dup_1729, modgen_ram_ix167_a_133__dup_1728, 
         modgen_ram_ix167_a_134__dup_1727, modgen_ram_ix167_a_135__dup_1726, 
         nx14878, modgen_ram_ix167_a_136__dup_1725, 
         modgen_ram_ix167_a_137__dup_1724, modgen_ram_ix167_a_138__dup_1723, 
         nx14920, modgen_ram_ix167_a_139__dup_1722, nx14938, 
         modgen_ram_ix167_a_140__dup_1721, modgen_ram_ix167_a_141__dup_1720, 
         modgen_ram_ix167_a_142__dup_1719, modgen_ram_ix167_a_143__dup_1718, 
         nx14986, nx14998, modgen_ram_ix167_a_144__dup_1717, 
         modgen_ram_ix167_a_145__dup_1716, modgen_ram_ix167_a_146__dup_1715, 
         modgen_ram_ix167_a_147__dup_1714, nx15046, 
         modgen_ram_ix167_a_148__dup_1713, modgen_ram_ix167_a_149__dup_1712, 
         modgen_ram_ix167_a_150__dup_1711, modgen_ram_ix167_a_151__dup_1710, 
         nx15098, modgen_ram_ix167_a_152__dup_1709, 
         modgen_ram_ix167_a_153__dup_1708, modgen_ram_ix167_a_154__dup_1707, 
         modgen_ram_ix167_a_155__dup_1706, nx15154, 
         modgen_ram_ix167_a_156__dup_1705, modgen_ram_ix167_a_157__dup_1704, 
         modgen_ram_ix167_a_158__dup_1703, modgen_ram_ix167_a_159__dup_1702, 
         nx15206, nx15214, modgen_ram_ix167_a_160__dup_1701, 
         modgen_ram_ix167_a_161__dup_1700, modgen_ram_ix167_a_162__dup_1699, 
         nx15256, modgen_ram_ix167_a_163__dup_1698, nx15274, 
         modgen_ram_ix167_a_164__dup_1697, modgen_ram_ix167_a_165__dup_1696, 
         modgen_ram_ix167_a_166__dup_1695, modgen_ram_ix167_a_167__dup_1694, 
         nx15322, modgen_ram_ix167_a_168__dup_1693, 
         modgen_ram_ix167_a_169__dup_1692, modgen_ram_ix167_a_170__dup_1691, 
         nx15364, modgen_ram_ix167_a_171__dup_1690, nx15382, 
         modgen_ram_ix167_a_172__dup_1689, modgen_ram_ix167_a_173__dup_1688, 
         modgen_ram_ix167_a_174__dup_1687, modgen_ram_ix167_a_175__dup_1686, 
         nx15430, nx15442, modgen_ram_ix167_a_176__dup_1685, 
         modgen_ram_ix167_a_177__dup_1684, modgen_ram_ix167_a_178__dup_1683, 
         modgen_ram_ix167_a_179__dup_1682, nx15490, 
         modgen_ram_ix167_a_180__dup_1681, modgen_ram_ix167_a_181__dup_1680, 
         modgen_ram_ix167_a_182__dup_1679, modgen_ram_ix167_a_183__dup_1678, 
         nx15542, modgen_ram_ix167_a_184__dup_1677, 
         modgen_ram_ix167_a_185__dup_1676, modgen_ram_ix167_a_186__dup_1675, 
         modgen_ram_ix167_a_187__dup_1674, nx15598, 
         modgen_ram_ix167_a_188__dup_1673, modgen_ram_ix167_a_189__dup_1672, 
         modgen_ram_ix167_a_190__dup_1671, modgen_ram_ix167_a_191__dup_1670, 
         nx15650, nx15658, nx15670, modgen_ram_ix167_a_192__dup_1669, 
         modgen_ram_ix167_a_193__dup_1668, modgen_ram_ix167_a_194__dup_1667, 
         nx15704, modgen_ram_ix167_a_195__dup_1666, nx15722, 
         modgen_ram_ix167_a_196__dup_1665, modgen_ram_ix167_a_197__dup_1664, 
         modgen_ram_ix167_a_198__dup_1663, modgen_ram_ix167_a_199__dup_1662, 
         nx15770, modgen_ram_ix167_a_200__dup_1661, 
         modgen_ram_ix167_a_201__dup_1660, modgen_ram_ix167_a_202__dup_1659, 
         nx15812, modgen_ram_ix167_a_203__dup_1658, nx15830, 
         modgen_ram_ix167_a_204__dup_1657, modgen_ram_ix167_a_205__dup_1656, 
         modgen_ram_ix167_a_206__dup_1655, modgen_ram_ix167_a_207__dup_1654, 
         nx15878, nx15890, modgen_ram_ix167_a_208__dup_1653, 
         modgen_ram_ix167_a_209__dup_1652, modgen_ram_ix167_a_210__dup_1651, 
         modgen_ram_ix167_a_211__dup_1650, nx15938, 
         modgen_ram_ix167_a_212__dup_1649, modgen_ram_ix167_a_213__dup_1648, 
         modgen_ram_ix167_a_214__dup_1647, modgen_ram_ix167_a_215__dup_1646, 
         nx15990, modgen_ram_ix167_a_216__dup_1645, 
         modgen_ram_ix167_a_217__dup_1644, modgen_ram_ix167_a_218__dup_1643, 
         modgen_ram_ix167_a_219__dup_1642, nx16046, 
         modgen_ram_ix167_a_220__dup_1641, modgen_ram_ix167_a_221__dup_1640, 
         modgen_ram_ix167_a_222__dup_1639, modgen_ram_ix167_a_223__dup_1638, 
         nx16098, nx16106, modgen_ram_ix167_a_224__dup_1637, 
         modgen_ram_ix167_a_225__dup_1636, modgen_ram_ix167_a_226__dup_1635, 
         nx16148, modgen_ram_ix167_a_227__dup_1634, nx16166, 
         modgen_ram_ix167_a_228__dup_1633, modgen_ram_ix167_a_229__dup_1632, 
         modgen_ram_ix167_a_230__dup_1631, modgen_ram_ix167_a_231__dup_1630, 
         nx16214, modgen_ram_ix167_a_232__dup_1629, 
         modgen_ram_ix167_a_233__dup_1628, modgen_ram_ix167_a_234__dup_1627, 
         nx16256, modgen_ram_ix167_a_235__dup_1626, nx16274, 
         modgen_ram_ix167_a_236__dup_1625, modgen_ram_ix167_a_237__dup_1624, 
         modgen_ram_ix167_a_238__dup_1623, modgen_ram_ix167_a_239__dup_1622, 
         nx16322, nx16334, modgen_ram_ix167_a_240__dup_1621, 
         modgen_ram_ix167_a_241__dup_1620, modgen_ram_ix167_a_242__dup_1619, 
         modgen_ram_ix167_a_243__dup_1618, nx16382, 
         modgen_ram_ix167_a_244__dup_1617, modgen_ram_ix167_a_245__dup_1616, 
         modgen_ram_ix167_a_246__dup_1615, modgen_ram_ix167_a_247__dup_1614, 
         nx16434, modgen_ram_ix167_a_248__dup_1613, 
         modgen_ram_ix167_a_249__dup_1612, modgen_ram_ix167_a_250__dup_1611, 
         modgen_ram_ix167_a_251__dup_1610, nx16490, 
         modgen_ram_ix167_a_252__dup_1609, modgen_ram_ix167_a_253__dup_1608, 
         modgen_ram_ix167_a_254__dup_1607, modgen_ram_ix167_a_255__dup_1606, 
         nx16542, nx16550, nx16560, nx16574, modgen_ram_ix167_a_0__dup_1597, 
         modgen_ram_ix167_a_1__dup_1596, modgen_ram_ix167_a_2__dup_1595, nx16612, 
         modgen_ram_ix167_a_3__dup_1594, nx16630, modgen_ram_ix167_a_4__dup_1593, 
         modgen_ram_ix167_a_5__dup_1592, modgen_ram_ix167_a_6__dup_1591, 
         modgen_ram_ix167_a_7__dup_1590, nx16678, modgen_ram_ix167_a_8__dup_1589, 
         modgen_ram_ix167_a_9__dup_1588, modgen_ram_ix167_a_10__dup_1587, 
         nx16720, modgen_ram_ix167_a_11__dup_1586, nx16738, 
         modgen_ram_ix167_a_12__dup_1585, modgen_ram_ix167_a_13__dup_1584, 
         modgen_ram_ix167_a_14__dup_1583, modgen_ram_ix167_a_15__dup_1582, 
         nx16786, nx16798, modgen_ram_ix167_a_16__dup_1581, 
         modgen_ram_ix167_a_17__dup_1580, modgen_ram_ix167_a_18__dup_1579, 
         modgen_ram_ix167_a_19__dup_1578, nx16846, 
         modgen_ram_ix167_a_20__dup_1577, modgen_ram_ix167_a_21__dup_1576, 
         modgen_ram_ix167_a_22__dup_1575, modgen_ram_ix167_a_23__dup_1574, 
         nx16898, modgen_ram_ix167_a_24__dup_1573, 
         modgen_ram_ix167_a_25__dup_1572, modgen_ram_ix167_a_26__dup_1571, 
         modgen_ram_ix167_a_27__dup_1570, nx16954, 
         modgen_ram_ix167_a_28__dup_1569, modgen_ram_ix167_a_29__dup_1568, 
         modgen_ram_ix167_a_30__dup_1567, modgen_ram_ix167_a_31__dup_1566, 
         nx17006, nx17014, modgen_ram_ix167_a_32__dup_1565, 
         modgen_ram_ix167_a_33__dup_1564, modgen_ram_ix167_a_34__dup_1563, 
         nx17056, modgen_ram_ix167_a_35__dup_1562, nx17074, 
         modgen_ram_ix167_a_36__dup_1561, modgen_ram_ix167_a_37__dup_1560, 
         modgen_ram_ix167_a_38__dup_1559, modgen_ram_ix167_a_39__dup_1558, 
         nx17122, modgen_ram_ix167_a_40__dup_1557, 
         modgen_ram_ix167_a_41__dup_1556, modgen_ram_ix167_a_42__dup_1555, 
         nx17164, modgen_ram_ix167_a_43__dup_1554, nx17182, 
         modgen_ram_ix167_a_44__dup_1553, modgen_ram_ix167_a_45__dup_1552, 
         modgen_ram_ix167_a_46__dup_1551, modgen_ram_ix167_a_47__dup_1550, 
         nx17230, nx17242, modgen_ram_ix167_a_48__dup_1549, 
         modgen_ram_ix167_a_49__dup_1548, modgen_ram_ix167_a_50__dup_1547, 
         modgen_ram_ix167_a_51__dup_1546, nx17290, 
         modgen_ram_ix167_a_52__dup_1545, modgen_ram_ix167_a_53__dup_1544, 
         modgen_ram_ix167_a_54__dup_1543, modgen_ram_ix167_a_55__dup_1542, 
         nx17342, modgen_ram_ix167_a_56__dup_1541, 
         modgen_ram_ix167_a_57__dup_1540, modgen_ram_ix167_a_58__dup_1539, 
         modgen_ram_ix167_a_59__dup_1538, nx17398, 
         modgen_ram_ix167_a_60__dup_1537, modgen_ram_ix167_a_61__dup_1536, 
         modgen_ram_ix167_a_62__dup_1535, modgen_ram_ix167_a_63__dup_1534, 
         nx17450, nx17458, nx17470, modgen_ram_ix167_a_64__dup_1533, 
         modgen_ram_ix167_a_65__dup_1532, modgen_ram_ix167_a_66__dup_1531, 
         nx17504, modgen_ram_ix167_a_67__dup_1530, nx17522, 
         modgen_ram_ix167_a_68__dup_1529, modgen_ram_ix167_a_69__dup_1528, 
         modgen_ram_ix167_a_70__dup_1527, modgen_ram_ix167_a_71__dup_1526, 
         nx17570, modgen_ram_ix167_a_72__dup_1525, 
         modgen_ram_ix167_a_73__dup_1524, modgen_ram_ix167_a_74__dup_1523, 
         nx17612, modgen_ram_ix167_a_75__dup_1522, nx17630, 
         modgen_ram_ix167_a_76__dup_1521, modgen_ram_ix167_a_77__dup_1520, 
         modgen_ram_ix167_a_78__dup_1519, modgen_ram_ix167_a_79__dup_1518, 
         nx17678, nx17690, modgen_ram_ix167_a_80__dup_1517, 
         modgen_ram_ix167_a_81__dup_1516, modgen_ram_ix167_a_82__dup_1515, 
         modgen_ram_ix167_a_83__dup_1514, nx17738, 
         modgen_ram_ix167_a_84__dup_1513, modgen_ram_ix167_a_85__dup_1512, 
         modgen_ram_ix167_a_86__dup_1511, modgen_ram_ix167_a_87__dup_1510, 
         nx17790, modgen_ram_ix167_a_88__dup_1509, 
         modgen_ram_ix167_a_89__dup_1508, modgen_ram_ix167_a_90__dup_1507, 
         modgen_ram_ix167_a_91__dup_1506, nx17846, 
         modgen_ram_ix167_a_92__dup_1505, modgen_ram_ix167_a_93__dup_1504, 
         modgen_ram_ix167_a_94__dup_1503, modgen_ram_ix167_a_95__dup_1502, 
         nx17898, nx17906, modgen_ram_ix167_a_96__dup_1501, 
         modgen_ram_ix167_a_97__dup_1500, modgen_ram_ix167_a_98__dup_1499, 
         nx17948, modgen_ram_ix167_a_99__dup_1498, nx17966, 
         modgen_ram_ix167_a_100__dup_1497, modgen_ram_ix167_a_101__dup_1496, 
         modgen_ram_ix167_a_102__dup_1495, modgen_ram_ix167_a_103__dup_1494, 
         nx18014, modgen_ram_ix167_a_104__dup_1493, 
         modgen_ram_ix167_a_105__dup_1492, modgen_ram_ix167_a_106__dup_1491, 
         nx18056, modgen_ram_ix167_a_107__dup_1490, nx18074, 
         modgen_ram_ix167_a_108__dup_1489, modgen_ram_ix167_a_109__dup_1488, 
         modgen_ram_ix167_a_110__dup_1487, modgen_ram_ix167_a_111__dup_1486, 
         nx18122, nx18134, modgen_ram_ix167_a_112__dup_1485, 
         modgen_ram_ix167_a_113__dup_1484, modgen_ram_ix167_a_114__dup_1483, 
         modgen_ram_ix167_a_115__dup_1482, nx18182, 
         modgen_ram_ix167_a_116__dup_1481, modgen_ram_ix167_a_117__dup_1480, 
         modgen_ram_ix167_a_118__dup_1479, modgen_ram_ix167_a_119__dup_1478, 
         nx18234, modgen_ram_ix167_a_120__dup_1477, 
         modgen_ram_ix167_a_121__dup_1476, modgen_ram_ix167_a_122__dup_1475, 
         modgen_ram_ix167_a_123__dup_1474, nx18290, 
         modgen_ram_ix167_a_124__dup_1473, modgen_ram_ix167_a_125__dup_1472, 
         modgen_ram_ix167_a_126__dup_1471, modgen_ram_ix167_a_127__dup_1470, 
         nx18342, nx18350, nx18358, nx18366, modgen_ram_ix167_a_128__dup_1469, 
         modgen_ram_ix167_a_129__dup_1468, modgen_ram_ix167_a_130__dup_1467, 
         nx18400, modgen_ram_ix167_a_131__dup_1466, nx18418, 
         modgen_ram_ix167_a_132__dup_1465, modgen_ram_ix167_a_133__dup_1464, 
         modgen_ram_ix167_a_134__dup_1463, modgen_ram_ix167_a_135__dup_1462, 
         nx18466, modgen_ram_ix167_a_136__dup_1461, 
         modgen_ram_ix167_a_137__dup_1460, modgen_ram_ix167_a_138__dup_1459, 
         nx18508, modgen_ram_ix167_a_139__dup_1458, nx18526, 
         modgen_ram_ix167_a_140__dup_1457, modgen_ram_ix167_a_141__dup_1456, 
         modgen_ram_ix167_a_142__dup_1455, modgen_ram_ix167_a_143__dup_1454, 
         nx18574, nx18586, modgen_ram_ix167_a_144__dup_1453, 
         modgen_ram_ix167_a_145__dup_1452, modgen_ram_ix167_a_146__dup_1451, 
         modgen_ram_ix167_a_147__dup_1450, nx18634, 
         modgen_ram_ix167_a_148__dup_1449, modgen_ram_ix167_a_149__dup_1448, 
         modgen_ram_ix167_a_150__dup_1447, modgen_ram_ix167_a_151__dup_1446, 
         nx18686, modgen_ram_ix167_a_152__dup_1445, 
         modgen_ram_ix167_a_153__dup_1444, modgen_ram_ix167_a_154__dup_1443, 
         modgen_ram_ix167_a_155__dup_1442, nx18742, 
         modgen_ram_ix167_a_156__dup_1441, modgen_ram_ix167_a_157__dup_1440, 
         modgen_ram_ix167_a_158__dup_1439, modgen_ram_ix167_a_159__dup_1438, 
         nx18794, nx18802, modgen_ram_ix167_a_160__dup_1437, 
         modgen_ram_ix167_a_161__dup_1436, modgen_ram_ix167_a_162__dup_1435, 
         nx18844, modgen_ram_ix167_a_163__dup_1434, nx18862, 
         modgen_ram_ix167_a_164__dup_1433, modgen_ram_ix167_a_165__dup_1432, 
         modgen_ram_ix167_a_166__dup_1431, modgen_ram_ix167_a_167__dup_1430, 
         nx18910, modgen_ram_ix167_a_168__dup_1429, 
         modgen_ram_ix167_a_169__dup_1428, modgen_ram_ix167_a_170__dup_1427, 
         nx18952, modgen_ram_ix167_a_171__dup_1426, nx18970, 
         modgen_ram_ix167_a_172__dup_1425, modgen_ram_ix167_a_173__dup_1424, 
         modgen_ram_ix167_a_174__dup_1423, modgen_ram_ix167_a_175__dup_1422, 
         nx19018, nx19030, modgen_ram_ix167_a_176__dup_1421, 
         modgen_ram_ix167_a_177__dup_1420, modgen_ram_ix167_a_178__dup_1419, 
         modgen_ram_ix167_a_179__dup_1418, nx19078, 
         modgen_ram_ix167_a_180__dup_1417, modgen_ram_ix167_a_181__dup_1416, 
         modgen_ram_ix167_a_182__dup_1415, modgen_ram_ix167_a_183__dup_1414, 
         nx19130, modgen_ram_ix167_a_184__dup_1413, 
         modgen_ram_ix167_a_185__dup_1412, modgen_ram_ix167_a_186__dup_1411, 
         modgen_ram_ix167_a_187__dup_1410, nx19186, 
         modgen_ram_ix167_a_188__dup_1409, modgen_ram_ix167_a_189__dup_1408, 
         modgen_ram_ix167_a_190__dup_1407, modgen_ram_ix167_a_191__dup_1406, 
         nx19238, nx19246, nx19258, modgen_ram_ix167_a_192__dup_1405, 
         modgen_ram_ix167_a_193__dup_1404, modgen_ram_ix167_a_194__dup_1403, 
         nx19292, modgen_ram_ix167_a_195__dup_1402, nx19310, 
         modgen_ram_ix167_a_196__dup_1401, modgen_ram_ix167_a_197__dup_1400, 
         modgen_ram_ix167_a_198__dup_1399, modgen_ram_ix167_a_199__dup_1398, 
         nx19358, modgen_ram_ix167_a_200__dup_1397, 
         modgen_ram_ix167_a_201__dup_1396, modgen_ram_ix167_a_202__dup_1395, 
         nx19400, modgen_ram_ix167_a_203__dup_1394, nx19418, 
         modgen_ram_ix167_a_204__dup_1393, modgen_ram_ix167_a_205__dup_1392, 
         modgen_ram_ix167_a_206__dup_1391, modgen_ram_ix167_a_207__dup_1390, 
         nx19466, nx19478, modgen_ram_ix167_a_208__dup_1389, 
         modgen_ram_ix167_a_209__dup_1388, modgen_ram_ix167_a_210__dup_1387, 
         modgen_ram_ix167_a_211__dup_1386, nx19526, 
         modgen_ram_ix167_a_212__dup_1385, modgen_ram_ix167_a_213__dup_1384, 
         modgen_ram_ix167_a_214__dup_1383, modgen_ram_ix167_a_215__dup_1382, 
         nx19578, modgen_ram_ix167_a_216__dup_1381, 
         modgen_ram_ix167_a_217__dup_1380, modgen_ram_ix167_a_218__dup_1379, 
         modgen_ram_ix167_a_219__dup_1378, nx19634, 
         modgen_ram_ix167_a_220__dup_1377, modgen_ram_ix167_a_221__dup_1376, 
         modgen_ram_ix167_a_222__dup_1375, modgen_ram_ix167_a_223__dup_1374, 
         nx19686, nx19694, modgen_ram_ix167_a_224__dup_1373, 
         modgen_ram_ix167_a_225__dup_1372, modgen_ram_ix167_a_226__dup_1371, 
         nx19736, modgen_ram_ix167_a_227__dup_1370, nx19754, 
         modgen_ram_ix167_a_228__dup_1369, modgen_ram_ix167_a_229__dup_1368, 
         modgen_ram_ix167_a_230__dup_1367, modgen_ram_ix167_a_231__dup_1366, 
         nx19802, modgen_ram_ix167_a_232__dup_1365, 
         modgen_ram_ix167_a_233__dup_1364, modgen_ram_ix167_a_234__dup_1363, 
         nx19844, modgen_ram_ix167_a_235__dup_1362, nx19862, 
         modgen_ram_ix167_a_236__dup_1361, modgen_ram_ix167_a_237__dup_1360, 
         modgen_ram_ix167_a_238__dup_1359, modgen_ram_ix167_a_239__dup_1358, 
         nx19910, nx19922, modgen_ram_ix167_a_240__dup_1357, 
         modgen_ram_ix167_a_241__dup_1356, modgen_ram_ix167_a_242__dup_1355, 
         modgen_ram_ix167_a_243__dup_1354, nx19970, 
         modgen_ram_ix167_a_244__dup_1353, modgen_ram_ix167_a_245__dup_1352, 
         modgen_ram_ix167_a_246__dup_1351, modgen_ram_ix167_a_247__dup_1350, 
         nx20022, modgen_ram_ix167_a_248__dup_1349, 
         modgen_ram_ix167_a_249__dup_1348, modgen_ram_ix167_a_250__dup_1347, 
         modgen_ram_ix167_a_251__dup_1346, nx20078, 
         modgen_ram_ix167_a_252__dup_1345, modgen_ram_ix167_a_253__dup_1344, 
         modgen_ram_ix167_a_254__dup_1343, modgen_ram_ix167_a_255__dup_1342, 
         nx20130, nx20138, nx20148, nx20162, modgen_ram_ix167_a_0__dup_1333, 
         modgen_ram_ix167_a_1__dup_1332, modgen_ram_ix167_a_2__dup_1331, nx20200, 
         modgen_ram_ix167_a_3__dup_1330, nx20218, modgen_ram_ix167_a_4__dup_1329, 
         modgen_ram_ix167_a_5__dup_1328, modgen_ram_ix167_a_6__dup_1327, 
         modgen_ram_ix167_a_7__dup_1326, nx20266, modgen_ram_ix167_a_8__dup_1325, 
         modgen_ram_ix167_a_9__dup_1324, modgen_ram_ix167_a_10__dup_1323, 
         nx20308, modgen_ram_ix167_a_11__dup_1322, nx20326, 
         modgen_ram_ix167_a_12__dup_1321, modgen_ram_ix167_a_13__dup_1320, 
         modgen_ram_ix167_a_14__dup_1319, modgen_ram_ix167_a_15__dup_1318, 
         nx20374, nx20386, modgen_ram_ix167_a_16__dup_1317, 
         modgen_ram_ix167_a_17__dup_1316, modgen_ram_ix167_a_18__dup_1315, 
         modgen_ram_ix167_a_19__dup_1314, nx20434, 
         modgen_ram_ix167_a_20__dup_1313, modgen_ram_ix167_a_21__dup_1312, 
         modgen_ram_ix167_a_22__dup_1311, modgen_ram_ix167_a_23__dup_1310, 
         nx20486, modgen_ram_ix167_a_24__dup_1309, 
         modgen_ram_ix167_a_25__dup_1308, modgen_ram_ix167_a_26__dup_1307, 
         modgen_ram_ix167_a_27__dup_1306, nx20542, 
         modgen_ram_ix167_a_28__dup_1305, modgen_ram_ix167_a_29__dup_1304, 
         modgen_ram_ix167_a_30__dup_1303, modgen_ram_ix167_a_31__dup_1302, 
         nx20594, nx20602, modgen_ram_ix167_a_32__dup_1301, 
         modgen_ram_ix167_a_33__dup_1300, modgen_ram_ix167_a_34__dup_1299, 
         nx20644, modgen_ram_ix167_a_35__dup_1298, nx20662, 
         modgen_ram_ix167_a_36__dup_1297, modgen_ram_ix167_a_37__dup_1296, 
         modgen_ram_ix167_a_38__dup_1295, modgen_ram_ix167_a_39__dup_1294, 
         nx20710, modgen_ram_ix167_a_40__dup_1293, 
         modgen_ram_ix167_a_41__dup_1292, modgen_ram_ix167_a_42__dup_1291, 
         nx20752, modgen_ram_ix167_a_43__dup_1290, nx20770, 
         modgen_ram_ix167_a_44__dup_1289, modgen_ram_ix167_a_45__dup_1288, 
         modgen_ram_ix167_a_46__dup_1287, modgen_ram_ix167_a_47__dup_1286, 
         nx20818, nx20830, modgen_ram_ix167_a_48__dup_1285, 
         modgen_ram_ix167_a_49__dup_1284, modgen_ram_ix167_a_50__dup_1283, 
         modgen_ram_ix167_a_51__dup_1282, nx20878, 
         modgen_ram_ix167_a_52__dup_1281, modgen_ram_ix167_a_53__dup_1280, 
         modgen_ram_ix167_a_54__dup_1279, modgen_ram_ix167_a_55__dup_1278, 
         nx20930, modgen_ram_ix167_a_56__dup_1277, 
         modgen_ram_ix167_a_57__dup_1276, modgen_ram_ix167_a_58__dup_1275, 
         modgen_ram_ix167_a_59__dup_1274, nx20986, 
         modgen_ram_ix167_a_60__dup_1273, modgen_ram_ix167_a_61__dup_1272, 
         modgen_ram_ix167_a_62__dup_1271, modgen_ram_ix167_a_63__dup_1270, 
         nx21038, nx21046, nx21058, modgen_ram_ix167_a_64__dup_1269, 
         modgen_ram_ix167_a_65__dup_1268, modgen_ram_ix167_a_66__dup_1267, 
         nx21092, modgen_ram_ix167_a_67__dup_1266, nx21110, 
         modgen_ram_ix167_a_68__dup_1265, modgen_ram_ix167_a_69__dup_1264, 
         modgen_ram_ix167_a_70__dup_1263, modgen_ram_ix167_a_71__dup_1262, 
         nx21158, modgen_ram_ix167_a_72__dup_1261, 
         modgen_ram_ix167_a_73__dup_1260, modgen_ram_ix167_a_74__dup_1259, 
         nx21200, modgen_ram_ix167_a_75__dup_1258, nx21218, 
         modgen_ram_ix167_a_76__dup_1257, modgen_ram_ix167_a_77__dup_1256, 
         modgen_ram_ix167_a_78__dup_1255, modgen_ram_ix167_a_79__dup_1254, 
         nx21266, nx21278, modgen_ram_ix167_a_80__dup_1253, 
         modgen_ram_ix167_a_81__dup_1252, modgen_ram_ix167_a_82__dup_1251, 
         modgen_ram_ix167_a_83__dup_1250, nx21326, 
         modgen_ram_ix167_a_84__dup_1249, modgen_ram_ix167_a_85__dup_1248, 
         modgen_ram_ix167_a_86__dup_1247, modgen_ram_ix167_a_87__dup_1246, 
         nx21378, modgen_ram_ix167_a_88__dup_1245, 
         modgen_ram_ix167_a_89__dup_1244, modgen_ram_ix167_a_90__dup_1243, 
         modgen_ram_ix167_a_91__dup_1242, nx21434, 
         modgen_ram_ix167_a_92__dup_1241, modgen_ram_ix167_a_93__dup_1240, 
         modgen_ram_ix167_a_94__dup_1239, modgen_ram_ix167_a_95__dup_1238, 
         nx21486, nx21494, modgen_ram_ix167_a_96__dup_1237, 
         modgen_ram_ix167_a_97__dup_1236, modgen_ram_ix167_a_98__dup_1235, 
         nx21536, modgen_ram_ix167_a_99__dup_1234, nx21554, 
         modgen_ram_ix167_a_100__dup_1233, modgen_ram_ix167_a_101__dup_1232, 
         modgen_ram_ix167_a_102__dup_1231, modgen_ram_ix167_a_103__dup_1230, 
         nx21602, modgen_ram_ix167_a_104__dup_1229, 
         modgen_ram_ix167_a_105__dup_1228, modgen_ram_ix167_a_106__dup_1227, 
         nx21644, modgen_ram_ix167_a_107__dup_1226, nx21662, 
         modgen_ram_ix167_a_108__dup_1225, modgen_ram_ix167_a_109__dup_1224, 
         modgen_ram_ix167_a_110__dup_1223, modgen_ram_ix167_a_111__dup_1222, 
         nx21710, nx21722, modgen_ram_ix167_a_112__dup_1221, 
         modgen_ram_ix167_a_113__dup_1220, modgen_ram_ix167_a_114__dup_1219, 
         modgen_ram_ix167_a_115__dup_1218, nx21770, 
         modgen_ram_ix167_a_116__dup_1217, modgen_ram_ix167_a_117__dup_1216, 
         modgen_ram_ix167_a_118__dup_1215, modgen_ram_ix167_a_119__dup_1214, 
         nx21822, modgen_ram_ix167_a_120__dup_1213, 
         modgen_ram_ix167_a_121__dup_1212, modgen_ram_ix167_a_122__dup_1211, 
         modgen_ram_ix167_a_123__dup_1210, nx21878, 
         modgen_ram_ix167_a_124__dup_1209, modgen_ram_ix167_a_125__dup_1208, 
         modgen_ram_ix167_a_126__dup_1207, modgen_ram_ix167_a_127__dup_1206, 
         nx21930, nx21938, nx21946, nx21954, modgen_ram_ix167_a_128__dup_1205, 
         modgen_ram_ix167_a_129__dup_1204, modgen_ram_ix167_a_130__dup_1203, 
         nx21988, modgen_ram_ix167_a_131__dup_1202, nx22006, 
         modgen_ram_ix167_a_132__dup_1201, modgen_ram_ix167_a_133__dup_1200, 
         modgen_ram_ix167_a_134__dup_1199, modgen_ram_ix167_a_135__dup_1198, 
         nx22054, modgen_ram_ix167_a_136__dup_1197, 
         modgen_ram_ix167_a_137__dup_1196, modgen_ram_ix167_a_138__dup_1195, 
         nx22096, modgen_ram_ix167_a_139__dup_1194, nx22114, 
         modgen_ram_ix167_a_140__dup_1193, modgen_ram_ix167_a_141__dup_1192, 
         modgen_ram_ix167_a_142__dup_1191, modgen_ram_ix167_a_143__dup_1190, 
         nx22162, nx22174, modgen_ram_ix167_a_144__dup_1189, 
         modgen_ram_ix167_a_145__dup_1188, modgen_ram_ix167_a_146__dup_1187, 
         modgen_ram_ix167_a_147__dup_1186, nx22222, 
         modgen_ram_ix167_a_148__dup_1185, modgen_ram_ix167_a_149__dup_1184, 
         modgen_ram_ix167_a_150__dup_1183, modgen_ram_ix167_a_151__dup_1182, 
         nx22274, modgen_ram_ix167_a_152__dup_1181, 
         modgen_ram_ix167_a_153__dup_1180, modgen_ram_ix167_a_154__dup_1179, 
         modgen_ram_ix167_a_155__dup_1178, nx22330, 
         modgen_ram_ix167_a_156__dup_1177, modgen_ram_ix167_a_157__dup_1176, 
         modgen_ram_ix167_a_158__dup_1175, modgen_ram_ix167_a_159__dup_1174, 
         nx22382, nx22390, modgen_ram_ix167_a_160__dup_1173, 
         modgen_ram_ix167_a_161__dup_1172, modgen_ram_ix167_a_162__dup_1171, 
         nx22432, modgen_ram_ix167_a_163__dup_1170, nx22450, 
         modgen_ram_ix167_a_164__dup_1169, modgen_ram_ix167_a_165__dup_1168, 
         modgen_ram_ix167_a_166__dup_1167, modgen_ram_ix167_a_167__dup_1166, 
         nx22498, modgen_ram_ix167_a_168__dup_1165, 
         modgen_ram_ix167_a_169__dup_1164, modgen_ram_ix167_a_170__dup_1163, 
         nx22540, modgen_ram_ix167_a_171__dup_1162, nx22558, 
         modgen_ram_ix167_a_172__dup_1161, modgen_ram_ix167_a_173__dup_1160, 
         modgen_ram_ix167_a_174__dup_1159, modgen_ram_ix167_a_175__dup_1158, 
         nx22606, nx22618, modgen_ram_ix167_a_176__dup_1157, 
         modgen_ram_ix167_a_177__dup_1156, modgen_ram_ix167_a_178__dup_1155, 
         modgen_ram_ix167_a_179__dup_1154, nx22666, 
         modgen_ram_ix167_a_180__dup_1153, modgen_ram_ix167_a_181__dup_1152, 
         modgen_ram_ix167_a_182__dup_1151, modgen_ram_ix167_a_183__dup_1150, 
         nx22718, modgen_ram_ix167_a_184__dup_1149, 
         modgen_ram_ix167_a_185__dup_1148, modgen_ram_ix167_a_186__dup_1147, 
         modgen_ram_ix167_a_187__dup_1146, nx22774, 
         modgen_ram_ix167_a_188__dup_1145, modgen_ram_ix167_a_189__dup_1144, 
         modgen_ram_ix167_a_190__dup_1143, modgen_ram_ix167_a_191__dup_1142, 
         nx22826, nx22834, nx22846, modgen_ram_ix167_a_192__dup_1141, 
         modgen_ram_ix167_a_193__dup_1140, modgen_ram_ix167_a_194__dup_1139, 
         nx22880, modgen_ram_ix167_a_195__dup_1138, nx22898, 
         modgen_ram_ix167_a_196__dup_1137, modgen_ram_ix167_a_197__dup_1136, 
         modgen_ram_ix167_a_198__dup_1135, modgen_ram_ix167_a_199__dup_1134, 
         nx22946, modgen_ram_ix167_a_200__dup_1133, 
         modgen_ram_ix167_a_201__dup_1132, modgen_ram_ix167_a_202__dup_1131, 
         nx22988, modgen_ram_ix167_a_203__dup_1130, nx23006, 
         modgen_ram_ix167_a_204__dup_1129, modgen_ram_ix167_a_205__dup_1128, 
         modgen_ram_ix167_a_206__dup_1127, modgen_ram_ix167_a_207__dup_1126, 
         nx23054, nx23066, modgen_ram_ix167_a_208__dup_1125, 
         modgen_ram_ix167_a_209__dup_1124, modgen_ram_ix167_a_210__dup_1123, 
         modgen_ram_ix167_a_211__dup_1122, nx23114, 
         modgen_ram_ix167_a_212__dup_1121, modgen_ram_ix167_a_213__dup_1120, 
         modgen_ram_ix167_a_214__dup_1119, modgen_ram_ix167_a_215__dup_1118, 
         nx23166, modgen_ram_ix167_a_216__dup_1117, 
         modgen_ram_ix167_a_217__dup_1116, modgen_ram_ix167_a_218__dup_1115, 
         modgen_ram_ix167_a_219__dup_1114, nx23222, 
         modgen_ram_ix167_a_220__dup_1113, modgen_ram_ix167_a_221__dup_1112, 
         modgen_ram_ix167_a_222__dup_1111, modgen_ram_ix167_a_223__dup_1110, 
         nx23274, nx23282, modgen_ram_ix167_a_224__dup_1109, 
         modgen_ram_ix167_a_225__dup_1108, modgen_ram_ix167_a_226__dup_1107, 
         nx23324, modgen_ram_ix167_a_227__dup_1106, nx23342, 
         modgen_ram_ix167_a_228__dup_1105, modgen_ram_ix167_a_229__dup_1104, 
         modgen_ram_ix167_a_230__dup_1103, modgen_ram_ix167_a_231__dup_1102, 
         nx23390, modgen_ram_ix167_a_232__dup_1101, 
         modgen_ram_ix167_a_233__dup_1100, modgen_ram_ix167_a_234__dup_1099, 
         nx23432, modgen_ram_ix167_a_235__dup_1098, nx23450, 
         modgen_ram_ix167_a_236__dup_1097, modgen_ram_ix167_a_237__dup_1096, 
         modgen_ram_ix167_a_238__dup_1095, modgen_ram_ix167_a_239__dup_1094, 
         nx23498, nx23510, modgen_ram_ix167_a_240__dup_1093, 
         modgen_ram_ix167_a_241__dup_1092, modgen_ram_ix167_a_242__dup_1091, 
         modgen_ram_ix167_a_243__dup_1090, nx23558, 
         modgen_ram_ix167_a_244__dup_1089, modgen_ram_ix167_a_245__dup_1088, 
         modgen_ram_ix167_a_246__dup_1087, modgen_ram_ix167_a_247__dup_1086, 
         nx23610, modgen_ram_ix167_a_248__dup_1085, 
         modgen_ram_ix167_a_249__dup_1084, modgen_ram_ix167_a_250__dup_1083, 
         modgen_ram_ix167_a_251__dup_1082, nx23666, 
         modgen_ram_ix167_a_252__dup_1081, modgen_ram_ix167_a_253__dup_1080, 
         modgen_ram_ix167_a_254__dup_1079, modgen_ram_ix167_a_255__dup_1078, 
         nx23718, nx23726, nx23736, nx23750, modgen_ram_ix167_a_0__dup_1069, 
         modgen_ram_ix167_a_1__dup_1068, modgen_ram_ix167_a_2__dup_1067, nx23788, 
         modgen_ram_ix167_a_3__dup_1066, nx23806, modgen_ram_ix167_a_4__dup_1065, 
         modgen_ram_ix167_a_5__dup_1064, modgen_ram_ix167_a_6__dup_1063, 
         modgen_ram_ix167_a_7__dup_1062, nx23854, modgen_ram_ix167_a_8__dup_1061, 
         modgen_ram_ix167_a_9__dup_1060, modgen_ram_ix167_a_10__dup_1059, 
         nx23896, modgen_ram_ix167_a_11__dup_1058, nx23914, 
         modgen_ram_ix167_a_12__dup_1057, modgen_ram_ix167_a_13__dup_1056, 
         modgen_ram_ix167_a_14__dup_1055, modgen_ram_ix167_a_15__dup_1054, 
         nx23962, nx23974, modgen_ram_ix167_a_16__dup_1053, 
         modgen_ram_ix167_a_17__dup_1052, modgen_ram_ix167_a_18__dup_1051, 
         modgen_ram_ix167_a_19__dup_1050, nx24022, 
         modgen_ram_ix167_a_20__dup_1049, modgen_ram_ix167_a_21__dup_1048, 
         modgen_ram_ix167_a_22__dup_1047, modgen_ram_ix167_a_23__dup_1046, 
         nx24074, modgen_ram_ix167_a_24__dup_1045, 
         modgen_ram_ix167_a_25__dup_1044, modgen_ram_ix167_a_26__dup_1043, 
         modgen_ram_ix167_a_27__dup_1042, nx24130, 
         modgen_ram_ix167_a_28__dup_1041, modgen_ram_ix167_a_29__dup_1040, 
         modgen_ram_ix167_a_30__dup_1039, modgen_ram_ix167_a_31__dup_1038, 
         nx24182, nx24190, modgen_ram_ix167_a_32__dup_1037, 
         modgen_ram_ix167_a_33__dup_1036, modgen_ram_ix167_a_34__dup_1035, 
         nx24232, modgen_ram_ix167_a_35__dup_1034, nx24250, 
         modgen_ram_ix167_a_36__dup_1033, modgen_ram_ix167_a_37__dup_1032, 
         modgen_ram_ix167_a_38__dup_1031, modgen_ram_ix167_a_39__dup_1030, 
         nx24298, modgen_ram_ix167_a_40__dup_1029, 
         modgen_ram_ix167_a_41__dup_1028, modgen_ram_ix167_a_42__dup_1027, 
         nx24340, modgen_ram_ix167_a_43__dup_1026, nx24358, 
         modgen_ram_ix167_a_44__dup_1025, modgen_ram_ix167_a_45__dup_1024, 
         modgen_ram_ix167_a_46__dup_1023, modgen_ram_ix167_a_47__dup_1022, 
         nx24406, nx24418, modgen_ram_ix167_a_48__dup_1021, 
         modgen_ram_ix167_a_49__dup_1020, modgen_ram_ix167_a_50__dup_1019, 
         modgen_ram_ix167_a_51__dup_1018, nx24466, 
         modgen_ram_ix167_a_52__dup_1017, modgen_ram_ix167_a_53__dup_1016, 
         modgen_ram_ix167_a_54__dup_1015, modgen_ram_ix167_a_55__dup_1014, 
         nx24518, modgen_ram_ix167_a_56__dup_1013, 
         modgen_ram_ix167_a_57__dup_1012, modgen_ram_ix167_a_58__dup_1011, 
         modgen_ram_ix167_a_59__dup_1010, nx24574, 
         modgen_ram_ix167_a_60__dup_1009, modgen_ram_ix167_a_61__dup_1008, 
         modgen_ram_ix167_a_62__dup_1007, modgen_ram_ix167_a_63__dup_1006, 
         nx24626, nx24634, nx24646, modgen_ram_ix167_a_64__dup_1005, 
         modgen_ram_ix167_a_65__dup_1004, modgen_ram_ix167_a_66__dup_1003, 
         nx24680, modgen_ram_ix167_a_67__dup_1002, nx24698, 
         modgen_ram_ix167_a_68__dup_1001, modgen_ram_ix167_a_69__dup_1000, 
         modgen_ram_ix167_a_70__dup_999, modgen_ram_ix167_a_71__dup_998, nx24746, 
         modgen_ram_ix167_a_72__dup_997, modgen_ram_ix167_a_73__dup_996, 
         modgen_ram_ix167_a_74__dup_995, nx24788, modgen_ram_ix167_a_75__dup_994, 
         nx24806, modgen_ram_ix167_a_76__dup_993, modgen_ram_ix167_a_77__dup_992, 
         modgen_ram_ix167_a_78__dup_991, modgen_ram_ix167_a_79__dup_990, nx24854, 
         nx24866, modgen_ram_ix167_a_80__dup_989, modgen_ram_ix167_a_81__dup_988, 
         modgen_ram_ix167_a_82__dup_987, modgen_ram_ix167_a_83__dup_986, nx24914, 
         modgen_ram_ix167_a_84__dup_985, modgen_ram_ix167_a_85__dup_984, 
         modgen_ram_ix167_a_86__dup_983, modgen_ram_ix167_a_87__dup_982, nx24966, 
         modgen_ram_ix167_a_88__dup_981, modgen_ram_ix167_a_89__dup_980, 
         modgen_ram_ix167_a_90__dup_979, modgen_ram_ix167_a_91__dup_978, nx25022, 
         modgen_ram_ix167_a_92__dup_977, modgen_ram_ix167_a_93__dup_976, 
         modgen_ram_ix167_a_94__dup_975, modgen_ram_ix167_a_95__dup_974, nx25074, 
         nx25082, modgen_ram_ix167_a_96__dup_973, modgen_ram_ix167_a_97__dup_972, 
         modgen_ram_ix167_a_98__dup_971, nx25124, modgen_ram_ix167_a_99__dup_970, 
         nx25142, modgen_ram_ix167_a_100__dup_969, 
         modgen_ram_ix167_a_101__dup_968, modgen_ram_ix167_a_102__dup_967, 
         modgen_ram_ix167_a_103__dup_966, nx25190, 
         modgen_ram_ix167_a_104__dup_965, modgen_ram_ix167_a_105__dup_964, 
         modgen_ram_ix167_a_106__dup_963, nx25232, 
         modgen_ram_ix167_a_107__dup_962, nx25250, 
         modgen_ram_ix167_a_108__dup_961, modgen_ram_ix167_a_109__dup_960, 
         modgen_ram_ix167_a_110__dup_959, modgen_ram_ix167_a_111__dup_958, 
         nx25298, nx25310, modgen_ram_ix167_a_112__dup_957, 
         modgen_ram_ix167_a_113__dup_956, modgen_ram_ix167_a_114__dup_955, 
         modgen_ram_ix167_a_115__dup_954, nx25358, 
         modgen_ram_ix167_a_116__dup_953, modgen_ram_ix167_a_117__dup_952, 
         modgen_ram_ix167_a_118__dup_951, modgen_ram_ix167_a_119__dup_950, 
         nx25410, modgen_ram_ix167_a_120__dup_949, 
         modgen_ram_ix167_a_121__dup_948, modgen_ram_ix167_a_122__dup_947, 
         modgen_ram_ix167_a_123__dup_946, nx25466, 
         modgen_ram_ix167_a_124__dup_945, modgen_ram_ix167_a_125__dup_944, 
         modgen_ram_ix167_a_126__dup_943, modgen_ram_ix167_a_127__dup_942, 
         nx25518, nx25526, nx25534, nx25542, modgen_ram_ix167_a_128__dup_941, 
         modgen_ram_ix167_a_129__dup_940, modgen_ram_ix167_a_130__dup_939, 
         nx25576, modgen_ram_ix167_a_131__dup_938, nx25594, 
         modgen_ram_ix167_a_132__dup_937, modgen_ram_ix167_a_133__dup_936, 
         modgen_ram_ix167_a_134__dup_935, modgen_ram_ix167_a_135__dup_934, 
         nx25642, modgen_ram_ix167_a_136__dup_933, 
         modgen_ram_ix167_a_137__dup_932, modgen_ram_ix167_a_138__dup_931, 
         nx25684, modgen_ram_ix167_a_139__dup_930, nx25702, 
         modgen_ram_ix167_a_140__dup_929, modgen_ram_ix167_a_141__dup_928, 
         modgen_ram_ix167_a_142__dup_927, modgen_ram_ix167_a_143__dup_926, 
         nx25750, nx25762, modgen_ram_ix167_a_144__dup_925, 
         modgen_ram_ix167_a_145__dup_924, modgen_ram_ix167_a_146__dup_923, 
         modgen_ram_ix167_a_147__dup_922, nx25810, 
         modgen_ram_ix167_a_148__dup_921, modgen_ram_ix167_a_149__dup_920, 
         modgen_ram_ix167_a_150__dup_919, modgen_ram_ix167_a_151__dup_918, 
         nx25862, modgen_ram_ix167_a_152__dup_917, 
         modgen_ram_ix167_a_153__dup_916, modgen_ram_ix167_a_154__dup_915, 
         modgen_ram_ix167_a_155__dup_914, nx25918, 
         modgen_ram_ix167_a_156__dup_913, modgen_ram_ix167_a_157__dup_912, 
         modgen_ram_ix167_a_158__dup_911, modgen_ram_ix167_a_159__dup_910, 
         nx25970, nx25978, modgen_ram_ix167_a_160__dup_909, 
         modgen_ram_ix167_a_161__dup_908, modgen_ram_ix167_a_162__dup_907, 
         nx26020, modgen_ram_ix167_a_163__dup_906, nx26038, 
         modgen_ram_ix167_a_164__dup_905, modgen_ram_ix167_a_165__dup_904, 
         modgen_ram_ix167_a_166__dup_903, modgen_ram_ix167_a_167__dup_902, 
         nx26086, modgen_ram_ix167_a_168__dup_901, 
         modgen_ram_ix167_a_169__dup_900, modgen_ram_ix167_a_170__dup_899, 
         nx26128, modgen_ram_ix167_a_171__dup_898, nx26146, 
         modgen_ram_ix167_a_172__dup_897, modgen_ram_ix167_a_173__dup_896, 
         modgen_ram_ix167_a_174__dup_895, modgen_ram_ix167_a_175__dup_894, 
         nx26194, nx26206, modgen_ram_ix167_a_176__dup_893, 
         modgen_ram_ix167_a_177__dup_892, modgen_ram_ix167_a_178__dup_891, 
         modgen_ram_ix167_a_179__dup_890, nx26254, 
         modgen_ram_ix167_a_180__dup_889, modgen_ram_ix167_a_181__dup_888, 
         modgen_ram_ix167_a_182__dup_887, modgen_ram_ix167_a_183__dup_886, 
         nx26306, modgen_ram_ix167_a_184__dup_885, 
         modgen_ram_ix167_a_185__dup_884, modgen_ram_ix167_a_186__dup_883, 
         modgen_ram_ix167_a_187__dup_882, nx26362, 
         modgen_ram_ix167_a_188__dup_881, modgen_ram_ix167_a_189__dup_880, 
         modgen_ram_ix167_a_190__dup_879, modgen_ram_ix167_a_191__dup_878, 
         nx26414, nx26422, nx26434, modgen_ram_ix167_a_192__dup_877, 
         modgen_ram_ix167_a_193__dup_876, modgen_ram_ix167_a_194__dup_875, 
         nx26468, modgen_ram_ix167_a_195__dup_874, nx26486, 
         modgen_ram_ix167_a_196__dup_873, modgen_ram_ix167_a_197__dup_872, 
         modgen_ram_ix167_a_198__dup_871, modgen_ram_ix167_a_199__dup_870, 
         nx26534, modgen_ram_ix167_a_200__dup_869, 
         modgen_ram_ix167_a_201__dup_868, modgen_ram_ix167_a_202__dup_867, 
         nx26576, modgen_ram_ix167_a_203__dup_866, nx26594, 
         modgen_ram_ix167_a_204__dup_865, modgen_ram_ix167_a_205__dup_864, 
         modgen_ram_ix167_a_206__dup_863, modgen_ram_ix167_a_207__dup_862, 
         nx26642, nx26654, modgen_ram_ix167_a_208__dup_861, 
         modgen_ram_ix167_a_209__dup_860, modgen_ram_ix167_a_210__dup_859, 
         modgen_ram_ix167_a_211__dup_858, nx26702, 
         modgen_ram_ix167_a_212__dup_857, modgen_ram_ix167_a_213__dup_856, 
         modgen_ram_ix167_a_214__dup_855, modgen_ram_ix167_a_215__dup_854, 
         nx26754, modgen_ram_ix167_a_216__dup_853, 
         modgen_ram_ix167_a_217__dup_852, modgen_ram_ix167_a_218__dup_851, 
         modgen_ram_ix167_a_219__dup_850, nx26810, 
         modgen_ram_ix167_a_220__dup_849, modgen_ram_ix167_a_221__dup_848, 
         modgen_ram_ix167_a_222__dup_847, modgen_ram_ix167_a_223__dup_846, 
         nx26862, nx26870, modgen_ram_ix167_a_224__dup_845, 
         modgen_ram_ix167_a_225__dup_844, modgen_ram_ix167_a_226__dup_843, 
         nx26912, modgen_ram_ix167_a_227__dup_842, nx26930, 
         modgen_ram_ix167_a_228__dup_841, modgen_ram_ix167_a_229__dup_840, 
         modgen_ram_ix167_a_230__dup_839, modgen_ram_ix167_a_231__dup_838, 
         nx26978, modgen_ram_ix167_a_232__dup_837, 
         modgen_ram_ix167_a_233__dup_836, modgen_ram_ix167_a_234__dup_835, 
         nx27020, modgen_ram_ix167_a_235__dup_834, nx27038, 
         modgen_ram_ix167_a_236__dup_833, modgen_ram_ix167_a_237__dup_832, 
         modgen_ram_ix167_a_238__dup_831, modgen_ram_ix167_a_239__dup_830, 
         nx27086, nx27098, modgen_ram_ix167_a_240__dup_829, 
         modgen_ram_ix167_a_241__dup_828, modgen_ram_ix167_a_242__dup_827, 
         modgen_ram_ix167_a_243__dup_826, nx27146, 
         modgen_ram_ix167_a_244__dup_825, modgen_ram_ix167_a_245__dup_824, 
         modgen_ram_ix167_a_246__dup_823, modgen_ram_ix167_a_247__dup_822, 
         nx27198, modgen_ram_ix167_a_248__dup_821, 
         modgen_ram_ix167_a_249__dup_820, modgen_ram_ix167_a_250__dup_819, 
         modgen_ram_ix167_a_251__dup_818, nx27254, 
         modgen_ram_ix167_a_252__dup_817, modgen_ram_ix167_a_253__dup_816, 
         modgen_ram_ix167_a_254__dup_815, modgen_ram_ix167_a_255__dup_814, 
         nx27306, nx27314, nx27324, nx27338, modgen_ram_ix167_a_0__dup_811, 
         modgen_ram_ix167_a_1__dup_810, modgen_ram_ix167_a_2__dup_809, nx27376, 
         modgen_ram_ix167_a_3__dup_808, nx27394, modgen_ram_ix167_a_4__dup_807, 
         modgen_ram_ix167_a_5__dup_806, modgen_ram_ix167_a_6__dup_805, 
         modgen_ram_ix167_a_7__dup_804, nx27442, modgen_ram_ix167_a_8, 
         modgen_ram_ix167_a_9, modgen_ram_ix167_a_10, nx27484, 
         modgen_ram_ix167_a_11, nx27502, modgen_ram_ix167_a_12, 
         modgen_ram_ix167_a_13, modgen_ram_ix167_a_14, modgen_ram_ix167_a_15, 
         nx27550, nx27562, modgen_ram_ix167_a_16, modgen_ram_ix167_a_17, 
         modgen_ram_ix167_a_18, modgen_ram_ix167_a_19, nx27610, 
         modgen_ram_ix167_a_20, modgen_ram_ix167_a_21, modgen_ram_ix167_a_22, 
         modgen_ram_ix167_a_23, nx27662, modgen_ram_ix167_a_24, 
         modgen_ram_ix167_a_25, modgen_ram_ix167_a_26, modgen_ram_ix167_a_27, 
         nx27718, modgen_ram_ix167_a_28, modgen_ram_ix167_a_29, 
         modgen_ram_ix167_a_30, modgen_ram_ix167_a_31, nx27770, nx27778, 
         modgen_ram_ix167_a_32, modgen_ram_ix167_a_33, modgen_ram_ix167_a_34, 
         nx27820, modgen_ram_ix167_a_35, nx27838, modgen_ram_ix167_a_36, 
         modgen_ram_ix167_a_37, modgen_ram_ix167_a_38, modgen_ram_ix167_a_39, 
         nx27886, modgen_ram_ix167_a_40, modgen_ram_ix167_a_41, 
         modgen_ram_ix167_a_42, nx27928, modgen_ram_ix167_a_43, nx27946, 
         modgen_ram_ix167_a_44, modgen_ram_ix167_a_45, modgen_ram_ix167_a_46, 
         modgen_ram_ix167_a_47, nx27994, nx28006, modgen_ram_ix167_a_48, 
         modgen_ram_ix167_a_49, modgen_ram_ix167_a_50, modgen_ram_ix167_a_51, 
         nx28054, modgen_ram_ix167_a_52, modgen_ram_ix167_a_53, 
         modgen_ram_ix167_a_54, modgen_ram_ix167_a_55, nx28106, 
         modgen_ram_ix167_a_56, modgen_ram_ix167_a_57, modgen_ram_ix167_a_58, 
         modgen_ram_ix167_a_59, nx28162, modgen_ram_ix167_a_60, 
         modgen_ram_ix167_a_61, modgen_ram_ix167_a_62, modgen_ram_ix167_a_63, 
         nx28214, nx28222, nx28234, modgen_ram_ix167_a_64, modgen_ram_ix167_a_65, 
         modgen_ram_ix167_a_66, nx28268, modgen_ram_ix167_a_67, nx28286, 
         modgen_ram_ix167_a_68, modgen_ram_ix167_a_69, modgen_ram_ix167_a_70, 
         modgen_ram_ix167_a_71, nx28334, modgen_ram_ix167_a_72, 
         modgen_ram_ix167_a_73, modgen_ram_ix167_a_74, nx28376, 
         modgen_ram_ix167_a_75, nx28394, modgen_ram_ix167_a_76, 
         modgen_ram_ix167_a_77, modgen_ram_ix167_a_78, modgen_ram_ix167_a_79, 
         nx28442, nx28454, modgen_ram_ix167_a_80, modgen_ram_ix167_a_81, 
         modgen_ram_ix167_a_82, modgen_ram_ix167_a_83, nx28502, 
         modgen_ram_ix167_a_84, modgen_ram_ix167_a_85, modgen_ram_ix167_a_86, 
         modgen_ram_ix167_a_87, nx28554, modgen_ram_ix167_a_88, 
         modgen_ram_ix167_a_89, modgen_ram_ix167_a_90, modgen_ram_ix167_a_91, 
         nx28610, modgen_ram_ix167_a_92, modgen_ram_ix167_a_93, 
         modgen_ram_ix167_a_94, modgen_ram_ix167_a_95, nx28662, nx28670, 
         modgen_ram_ix167_a_96, modgen_ram_ix167_a_97, modgen_ram_ix167_a_98, 
         nx28712, modgen_ram_ix167_a_99, nx28730, modgen_ram_ix167_a_100, 
         modgen_ram_ix167_a_101, modgen_ram_ix167_a_102, modgen_ram_ix167_a_103, 
         nx28778, modgen_ram_ix167_a_104, modgen_ram_ix167_a_105, 
         modgen_ram_ix167_a_106, nx28820, modgen_ram_ix167_a_107, nx28838, 
         modgen_ram_ix167_a_108, modgen_ram_ix167_a_109, modgen_ram_ix167_a_110, 
         modgen_ram_ix167_a_111, nx28886, nx28898, modgen_ram_ix167_a_112, 
         modgen_ram_ix167_a_113, modgen_ram_ix167_a_114, modgen_ram_ix167_a_115, 
         nx28946, modgen_ram_ix167_a_116, modgen_ram_ix167_a_117, 
         modgen_ram_ix167_a_118, modgen_ram_ix167_a_119, nx28998, 
         modgen_ram_ix167_a_120, modgen_ram_ix167_a_121, modgen_ram_ix167_a_122, 
         modgen_ram_ix167_a_123, nx29054, modgen_ram_ix167_a_124, 
         modgen_ram_ix167_a_125, modgen_ram_ix167_a_126, modgen_ram_ix167_a_127, 
         nx29106, nx29114, nx29122, nx29130, modgen_ram_ix167_a_128, 
         modgen_ram_ix167_a_129, modgen_ram_ix167_a_130, nx29164, 
         modgen_ram_ix167_a_131, nx29182, modgen_ram_ix167_a_132, 
         modgen_ram_ix167_a_133, modgen_ram_ix167_a_134, modgen_ram_ix167_a_135, 
         nx29230, modgen_ram_ix167_a_136, modgen_ram_ix167_a_137, 
         modgen_ram_ix167_a_138, nx29272, modgen_ram_ix167_a_139, nx29290, 
         modgen_ram_ix167_a_140, modgen_ram_ix167_a_141, modgen_ram_ix167_a_142, 
         modgen_ram_ix167_a_143, nx29338, nx29350, modgen_ram_ix167_a_144, 
         modgen_ram_ix167_a_145, modgen_ram_ix167_a_146, modgen_ram_ix167_a_147, 
         nx29398, modgen_ram_ix167_a_148, modgen_ram_ix167_a_149, 
         modgen_ram_ix167_a_150, modgen_ram_ix167_a_151, nx29450, 
         modgen_ram_ix167_a_152, modgen_ram_ix167_a_153, modgen_ram_ix167_a_154, 
         modgen_ram_ix167_a_155, nx29506, modgen_ram_ix167_a_156, 
         modgen_ram_ix167_a_157, modgen_ram_ix167_a_158, modgen_ram_ix167_a_159, 
         nx29558, nx29566, modgen_ram_ix167_a_160, modgen_ram_ix167_a_161, 
         modgen_ram_ix167_a_162, nx29608, modgen_ram_ix167_a_163, nx29626, 
         modgen_ram_ix167_a_164, modgen_ram_ix167_a_165, modgen_ram_ix167_a_166, 
         modgen_ram_ix167_a_167, nx29674, modgen_ram_ix167_a_168, 
         modgen_ram_ix167_a_169, modgen_ram_ix167_a_170, nx29716, 
         modgen_ram_ix167_a_171, nx29734, modgen_ram_ix167_a_172, 
         modgen_ram_ix167_a_173, modgen_ram_ix167_a_174, modgen_ram_ix167_a_175, 
         nx29782, nx29794, modgen_ram_ix167_a_176, modgen_ram_ix167_a_177, 
         modgen_ram_ix167_a_178, modgen_ram_ix167_a_179, nx29842, 
         modgen_ram_ix167_a_180, modgen_ram_ix167_a_181, modgen_ram_ix167_a_182, 
         modgen_ram_ix167_a_183, nx29894, modgen_ram_ix167_a_184, 
         modgen_ram_ix167_a_185, modgen_ram_ix167_a_186, modgen_ram_ix167_a_187, 
         nx29950, modgen_ram_ix167_a_188, modgen_ram_ix167_a_189, 
         modgen_ram_ix167_a_190, modgen_ram_ix167_a_191, nx30002, nx30010, 
         nx30022, modgen_ram_ix167_a_192, modgen_ram_ix167_a_193, 
         modgen_ram_ix167_a_194, nx30056, modgen_ram_ix167_a_195, nx30074, 
         modgen_ram_ix167_a_196, modgen_ram_ix167_a_197, modgen_ram_ix167_a_198, 
         modgen_ram_ix167_a_199, nx30122, modgen_ram_ix167_a_200, 
         modgen_ram_ix167_a_201, modgen_ram_ix167_a_202, nx30164, 
         modgen_ram_ix167_a_203, nx30182, modgen_ram_ix167_a_204, 
         modgen_ram_ix167_a_205, modgen_ram_ix167_a_206, modgen_ram_ix167_a_207, 
         nx30230, nx30242, modgen_ram_ix167_a_208, modgen_ram_ix167_a_209, 
         modgen_ram_ix167_a_210, modgen_ram_ix167_a_211, nx30290, 
         modgen_ram_ix167_a_212, modgen_ram_ix167_a_213, modgen_ram_ix167_a_214, 
         modgen_ram_ix167_a_215, nx30342, modgen_ram_ix167_a_216, 
         modgen_ram_ix167_a_217, modgen_ram_ix167_a_218, modgen_ram_ix167_a_219, 
         nx30398, modgen_ram_ix167_a_220, modgen_ram_ix167_a_221, 
         modgen_ram_ix167_a_222, modgen_ram_ix167_a_223, nx30450, nx30458, 
         modgen_ram_ix167_a_224, modgen_ram_ix167_a_225, modgen_ram_ix167_a_226, 
         nx30500, modgen_ram_ix167_a_227, nx30518, modgen_ram_ix167_a_228, 
         modgen_ram_ix167_a_229, modgen_ram_ix167_a_230, modgen_ram_ix167_a_231, 
         nx30566, modgen_ram_ix167_a_232, modgen_ram_ix167_a_233, 
         modgen_ram_ix167_a_234, nx30608, modgen_ram_ix167_a_235, nx30626, 
         modgen_ram_ix167_a_236, modgen_ram_ix167_a_237, modgen_ram_ix167_a_238, 
         modgen_ram_ix167_a_239, nx30674, nx30686, modgen_ram_ix167_a_240, 
         modgen_ram_ix167_a_241, modgen_ram_ix167_a_242, modgen_ram_ix167_a_243, 
         nx30734, modgen_ram_ix167_a_244, modgen_ram_ix167_a_245, 
         modgen_ram_ix167_a_246, modgen_ram_ix167_a_247, nx30786, 
         modgen_ram_ix167_a_248, modgen_ram_ix167_a_249, modgen_ram_ix167_a_250, 
         modgen_ram_ix167_a_251, nx30842, modgen_ram_ix167_a_252, 
         modgen_ram_ix167_a_253, modgen_ram_ix167_a_254, modgen_ram_ix167_a_255, 
         nx30894, nx30902, nx30912, nx30926, NOT_nx50, nx3286, nx3287, nx443, 
         nx3288, nx3289, nx3290, nx490, nx503, nx529, nx557, nx3291, nx673, 
         nx763, nx863, nx3292, nx869, nx3293, nx3294, nx886, nx889, nx3295, 
         nx3297, nx3298, nx911, nx917, nx3299, nx3300, nx928, nx3301, nx933, 
         nx3303, nx947, nx951, nx3304, nx3305, nx961, nx3307, nx967, nx3309, 
         nx3310, nx3311, nx3312, nx3313, nx3314, nx3315, nx3316, nx1011, nx3317, 
         nx1018, nx1021, nx1027, nx1029, nx1033, nx1043, nx1049, nx1051, nx3319, 
         nx3321, nx3322, nx1067, nx3323, nx1081, nx1083, nx1087, nx1093, nx1095, 
         nx1099, nx1107, nx1111, nx1113, nx1117, nx1121, nx1123, nx1127, nx1131, 
         nx1133, nx1142, nx3325, nx3326, nx3327, nx1158, nx1169, nx3328, nx3329, 
         nx1181, nx1185, nx1187, nx1191, nx1202, nx1207, nx1209, nx1213, nx1218, 
         nx1220, nx1225, nx3330, nx3331, nx3332, nx3333, nx3334, nx3335, nx3336, 
         nx1267, nx1273, nx1275, nx1279, nx1284, nx1286, nx1291, nx1295, nx3337, 
         nx1309, nx1311, nx1315, nx1321, nx1323, nx1326, nx1335, nx1339, nx1341, 
         nx1344, nx1349, nx1351, nx1357, nx1367, nx3339, nx1374, nx1377, nx1383, 
         nx1385, nx1389, nx1399, nx1405, nx1407, nx1411, nx1415, nx1417, nx1423, 
         nx1425, nx1429, nx1439, nx1445, nx1447, nx1451, nx3340, nx1458, nx1461, 
         nx3341, nx3342, nx3343, nx3345, nx3346, nx3347, nx3348, nx3349, nx3350, 
         nx3351, nx3352, nx3353, nx3354, nx3355, nx3356, nx3357, nx1545, nx1549, 
         nx1555, nx3358, nx1562, nx3359, nx1575, nx3361, nx1582, nx3362, nx3363, 
         nx3364, nx1597, nx1606, nx3365, nx1613, nx1617, nx1621, nx3366, nx3367, 
         nx3369, nx3370, nx3371, nx1648, nx3372, nx1655, nx1659, nx1669, nx1675, 
         nx1677, nx3373, nx1686, nx1688, nx3374, nx1695, nx1699, nx1709, nx1715, 
         nx1717, nx1721, nx3375, nx1729, nx3377, nx1741, nx1745, nx1747, nx1751, 
         nx1755, nx3378, nx3379, nx3380, nx1777, nx1779, nx1783, nx1789, nx3381, 
         nx3382, nx3383, nx3384, nx3385, nx3386, nx3387, nx3388, nx3389, nx3390, 
         nx3391, nx3392, nx3393, nx3394, nx3395, nx3396, nx3397, nx3398, nx3399, 
         nx3401, nx3402, nx3403, nx3404, nx3405, nx3406, nx3407, nx3408, nx3409, 
         nx3411, nx3412, nx1929, nx1939, nx3413, nx3414, nx1951, nx1955, nx1957, 
         nx3415, nx1965, nx1969, nx1979, nx1985, nx1987, nx3416, nx1996, nx1998, 
         nx3417, nx2011, nx3418, nx3419, nx3420, nx2025, nx2027, nx3421, nx2041, 
         nx2047, nx2049, nx2053, nx2057, nx3422, nx3423, nx2075, nx3424, nx3425, 
         nx3427, nx3428, nx3429, nx3430, nx3431, nx3433, nx3434, nx3435, nx3436, 
         nx3437, nx3439, nx3440, nx3441, nx3442, nx3443, nx3444, nx3445, nx3446, 
         nx3447, nx3448, nx3449, nx2181, nx2185, nx3451, nx2191, nx3452, nx2205, 
         nx3453, nx2211, nx2215, nx2219, nx2221, nx3454, nx2229, nx2233, nx3455, 
         nx2253, nx2255, nx3456, nx3457, nx2267, nx3459, nx2281, nx2285, nx2287, 
         nx2291, nx2295, nx2297, nx3460, nx2311, nx3461, nx2319, nx2323, nx2327, 
         nx2329, nx3462, nx3463, nx3464, nx2349, nx3465, nx3466, nx3467, nx3468, 
         nx3469, nx3470, nx3471, nx3473, nx3474, nx3475, nx3477, nx3478, nx3479, 
         nx3480, nx3481, nx3482, nx3483, nx3485, nx3487, nx3488, nx3489, nx3490, 
         nx2451, nx2456, nx3491, nx2461, nx3492, nx2475, nx2477, nx2480, nx2485, 
         nx2487, nx2493, nx3493, nx2498, nx2511, nx3494, nx2517, nx3495, nx2525, 
         nx2527, nx2531, nx2541, nx2545, nx2547, nx2551, nx2555, nx3497, nx3498, 
         nx2571, nx2577, nx2579, nx3499, nx3500, nx3501, nx2593, nx2605, nx2609, 
         nx2611, nx2615, nx3503, nx3504, nx2627, nx2631, nx2639, nx2645, nx3505, 
         nx3506, nx3507, nx3509, nx2661, nx2671, nx2675, nx3510, nx3511, nx2687, 
         nx2689, nx2693, nx3512, nx3513, nx3514, nx2713, nx3515, nx2720, nx2723, 
         nx2733, nx3516, nx3517, nx2742, nx2747, nx2749, nx2755, nx2757, nx2760, 
         nx2773, nx2777, nx2779, nx2783, nx2788, nx2790, nx2793, nx2803, nx2807, 
         nx2809, nx2813, nx2817, nx2819, nx2825, nx2833, nx2839, nx2841, nx2845, 
         nx2849, nx2851, nx2855, nx2865, nx2869, nx2871, nx3518, nx2879, nx2881, 
         nx2887, nx2890, nx2901, nx2905, nx2907, nx2911, nx2915, nx2917, nx2921, 
         nx2931, nx2935, nx2937, nx2941, nx2947, nx2949, nx2955, nx2969, nx2975, 
         nx2977, nx2981, nx2985, nx2987, nx2991, nx3001, nx3005, nx3007, nx3011, 
         nx3015, nx3017, NOT_nx5764, NOT_nx5746, NOT_nx5724, NOT_nx5706, 
         NOT_nx5680, NOT_nx5662, NOT_nx5640, NOT_nx5622, NOT_nx5592, NOT_nx5574, 
         NOT_nx5552, NOT_nx5534, NOT_nx5508, NOT_nx5490, NOT_nx5468, NOT_nx5450, 
         NOT_nx5414, NOT_nx5396, NOT_nx5374, NOT_nx5356, NOT_nx5330, NOT_nx5312, 
         NOT_nx5290, NOT_nx5272, NOT_nx5242, NOT_nx5224, NOT_nx5202, NOT_nx5184, 
         NOT_nx5158, NOT_nx5140, NOT_nx5118, NOT_nx5100, NOT_nx5060, NOT_nx5042, 
         NOT_nx5020, NOT_nx5002, NOT_nx4976, NOT_nx4958, NOT_nx4936, NOT_nx4918, 
         NOT_nx4888, NOT_nx4870, NOT_nx4848, NOT_nx4830, NOT_nx4804, NOT_nx4786, 
         NOT_nx4764, NOT_nx4746, NOT_nx4710, NOT_nx4692, NOT_nx4670, NOT_nx4652, 
         NOT_nx4626, NOT_nx4608, NOT_nx4586, NOT_nx4568, NOT_nx4538, NOT_nx4520, 
         NOT_nx4498, NOT_nx4480, NOT_nx4454, NOT_nx4436, NOT_nx4414, NOT_nx4396, 
         NOT_nx4346, NOT_nx4328, NOT_nx4306, NOT_nx4288, NOT_nx4262, NOT_nx4244, 
         NOT_nx4222, NOT_nx4204, NOT_nx4174, NOT_nx4156, NOT_nx4134, NOT_nx4116, 
         NOT_nx4090, NOT_nx4072, NOT_nx4050, NOT_nx4032, NOT_nx3996, NOT_nx3978, 
         NOT_nx3956, NOT_nx3938, NOT_nx3912, NOT_nx3894, NOT_nx3872, NOT_nx3854, 
         NOT_nx3824, NOT_nx3806, NOT_nx3784, NOT_nx3766, NOT_nx3740, NOT_nx3722, 
         NOT_nx3700, NOT_nx3682, NOT_nx3642, NOT_nx3624, NOT_nx3602, NOT_nx3584, 
         NOT_nx3558, NOT_nx3540, NOT_nx3518, NOT_nx3500, NOT_nx3470, NOT_nx3452, 
         NOT_nx3430, NOT_nx3412, NOT_nx3386, NOT_nx3368, NOT_nx3346, NOT_nx3328, 
         NOT_nx3292, NOT_nx3274, NOT_nx3252, NOT_nx3234, NOT_nx3208, NOT_nx3190, 
         NOT_nx3168, NOT_nx3150, NOT_nx3120, NOT_nx3102, NOT_nx3080, NOT_nx3062, 
         NOT_nx3036, NOT_nx3018, NOT_nx2996, NOT_nx2978, NOT_nx2926, NOT_nx2908, 
         NOT_nx2886, NOT_nx2868, NOT_nx2842, NOT_nx2824, NOT_nx2802, NOT_nx2784, 
         NOT_nx2754, NOT_nx2736, NOT_nx2714, NOT_nx2696, NOT_nx2670, NOT_nx2652, 
         NOT_nx2630, NOT_nx2612, NOT_nx2576, NOT_nx2558, NOT_nx2536, NOT_nx2518, 
         NOT_nx2492, NOT_nx2474, NOT_nx2452, NOT_nx2434, NOT_nx2404, NOT_nx2386, 
         NOT_nx2364, NOT_nx2346, NOT_nx2320, NOT_nx2302, NOT_nx2280, NOT_nx2262, 
         NOT_nx2222, NOT_nx2204, NOT_nx2182, NOT_nx2164, NOT_nx2138, NOT_nx2120, 
         NOT_nx2098, NOT_nx2080, NOT_nx2050, NOT_nx2032, NOT_nx2010, NOT_nx1992, 
         NOT_nx1966, NOT_nx1948, NOT_nx1926, NOT_nx1908, NOT_nx1872, NOT_nx1854, 
         NOT_nx1832, NOT_nx1814, NOT_nx1788, NOT_nx1770, NOT_nx1748, NOT_nx1730, 
         NOT_nx1700, NOT_nx1682, NOT_nx1660, NOT_nx1642, NOT_nx1616, NOT_nx1598, 
         NOT_nx1576, NOT_nx1558, NOT_nx1510, NOT_nx1492, NOT_nx1470, NOT_nx1452, 
         NOT_nx1426, NOT_nx1408, NOT_nx1386, NOT_nx1368, NOT_nx1338, NOT_nx1320, 
         NOT_nx1298, NOT_nx1280, NOT_nx1254, NOT_nx1236, NOT_nx1214, NOT_nx1196, 
         NOT_nx1154, NOT_nx1136, NOT_nx1114, NOT_nx1096, NOT_nx1070, NOT_nx1052, 
         NOT_nx1030, NOT_nx1012, NOT_nx982, NOT_nx964, NOT_nx942, NOT_nx924, 
         NOT_nx898, NOT_nx880, NOT_nx858, NOT_nx840, NOT_nx796, NOT_nx778, 
         NOT_nx756, NOT_nx738, NOT_nx712, NOT_nx694, NOT_nx672, NOT_nx654, 
         NOT_nx624, NOT_nx606, NOT_nx584, NOT_nx566, NOT_nx540, NOT_nx522, 
         NOT_nx500, NOT_nx482, NOT_nx442, NOT_nx422, NOT_nx398, NOT_nx378, 
         NOT_nx344, NOT_nx324, NOT_nx340, NOT_nx280, NOT_nx244, NOT_nx224, 
         NOT_nx200, NOT_nx180, NOT_nx148, nx3519, nx3520, NOT_nx70, nx28497, 
         nx28499, nx28501, nx28503, nx28509, nx28511, nx28513, nx28515, nx28517, 
         nx28519, nx28521, nx28523, nx3581, nx3583, nx3584, nx3585, nx3586, nx68, 
         nx3587, nx3588, nx100, nx421, nx3589, nx3590, nx422, nx3591, nx3592, 
         nx3593, nx425, nx3594, nx3595, nx3596, nx3597, nx3598, nx3599, nx3600, 
         nx3601, nx457, nx3602, nx3603, nx3604, nx3605, nx3606, nx3607, nx477, 
         nx3608, nx3609, nx3611, nx497, nx499, nx3612, nx3613, nx3614, nx3615, 
         nx3616, nx3617, nx3618, nx523, nx525, nx3619, nx3620, nx3621, nx3622, 
         nx3675, nx3676, nx38, nx3677, nx3679, nx3680, nx3681, nx3682, nx3683, 
         nx3684, nx3685, nx3686, nx3687, nx3689, nx512, nx522, nx534, nx3690, 
         nx3691, nx3692, nx3693, nx3695, nx3696, nx3697, nx3698, nx3699, nx3701, 
         nx569, nx571, nx574, nx3702, nx3703, nx3704, nx3705, nx3706, nx592, 
         nx3707, nx3708, nx600, nx604, nx606, nx3709, nx3710, nx615, 
         sp_7__dup_3799, nx3800, nx3801, nx30, nx3803, sp_6__dup_3804, 
         sp_5__dup_3805, sp_4__dup_3806, sp_3__dup_3807, sp_2__dup_3808, 
         sp_1__dup_3809, sp_0__dup_3810, pop, nx3811, nx3812, NOT_nx30, nx3813, 
         nx303, nx3814, nx305, nx3815, nx309, nx3817, nx3818, nx3819, nx3820, 
         nx3821, nx3823, nx382, nx323, nx331, nx345, nx3824, nx3825, nx355, 
         nx357, nx359, nx3826, nx3827, nx3829, nx377, nx381, nx3830, nx385, 
         nx3831, nx393, nx399, nx3832, nx405, nx407, nx3833, nx3834, nx3835, 
         nx429, nx431, nx3836, nx3837, nx441, nx3839, nx3841, nx448, nx3842, 
         nx3843, nx3844, nx465, nx3845, nx3846, nx473, nx3847, nx479, nx3849, 
         nx3850, nx486, nx3851, nx3880, nx3881, nx3883, nx3884, nx3885, nx3888, 
         nx3889, nx3890, nx3891, nx3892, nx3893, nx549, nx3895, NOT_nx158, nx652, 
         nx655, nx657, nx659, nx3896, nx3898, nx670, nx3899, nx3900, nx3901, 
         nx690, nx3902, nx3903, nx700, nx702, nx706, nx708, nx712, nx3905, nx718, 
         nx720, nx724, nx3906, nx3972, nx3973, nx3974, nx3975, nx3977, nx3978, 
         nx3979, nx3980, nx3981, nx3982, nx3983, nx3984, nx3985, nx180, nx3986, 
         nx3988, nx3989, nx404, nx3990, nx3991, nx3992, nx3993, nx3994, nx3995, 
         nx478, nx3996, nx483, nx3997, nx3998, nx493, nx3999, nx4000, nx4001, 
         nx4002, nx505, nx511, nx4003, nx521, nx4004, nx4005, nx4006, nx4008, 
         nx4009, nx4011, nx4012, nx4013, nx4014, nx4015, nx4016, nx4018, nx4203, 
         nx4205, nx16, nx4206, nx4208, nx4209, nx4211, nx92, nx4213, nx4215, 
         nx4217, nx4218, nx4219, nx4220, nx4222, nx4223, nx220, nx4224, nx248, 
         nx4225, nx4227, nx4228, nx4229, nx4231, nx4232, nx432, nx4233, nx4234, 
         nx4235, nx562, nx4236, nx4237, nx4238, nx4239, nx4241, nx4242, nx4243, 
         nx4244, nx4245, nx4247, nx1673, nx1683, nx4248, nx1703, nx1713, nx1723, 
         nx4249, nx4250, nx1753, nx4251, nx4252, nx4253, nx4254, nx4256, nx4258, 
         nx4260, nx4261, nx4262, nx4263, nx4264, nx4265, nx4266, nx4268, nx4269, 
         nx4270, nx4272, nx4274, nx4277, nx4279, nx1934, nx4280, nx4282, nx1949, 
         nx1956, nx1962, nx4284, nx1971, nx4286, nx4287, nx4289, nx1993, nx4290, 
         nx4291, nx4292, nx4293, nx4295, nx4296, nx4298, nx4300, nx4301, nx4303, 
         nx4304, nx4305, nx4307, nx4309, nx4311, nx4312, rx_done, nx4622, nx4623, 
         nx4624, nx4625, nx32, nx4627, nx4629, nx4631, nx52, nx4632, nx4634, 
         nx4635, receive, nx4636, nx4638, nx112, tx_done, nx4639, trans, nx4640, 
         nx4641, nx4643, sbuf_txd_2, sbuf_txd_1, nx4645, nx4646, nx4647, nx4648, 
         sbuf_txd_10, sbuf_txd_9, nx4650, nx4651, nx4652, nx4654, sbuf_txd_8, 
         nx4655, sbuf_txd_7, nx4656, sbuf_txd_6, sbuf_txd_5, sbuf_txd_4, 
         sbuf_txd_3, nx4658, nx4659, nx344, sbuf_txd_0, nx4660, shift_tr, 
         t1_ow_buf, nx418, smod_clk_tr, nx4661, nx4663, nx4665, tr_count_3, 
         tr_count_2, tr_count_1, tr_count_0, nx2326, nx4666, nx568, nx4668, 
         sbuf_rxd_tmp_11, nx4669, nx4671, shift_re, nx4672, smod_clk_re, nx4674, 
         nx4676, nx4677, nx636, nx4678, rx_sam_0, re_count_3, nx2331, nx644, 
         re_count_2, re_count_1, re_count_0, nx4679, nx4680, nx4681, rx_sam_1, 
         nx4682, nx4684, nx752, nx4686, nx4687, rxd_r, nx4689, sbuf_rxd_tmp_0, 
         sbuf_rxd_tmp_1, sbuf_rxd_tmp_2, sbuf_rxd_tmp_3, sbuf_rxd_tmp_4, 
         sbuf_rxd_tmp_5, sbuf_rxd_tmp_6, sbuf_rxd_tmp_7, sbuf_rxd_tmp_8, 
         sbuf_rxd_tmp_9, sbuf_rxd_tmp_10, nx4690, nx4691, nx1026, nx4693, nx4695, 
         nx4697, nx4698, NOT_nx2324, nx4700, nx4701, nx4702, nx4703, nx4705, 
         nx4706, nx4708, nx4709, nx2470, nx4711, nx4713, NOT_nx444, nx4715, 
         nx2520, nx2530, nx2540, nx4716, nx2560, nx2570, nx4717, nx4718, nx2600, 
         nx4719, nx2620, nx2630, nx4720, nx2650, nx2660, nx4722, nx2680, nx2690, 
         nx4725, nx4727, nx4728, nx4729, nx2740, nx2750, nx4730, nx4731, nx2780, 
         nx4732, nx2800, nx4733, nx4734, nx2980, nx2994, nx2998, nx3000, nx3003, 
         nx3008, nx4735, nx3012, nx3014, nx4739, nx3019, nx3024, nx3027, nx4740, 
         nx3037, nx3040, nx3046, nx3048, nx3052, nx4742, nx3057, nx3061, nx3063, 
         nx3067, nx3069, nx3081, nx3083, nx3085, nx3090, nx3094, nx3098, nx4744, 
         nx3102, nx3105, nx3110, nx3112, nx3119, nx3121, nx3123, nx3127, nx3129, 
         nx3132, nx4746, nx3136, nx3140, nx3143, nx3149, nx3151, nx4747, nx4748, 
         nx3161, nx3165, nx3167, nx3170, nx3174, nx3178, nx3180, nx3187, nx3190, 
         nx3194, nx3198, nx4750, nx4751, nx4752, nx4753, nx4754, nx4756, nx4757, 
         nx4758, nx4759, nx4760, nx4762, nx4763, nx4764, nx4765, nx4767, nx4768, 
         nx4769, nx4770, nx4772, nx4774, nx4775, nx4776, nx4778, nx4780, nx4781, 
         nx4782, nx4783, nx4784, nx4786, nx4787, nx4788, nx4789, nx4790, nx4792, 
         nx4793, nx4795, nx4796, nx4797, nx4799, nx4801, nx4803, nx4804, nx4806, 
         nx4808, nx4809, nx4810, nx4811, nx4813, nx4814, nx4815, nx4816, nx4820, 
         nx4821, nx4822, nx4824, nx4826, nx4828, nx4829, nx4831, nx4833, nx4835, 
         nx4836, nx4837, nx4839, nx4840, nx4841, nx4842, nx4843, nx4845, nx4846, 
         nx4848, nx4850, nx4851, nx5127, nx5128, nx5129, isrc_1__2, nx2822, 
         nx2823, nx2824, int_proc, nx5130, nx5131, nx5132, nx5133, nx5134, 
         nx5135, nx5136, nx108, nx5137, nx5138, nx5139, isrc_1__1, nx5140, 
         nx5141, nx5142, nx5143, nx5144, nx2829, nx5145, nx2830, nx208, nx2832, 
         isrc_1__0, nx5146, nx5147, nx5148, ie1_buff, nx5149, nx5151, nx5152, 
         nx268, nx5153, nx286, nx5154, nx310, nx324, nx5155, nx5156, nx5157, 
         nx5158, nx5159, nx366, nx2834, nx5160, nx5161, nx2835, nx5162, nx5163, 
         int_dept_0, nx2837, nx5164, isrc_0__0, int_dept_1, nx5165, nx5166, 
         nx5167, nx5168, nx5169, nx5170, nx5171, nx5172, nx5173, nx496, nx5174, 
         nx5175, nx5177, nx5178, nx5179, nx5180, nx5181, nx2840, nx5182, nx584, 
         nx5183, nx5184, nx5185, nx5186, nx626, nx5187, nx5188, nx2842, nx650, 
         tf1_buff, nx5189, nx5190, nx748, isrc_0__1, tf0_buff, nx788, nx5191, 
         nx5192, nx838, nx5193, nx5194, nx5195, nx898, nx912, nx5196, isrc_0__2, 
         ie0_buff, nx5197, nx5198, nx5199, nx5200, nx5201, int_lev_1__0, 
         int_lev_0__0, nx1054, nx5202, nx1096, nx5203, nx5204, nx5205, nx5206, 
         nx5207, nx1182, nx1186, nx5208, nx5209, nx1210, nx5210, nx5211, nx2859, 
         nx5212, nx5213, nx2889, nx2899, nx2909, nx2919, nx2929, NOT_nx2836, 
         nx2939, nx2959, nx5214, nx2979, nx2989, nx2999, nx3009, nx5215, nx3029, 
         nx3039, nx3049, nx3059, nx5216, nx3079, nx3089, nx3099, nx3109, nx5217, 
         nx5218, nx3139, NOT_nx2822, nx5219, nx3159, nx3169, nx3189, nx3199, 
         nx5220, nx5221, nx5222, nx5223, nx5224, nx5225, nx5226, nx5227, nx5228, 
         nx5229, nx5230, nx5231, nx5232, nx5233, nx5234, nx5235, nx5236, nx5237, 
         nx5238, nx5239, nx5240, nx5241, nx5242, nx5243, nx5244, nx5245, nx5246, 
         nx5247, nx5248, nx5249, nx5250, nx5251, nx5252, nx5253, nx5254, nx5255, 
         nx5257, nx5258, nx5259, nx5260, nx5261, nx5262, nx5263, nx5264, nx5265, 
         nx5266, nx5267, nx5268, nx5269, nx5270, nx5271, nx5272, nx5273, nx5274, 
         nx5275, nx5276, nx5277, nx5278, nx5279, nx5280, nx5281, nx5282, nx5283, 
         nx5284, nx5285, nx5286, nx5287, nx5288, nx5289, nx5290, nx5291, nx5292, 
         nx3523, nx3526, nx3530, nx3534, nx3537, nx3541, nx3553, nx5293, nx3567, 
         nx3569, nx3571, nx3578, nx5294, nx5295, nx5296, nx5297, nx5298, nx5299, 
         nx3628, nx3632, nx3643, nx5300, nx3660, nx3666, nx3668, nx5301, nx5659, 
         nx5660, nx5661, nx5662, nx5663, nx5664, t1_buff, nx5665, nx5666, nx5667, 
         nx5668, nx5669, nx5670, nx5671, nx156, nx5673, nx5674, nx5676, nx5678, 
         nx5679, nx5680, nx5681, nx5682, nx5683, nx5684, nx228, nx5685, nx5686, 
         nx5687, nx2169, nx5688, nx5689, nx5690, nx5691, nx5692, nx5693, nx348, 
         nx5695, nx2170, nx5696, nx5697, nx5698, nx5699, nx5700, nx5701, nx5702, 
         nx5703, nx5704, nx5705, nx5706, nx5707, t0_buff, nx586, nx5708, nx5709, 
         nx5710, nx5711, nx654, nx5712, nx672, nx5713, nx2174, nx5714, nx5715, 
         nx5716, nx732, nx5717, nx5718, nx5719, nx5720, nx764, nx5721, nx5722, 
         nx2177, nx802, nx5723, nx2178, nx5725, nx5726, nx5727, nx840, nx846, 
         nx864, nx874, nx5728, nx5729, nx5730, nx908, nx5731, nx5732, nx922, 
         nx5733, nx5734, nx5735, nx5736, nx5737, nx5738, nx5739, nx5740, nx5741, 
         nx5742, nx1036, nx2180, nx5743, nx5745, nx5746, nx5747, nx1078, nx5748, 
         nx1102, nx1112, nx1122, nx5749, nx5750, nx5751, nx5752, nx5753, nx1160, 
         nx5755, nx5756, nx1198, nx5757, nx1232, nx5758, nx5759, nx5760, nx5761, 
         tf1_0, tf1_1, nx1322, nx5762, nx5763, NOT_nx106, NOT_nx88, NOT_nx120, 
         NOT_nx680, nx5764, NOT_nx608, NOT_nx626, nx5765, nx5766, nx5767, nx5768, 
         nx2622, nx2625, nx5769, nx5770, nx2633, nx2635, nx5771, nx5772, nx5773, 
         nx2646, nx5775, nx2655, nx2657, nx5776, nx5777, nx2669, nx5779, nx5780, 
         nx5781, nx2683, nx5782, nx5783, nx5784, nx5785, nx2706, nx2708, nx5787, 
         nx2715, nx5788, nx5789, nx2727, nx5790, nx5791, nx2736, nx5792, nx2743, 
         nx5793, nx5795, nx2752, nx5797, nx5798, nx2764, nx2771, nx5799, nx2775, 
         nx5800, nx2782, nx2784, nx2786, nx2789, nx2792, nx2795, nx2797, nx2799, 
         nx2801, nx5801, nx2805, nx5802, nx2812, nx2814, nx5803, nx2821, nx5804, 
         nx2827, nx5805, nx2831, nx5806, nx2843, nx2846, nx2848, nx5807, nx2852, 
         nx2854, nx5808, nx5809, nx2860, nx2862, nx2864, nx2866, nx5811, nx2873, 
         nx2877, nx2882, nx5812, nx2888, nx5813, nx2895, nx2897, nx2902, nx5815, 
         nx5816, nx5817, nx2922, nx2926, nx2928, nx5818, nx2934, nx5819, nx5820, 
         nx5821, nx2950, nx2953, nx5822, nx2958, nx2960, nx2968, nx2972, nx5823, 
         nx5825, nx5826, nx5827, nx2997, nx5828, nx5829, nx3006, nx5830, nx5831, 
         nx3018, nx3023, nx3025, nx5832, nx3030, nx3035, nx5833, nx5835, nx3047, 
         nx5836, nx5837, nx3056, nx3060, nx3062, nx3064, nx3066, nx5838, nx3078, 
         nx5839, nx5840, nx5841, nx3087, nx3092, nx5842, nx3096, nx5843, nx3101, 
         nx3104, nx3106, nx5844, nx3113, nx5845, nx5846, nx3128, nx3133, nx3135, 
         nx5847, nx3147, nx5849, nx3153, nx3155, nx3160, nx6121, nx6122, nx6123, 
         nx6124, nx6125, nx6126, nx6127, nx6128, nx6129, nx6130, nx6131, nx70, 
         neg_trans, t2ex_r, nx6132, nx6133, nx6135, nx6136, nx6137, nx6138, 
         nx6139, nx6140, nx6141, nx6142, NOT_nx188, nx6143, nx6145, nx6146, 
         nx218, tc2_event, t2_r, nx2007, nx6147, nx6148, nx2008, nx2009, nx6149, 
         nx322, nx6150, nx6151, nx6152, nx360, nx2012, nx6153, nx6154, nx6155, 
         nx412, nx6156, nx2014, nx6157, nx6158, nx6159, nx476, nx6160, nx6161, 
         nx6162, nx6163, nx6165, nx540, nx6166, nx6167, nx2018, nx6168, nx6169, 
         nx6170, nx6171, nx6172, nx6173, nx6174, nx6175, nx6176, nx6177, nx686, 
         nx2022, nx6178, nx6179, nx6180, nx738, nx6181, nx770, nx782, nx6182, 
         nx6183, nx6184, nx6185, tf2_set, nx842, nx854, nx6186, nx6187, nx896, 
         nx6188, nx6189, nx6191, nx6192, nx6193, nx6195, nx6196, nx6197, 
         NOT_nx252, nx6198, nx6199, nx6200, nx6201, nx6202, nx6203, nx6204, 
         NOT_nx264, nx2271, nx6205, nx6206, nx6207, nx6208, nx6209, nx6210, 
         nx6211, nx6212, nx6213, nx6215, nx2473, nx6216, nx2479, nx2482, nx6217, 
         nx6218, nx2489, nx2491, nx6219, nx2501, nx2503, nx6220, nx2513, nx6221, 
         nx2518, nx6222, nx6223, nx2533, nx2535, nx6224, nx6225, nx6226, nx2553, 
         nx6227, nx6228, nx6229, nx2563, nx6230, nx2585, nx2592, nx6231, nx6232, 
         nx6233, nx6235, nx6236, nx6237, nx2616, nx2618, nx6238, nx6239, nx6240, 
         nx6241, nx2637, nx6243, nx6244, nx6245, nx6246, nx6247, nx6248, nx6249, 
         nx6251, nx2673, nx2678, nx2682, nx2685, nx6252, nx6253, nx6255, nx2705, 
         nx6256, nx6257, nx2717, nx6258, nx6259, nx2729, nx6260, nx2738, nx6261, 
         nx6262, nx6263, nx2753, nx2758, nx2762, nx2765, nx6264, nx2774, nx6265, 
         nx2781, nx6266, nx6267, nx6268, nx2798, nx6269, nx2802, nx2806, nx6270, 
         nx2811, nx6271, nx2815, nx6272, nx6273, nx6275, nx6276, nx2828, nx6277, 
         nx6278, nx6279, nx2836, nx6280, nx6281, nx6282, nx2853, nx6283, nx6284;



    assign wbi_cyc_o = wbi_stb_o ;
    assign wbd_cyc_o = wbd_stb_o ;
    TIELO_X1M_A12TS ix736 (.Y (ea_int)) ;
    TIEHI_X1M_A12TS ix734 (.Y (wbi_stb_o)) ;
    NOR2B_X0P7M_A12TS ix3 (.Y (we), .AN (wr), .B (wr_ind)) ;
    AND2_X0P5M_A12TS ix5 (.Y (pc_wr_dup_1371), .A (comp_wait), .B (pc_wr)) ;
    AOI21_X0P5M_A12TS ix11 (.Y (wr_dup_1054), .A0 (wr_addr_7), .A1 (nx747), .B0 (
                      nx749)) ;
    INV_X0P5B_A12TS ix748 (.Y (nx747), .A (wr_ind)) ;
    INV_X0P5B_A12TS ix750 (.Y (nx749), .A (wr)) ;
    OAI211_X1M_A12TS ix2367 (.Y (rmw), .A0 (nx4188), .A1 (nx4230), .B0 (nx4283)
                     , .C0 (nx4334)) ;
    AOI22_X0P5M_A12TS ix4189 (.Y (nx4188), .A0 (op_6), .A1 (nx102), .B0 (op1_n_6
                      ), .B1 (nx110)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_6 (.Q (op_6), .CK (wb_clk_i), .D (op1_n_6), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_6)) ;
    INV_X0P5B_A12TS ix4194 (.Y (nx4193), .A (state_1)) ;
    DFFSQ_X0P5M_A12TS reg_state_1 (.Q (state_1), .CK (wb_clk_i), .D (nx3887), .SN (
                      nx4221)) ;
    OAI21_X0P5M_A12TS ix3888 (.Y (nx3887), .A0 (nx4193), .A1 (nx4), .B0 (nx4198)
                      ) ;
    NOR2_X0P5A_A12TS ix806 (.Y (nx4), .A (mem_wait), .B (wait_data)) ;
    AO21A1AI2_X0P5M_A12TS ix4199 (.Y (nx4198), .A0 (state_1), .A1 (state_0), .B0 (
                          nx10), .C0 (nx4)) ;
    DFFSQ_X0P5M_A12TS reg_state_0 (.Q (state_0), .CK (wb_clk_i), .D (nx3897), .SN (
                      nx4221)) ;
    OAI21_X0P5M_A12TS ix3898 (.Y (nx3897), .A0 (nx4202), .A1 (nx4), .B0 (nx4204)
                      ) ;
    INV_X0P5B_A12TS ix4203 (.Y (nx4202), .A (state_0)) ;
    OAI211_X0P5M_A12TS ix4205 (.Y (nx4204), .A0 (nx64), .A1 (state_1), .B0 (
                       nx4202), .C0 (nx4)) ;
    AOI211_X0P5M_A12TS ix65 (.Y (nx64), .A0 (nx4207), .A1 (nx4216), .B0 (op1_n_3
                       ), .C0 (op1_n_6)) ;
    NAND3_X0P5A_A12TS ix4208 (.Y (nx4207), .A (nx48), .B (op1_n_1), .C (nx4214)
                      ) ;
    OAI31_X0P5M_A12TS ix49 (.Y (nx48), .A0 (op1_n_7), .A1 (op1_n_0), .A2 (nx4210
                      ), .B0 (nx4212)) ;
    INV_X0P5B_A12TS ix4211 (.Y (nx4210), .A (op1_n_5)) ;
    NAND3_X0P5A_A12TS ix4213 (.Y (nx4212), .A (op1_n_7), .B (op1_n_0), .C (
                      nx4210)) ;
    INV_X0P5B_A12TS ix4215 (.Y (nx4214), .A (op1_n_2)) ;
    NOR2_X0P5A_A12TS ix25 (.Y (nx24), .A (op1_n_0), .B (op1_n_1)) ;
    INV_X0P5B_A12TS ix4222 (.Y (nx4221), .A (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix807 (.Y (nx10), .A (state_1), .B (state_0)) ;
    AOI21_X0P5M_A12TS ix103 (.Y (nx102), .A0 (rd), .A1 (nx4226), .B0 (mem_wait)
                      ) ;
    NOR2_X1M_A12TS ix93 (.Y (rd), .A (wait_data), .B (NOT_nx10)) ;
    INV_X0P5B_A12TS ix4227 (.Y (nx4226), .A (wait_data)) ;
    NOR2_X0P5A_A12TS ix111 (.Y (nx110), .A (mem_wait), .B (nx98)) ;
    NAND2_X0P5A_A12TS ix99 (.Y (nx98), .A (rd), .B (nx4)) ;
    AOI32_X0P5M_A12TS ix4231 (.Y (nx4230), .A0 (nx2292), .A1 (nx756), .A2 (
                      nx4259), .B0 (nx834), .B1 (nx2304)) ;
    NOR2_X0P5A_A12TS ix2293 (.Y (nx2292), .A (op1_cur_0), .B (op1_cur_2)) ;
    INV_X0P5B_A12TS ix4241 (.Y (nx4240), .A (op_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_0 (.Q (op_0), .CK (wb_clk_i), .D (op1_n_0), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_0)) ;
    INV_X0P5B_A12TS ix4247 (.Y (nx4246), .A (op_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_2 (.Q (op_2), .CK (wb_clk_i), .D (op1_n_2), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_5 (.Q (op_5), .CK (wb_clk_i), .D (op1_n_5), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_5)) ;
    NAND2_X0P5A_A12TS ix85 (.Y (nx84), .A (nx4255), .B (nx4257)) ;
    NAND2_X0P5A_A12TS ix4256 (.Y (nx4255), .A (nx4226), .B (state_1)) ;
    NAND2_X0P5A_A12TS ix4258 (.Y (nx4257), .A (nx4226), .B (state_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_1 (.Q (op_1), .CK (wb_clk_i), .D (op1_n_1), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_1)) ;
    AOI22_X0P5M_A12TS ix4268 (.Y (nx4267), .A0 (op_4), .A1 (nx102), .B0 (op1_n_4
                      ), .B1 (nx110)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_4 (.Q (op_4), .CK (wb_clk_i), .D (op1_n_4), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_4)) ;
    NOR2_X0P5A_A12TS ix835 (.Y (nx834), .A (nx4267), .B (nx4271)) ;
    NAND2_X0P5A_A12TS ix4272 (.Y (nx4271), .A (nx4273), .B (nx4275)) ;
    AOI22_X0P5M_A12TS ix4274 (.Y (nx4273), .A0 (op_5), .A1 (nx102), .B0 (op1_n_5
                      ), .B1 (nx110)) ;
    AO1B2_X0P5M_A12TS ix2305 (.Y (nx2304), .A0N (nx4278), .B0 (op1_cur_2), .B1 (
                      nx4281)) ;
    AOI22_X0P5M_A12TS ix4279 (.Y (nx4278), .A0 (op_3), .A1 (nx102), .B0 (op1_n_3
                      ), .B1 (nx110)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_3 (.Q (op_3), .CK (wb_clk_i), .D (op1_n_3), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_3)) ;
    AOI31_X0P5M_A12TS ix4284 (.Y (nx4283), .A0 (op1_cur_2), .A1 (nx4285), .A2 (
                      nx834), .B0 (nx2360)) ;
    NOR2_X0P5A_A12TS ix4286 (.Y (nx4285), .A (nx194), .B (nx4188)) ;
    INV_X0P5B_A12TS ix4289 (.Y (nx4288), .A (op1_n_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_op_7 (.Q (op_7), .CK (wb_clk_i), .D (op1_n_7), .R (
                        wb_rst_i), .SE (NOT_nx10), .SI (op_7)) ;
    AOI31_X0P5M_A12TS ix2361 (.Y (nx2360), .A0 (nx4294), .A1 (nx4306), .A2 (
                      nx4322), .B0 (nx84)) ;
    NAND2_X0P5A_A12TS ix4295 (.Y (nx4294), .A (nx4285), .B (nx250)) ;
    NOR2_X0P5A_A12TS ix251 (.Y (nx250), .A (op1_cur_0), .B (nx4297)) ;
    NAND2_X0P5A_A12TS ix4298 (.Y (nx4297), .A (op1_cur_1), .B (nx4299)) ;
    NOR2_X0P5A_A12TS ix4300 (.Y (nx4299), .A (nx124), .B (op1_cur_2)) ;
    INV_X0P5B_A12TS ix4303 (.Y (nx4302), .A (op1_n_3)) ;
    AOI32_X0P5M_A12TS ix4307 (.Y (nx4306), .A0 (nx4308), .A1 (nx170), .A2 (
                      nx4317), .B0 (nx4267), .B1 (nx1396)) ;
    AOI22_X0P5M_A12TS ix4311 (.Y (nx4310), .A0 (op_7), .A1 (nx102), .B0 (op1_n_7
                      ), .B1 (nx110)) ;
    OA21A1OI2_X0P5M_A12TS ix4323 (.Y (nx4322), .A0 (nx2342), .A1 (nx4325), .B0 (
                          nx4285), .C0 (nx2336)) ;
    AND3_X0P5M_A12TS ix2343 (.Y (nx2342), .A (op1_cur_2), .B (nx4267), .C (
                     op1_cur_0)) ;
    NOR2_X0P5A_A12TS ix4326 (.Y (nx4325), .A (nx4278), .B (nx160)) ;
    NOR3_X0P5A_A12TS ix2337 (.Y (nx2336), .A (nx126), .B (op1_cur_0), .C (nx242)
                     ) ;
    NAND2_X0P5A_A12TS ix243 (.Y (nx242), .A (nx4332), .B (nx4308)) ;
    NOR2_X0P5A_A12TS ix4333 (.Y (nx4332), .A (nx4273), .B (nx4267)) ;
    AOI31_X0P5M_A12TS ix4335 (.Y (nx4334), .A0 (nx760), .A1 (nx194), .A2 (nx250)
                      , .B0 (nx2322)) ;
    NOR2_X0P5A_A12TS ix761 (.Y (nx760), .A (nx160), .B (nx4271)) ;
    OA21A1OI2_X0P5M_A12TS ix2323 (.Y (nx2322), .A0 (nx194), .A1 (nx4338), .B0 (
                          nx4340), .C0 (nx4271)) ;
    NAND2_X0P5A_A12TS ix4341 (.Y (nx4340), .A (op1_cur_1), .B (nx4285)) ;
    DFFSQ_X0P5M_A12TS reg_mem_act_0 (.Q (mem_act_0), .CK (wb_clk_i), .D (nx1660)
                      , .SN (nx4221)) ;
    NAND2_X0P5A_A12TS ix1661 (.Y (nx1660), .A (nx4344), .B (nx4346)) ;
    AOI211_X0P5M_A12TS ix4345 (.Y (nx4344), .A0 (nx4346), .A1 (nx4354), .B0 (
                       wait_data), .C0 (NOT_nx10)) ;
    AOI31_X0P5M_A12TS ix4347 (.Y (nx4346), .A0 (nx4332), .A1 (nx4317), .A2 (
                      nx4348), .B0 (nx4350)) ;
    NOR2_X0P5A_A12TS ix4349 (.Y (nx4348), .A (nx4310), .B (nx4188)) ;
    NOR3_X0P5A_A12TS ix4351 (.Y (nx4350), .A (nx126), .B (nx1080), .C (nx506)) ;
    NAND2_X0P5A_A12TS ix1081 (.Y (nx1080), .A (nx4348), .B (nx170)) ;
    AOI31_X0P5M_A12TS ix4355 (.Y (nx4354), .A0 (nx4308), .A1 (nx4273), .A2 (
                      nx4356), .B0 (nx1252)) ;
    NOR2_X0P5A_A12TS ix4357 (.Y (nx4356), .A (nx396), .B (nx126)) ;
    NAND2_X0P5A_A12TS ix397 (.Y (nx396), .A (op1_cur_0), .B (op1_cur_1)) ;
    OAI21_X0P5M_A12TS ix1253 (.Y (nx1252), .A0 (nx150), .A1 (nx1242), .B0 (
                      nx1240)) ;
    NAND2_X0P5A_A12TS ix151 (.Y (nx150), .A (nx4361), .B (nx4299)) ;
    NOR2_X0P5A_A12TS ix4362 (.Y (nx4361), .A (op1_cur_0), .B (op1_cur_1)) ;
    NAND2_X0P5A_A12TS ix1243 (.Y (nx1242), .A (nx4348), .B (nx4364)) ;
    NOR2_X0P5A_A12TS ix4365 (.Y (nx4364), .A (nx4273), .B (nx160)) ;
    DFFSQ_X0P5M_A12TS reg_mem_act_1 (.Q (mem_act_1), .CK (wb_clk_i), .D (nx1672)
                      , .SN (nx4221)) ;
    OAI31_X0P5M_A12TS ix1673 (.Y (nx1672), .A0 (nx126), .A1 (nx1080), .A2 (
                      nx4372), .B0 (nx4344)) ;
    AOI22_X0P5M_A12TS ix4373 (.Y (nx4372), .A0 (op_1), .A1 (nx102), .B0 (op1_n_1
                      ), .B1 (nx110)) ;
    DFFSQ_X0P5M_A12TS reg_mem_act_2 (.Q (mem_act_2), .CK (wb_clk_i), .D (nx1684)
                      , .SN (nx4221)) ;
    NAND3_X0P5A_A12TS ix1685 (.Y (nx1684), .A (nx1256), .B (nx1254), .C (nx4344)
                      ) ;
    NAND2_X0P5A_A12TS ix1257 (.Y (nx1256), .A (nx4377), .B (nx4356)) ;
    NOR2_X0P5A_A12TS ix4378 (.Y (nx4377), .A (nx234), .B (nx174)) ;
    NAND2_X0P5A_A12TS ix235 (.Y (nx234), .A (nx194), .B (nx4188)) ;
    NAND2_X0P5A_A12TS ix175 (.Y (nx174), .A (nx4273), .B (nx160)) ;
    NAND2_X0P5A_A12TS ix1255 (.Y (nx1254), .A (nx4382), .B (nx4356)) ;
    NOR2_X0P5A_A12TS ix4383 (.Y (nx4382), .A (nx234), .B (nx266)) ;
    NAND2_X0P5A_A12TS ix267 (.Y (nx266), .A (nx4273), .B (nx4267)) ;
    NAND2_X0P5A_A12TS ix425 (.Y (nx424), .A (nx4278), .B (op1_cur_2)) ;
    NAND2_X0P5A_A12TS ix495 (.Y (nx494), .A (nx4395), .B (nx4398)) ;
    NOR2_X0P5A_A12TS ix4396 (.Y (nx4395), .A (nx488), .B (nx4310)) ;
    NAND2_X0P5A_A12TS ix489 (.Y (nx488), .A (nx4273), .B (nx184)) ;
    NOR2_X0P5A_A12TS ix4399 (.Y (nx4398), .A (nx4278), .B (nx4267)) ;
    OAI21_X0P5M_A12TS ix4401 (.Y (nx4400), .A0 (nx4398), .A1 (nx4402), .B0 (
                      nx4404)) ;
    NOR2_X0P5A_A12TS ix4403 (.Y (nx4402), .A (nx506), .B (nx424)) ;
    NAND3_X0P5A_A12TS ix353 (.Y (nx352), .A (nx4299), .B (nx160), .C (nx4281)) ;
    NAND2_X0P5A_A12TS ix4416 (.Y (nx4415), .A (nx250), .B (nx406)) ;
    NOR2_X0P5A_A12TS ix407 (.Y (nx406), .A (nx196), .B (nx4273)) ;
    NAND2_X0P5A_A12TS ix197 (.Y (nx196), .A (nx4310), .B (nx4188)) ;
    NAND2_X0P5A_A12TS ix369 (.Y (nx368), .A (nx250), .B (nx4420)) ;
    NOR2_X0P5A_A12TS ix4421 (.Y (nx4420), .A (nx196), .B (nx266)) ;
    OAI211_X0P5M_A12TS ix555 (.Y (nx554), .A0 (nx532), .A1 (nx276), .B0 (nx4434)
                       , .C0 (nx4451)) ;
    NAND2_X0P5A_A12TS ix533 (.Y (nx532), .A (nx4281), .B (nx4429)) ;
    AOI211_X0P5M_A12TS ix4435 (.Y (nx4434), .A0 (nx4436), .A1 (nx4439), .B0 (
                       nx530), .C0 (nx4448)) ;
    OAI22_X0P5M_A12TS ix531 (.Y (nx530), .A0 (nx484), .A1 (nx516), .B0 (nx242), 
                      .B1 (nx4446)) ;
    NAND2_X0P5A_A12TS ix517 (.Y (nx516), .A (nx4444), .B (nx194)) ;
    NOR2_X0P5A_A12TS ix4445 (.Y (nx4444), .A (nx4273), .B (nx184)) ;
    NAND2_X0P5A_A12TS ix4447 (.Y (nx4446), .A (nx4361), .B (nx4429)) ;
    NOR2_X0P5A_A12TS ix4449 (.Y (nx4448), .A (nx516), .B (nx508)) ;
    NOR2_X0P5A_A12TS ix4457 (.Y (nx4456), .A (nx196), .B (nx174)) ;
    OAI211_X0P5M_A12TS ix693 (.Y (pc_wr_sel_0), .A0 (nx198), .A1 (nx4466), .B0 (
                       nx4468), .C0 (nx4476)) ;
    NAND2_X0P5A_A12TS ix4467 (.Y (nx4466), .A (nx4275), .B (nx250)) ;
    AOI22_X0P5M_A12TS ix4469 (.Y (nx4468), .A0 (nx4257), .A1 (nx564), .B0 (
                      nx4471), .B1 (nx4275)) ;
    NOR3_X0P5A_A12TS ix565 (.Y (nx564), .A (nx150), .B (nx196), .C (nx4273)) ;
    AOI21_X0P5M_A12TS ix4477 (.Y (nx4476), .A0 (nx4478), .A1 (nx554), .B0 (nx674
                      )) ;
    NOR2_X0P5A_A12TS ix4479 (.Y (nx4478), .A (nx4255), .B (nx78)) ;
    NOR2_X0P5A_A12TS ix675 (.Y (nx674), .A (nx4482), .B (nx4478)) ;
    NAND2_X0P5A_A12TS ix4483 (.Y (nx4482), .A (nx82), .B (nx656)) ;
    OAI22_X0P5M_A12TS ix657 (.Y (nx656), .A0 (nx4486), .A1 (nx4488), .B0 (nx4492
                      ), .B1 (nx4495)) ;
    NOR3_X0P5A_A12TS ix609 (.Y (nx608), .A (op_6), .B (mem_wait), .C (op_7)) ;
    NAND4B_X0P5M_A12TS ix4496 (.Y (nx4495), .AN (rd), .B (nx4246), .C (op_1), .D (
                       nx4240)) ;
    OAI21_X0P5M_A12TS ix711 (.Y (pc_wr_sel_1), .A0 (nx4422), .A1 (nx84), .B0 (
                      nx4498)) ;
    NAND4_X0P5A_A12TS ix571 (.Y (nx570), .A (nx4503), .B (nx494), .C (nx4390), .D (
                      nx4507)) ;
    NOR3_X0P5A_A12TS ix4504 (.Y (nx4503), .A (nx564), .B (nx420), .C (nx554)) ;
    OAI211_X0P5M_A12TS ix421 (.Y (nx420), .A0 (nx150), .A1 (nx308), .B0 (nx4415)
                       , .C0 (nx400)) ;
    NAND2_X0P5A_A12TS ix4508 (.Y (nx4507), .A (nx4317), .B (nx4285)) ;
    OAI22_X0P5M_A12TS ix723 (.Y (pc_wr_sel_2), .A0 (nx400), .A1 (nx224), .B0 (
                      nx82), .B1 (nx4511)) ;
    AO21A1AI2_X0P5M_A12TS ix4512 (.Y (nx4511), .A0 (nx4299), .A1 (nx4281), .B0 (
                          nx380), .C0 (nx4257)) ;
    NAND2_X0P5A_A12TS ix381 (.Y (nx380), .A (nx4514), .B (nx368)) ;
    OAI222_X0P5M_A12TS ix665 (.Y (pc_wr), .A0 (nx4257), .A1 (nx4482), .B0 (nx82)
                       , .B1 (nx4511), .C0 (nx224), .C1 (nx4519)) ;
    AOI211_X0P5M_A12TS ix4520 (.Y (nx4519), .A0 (eq), .A1 (nx582), .B0 (nx588), 
                       .C0 (nx420)) ;
    NOR3_X0P5A_A12TS ix589 (.Y (nx588), .A (eq), .B (nx442), .C (nx4524)) ;
    NOR3_X0P5A_A12TS ix443 (.Y (nx442), .A (nx234), .B (nx160), .C (nx4446)) ;
    NAND2_X0P5A_A12TS ix4525 (.Y (nx4524), .A (nx570), .B (nx4526)) ;
    AOI31_X0P5M_A12TS ix4527 (.Y (nx4526), .A0 (nx4317), .A1 (nx4285), .A2 (
                      nx4267), .B0 (nx216)) ;
    AOI21_X0P5M_A12TS ix217 (.Y (nx216), .A0 (nx206), .A1 (nx198), .B0 (nx150)
                      ) ;
    NAND2_X0P5A_A12TS ix207 (.Y (nx206), .A (nx4424), .B (nx4364)) ;
    NAND3_X0P5A_A12TS ix2287 (.Y (comp_sel_0), .A (nx4478), .B (nx4317), .C (
                      nx4285)) ;
    AO21A1AI2_X0P5M_A12TS ix747 (.Y (comp_sel_1), .A0 (nx4422), .A1 (nx200), .B0 (
                          nx84), .C0 (nx4533)) ;
    NAND2_X0P5A_A12TS ix201 (.Y (nx200), .A (nx4456), .B (nx4317)) ;
    OAI31_X0P5M_A12TS ix4534 (.Y (nx4533), .A0 (nx734), .A1 (nx216), .A2 (nx4538
                      ), .B0 (nx4478)) ;
    NOR2_X0P5A_A12TS ix735 (.Y (nx734), .A (nx150), .B (nx4536)) ;
    NAND2_X0P5A_A12TS ix4537 (.Y (nx4536), .A (nx4273), .B (nx4285)) ;
    NOR2_X0P5A_A12TS ix4539 (.Y (nx4538), .A (nx330), .B (nx150)) ;
    NAND2_X0P5A_A12TS ix331 (.Y (nx330), .A (nx4332), .B (nx4424)) ;
    DFFRPQ_X0P5M_A12TS reg_cy_sel_0 (.Q (cy_sel_0), .CK (wb_clk_i), .D (nx4157)
                       , .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4158 (.Y (nx4157), .A0 (nx1568), .A1 (nx4544), .A2 (
                      wait_data), .B0 (nx4563)) ;
    NAND2_X0P5A_A12TS ix1569 (.Y (nx1568), .A (nx4255), .B (nx4257)) ;
    AOI211_X0P5M_A12TS ix4545 (.Y (nx4544), .A0 (nx4546), .A1 (nx794), .B0 (
                       nx2204), .C0 (nx2192)) ;
    NOR2_X0P5A_A12TS ix4547 (.Y (nx4546), .A (nx272), .B (nx266)) ;
    OA21A1OI2_X0P5M_A12TS ix2205 (.Y (nx2204), .A0 (nx4273), .A1 (nx4294), .B0 (
                          nx4550), .C0 (nx4267)) ;
    OAI21_X0P5M_A12TS ix2193 (.Y (nx2192), .A0 (nx170), .A1 (nx4553), .B0 (
                      nx4556)) ;
    AOI222_X0P5M_A12TS ix4554 (.Y (nx4553), .A0 (nx194), .A1 (nx4398), .B0 (
                       nx4348), .B1 (nx2148), .C0 (nx4308), .C1 (nx250)) ;
    OAI21_X0P5M_A12TS ix2149 (.Y (nx2148), .A0 (op1_cur_2), .A1 (nx506), .B0 (
                      nx4278)) ;
    AOI31_X0P5M_A12TS ix4557 (.Y (nx4556), .A0 (nx2172), .A1 (op1_cur_2), .A2 (
                      nx4432), .B0 (nx2188)) ;
    OAI21_X0P5M_A12TS ix2173 (.Y (nx2172), .A0 (nx4310), .A1 (op1_cur_1), .B0 (
                      nx184)) ;
    AOI211_X0P5M_A12TS ix2189 (.Y (nx2188), .A0 (nx4560), .A1 (nx150), .B0 (
                       nx4273), .C0 (nx234)) ;
    NAND2_X0P5A_A12TS ix4564 (.Y (nx4563), .A (cy_sel_0), .B (wait_data)) ;
    SDFFRPQ_X0P5M_A12TS reg_cy_sel_1 (.Q (cy_sel_1), .CK (wb_clk_i), .D (nx2250)
                        , .R (wb_rst_i), .SE (wait_data), .SI (cy_sel_1)) ;
    OA21A1OI2_X0P5M_A12TS ix2251 (.Y (nx2250), .A0 (nx198), .A1 (nx4446), .B0 (
                          nx4567), .C0 (nx1568)) ;
    AND4_X0P5M_A12TS ix4568 (.Y (nx4567), .A (nx4569), .B (nx4574), .C (nx4582)
                     , .D (nx4588)) ;
    OAI21_X0P5M_A12TS ix4570 (.Y (nx4569), .A0 (nx4571), .A1 (nx4395), .B0 (
                      nx4398)) ;
    NOR2_X0P5A_A12TS ix4572 (.Y (nx4571), .A (nx948), .B (nx194)) ;
    NAND2_X0P5A_A12TS ix949 (.Y (nx948), .A (nx4273), .B (nx4188)) ;
    OA21A1OI2_X0P5M_A12TS ix4575 (.Y (nx4574), .A0 (nx4325), .A1 (nx4576), .B0 (
                          nx4395), .C0 (nx4578)) ;
    NOR2_X0P5A_A12TS ix4579 (.Y (nx4578), .A (nx398), .B (nx290)) ;
    NAND2_X0P5A_A12TS ix291 (.Y (nx290), .A (nx4308), .B (nx4364)) ;
    AOI222_X0P5M_A12TS ix4589 (.Y (nx4588), .A0 (nx4402), .A1 (nx4571), .B0 (
                       nx4590), .B1 (nx250), .C0 (nx4592), .C1 (nx914)) ;
    NOR2_X0P5A_A12TS ix4593 (.Y (nx4592), .A (nx272), .B (nx174)) ;
    DFFRPQ_X0P5M_A12TS reg_psw_set_0 (.Q (psw_set_0), .CK (wb_clk_i), .D (nx4137
                       ), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4138 (.Y (nx4137), .A0 (nx4597), .A1 (nx4630), .B0 (
                          wait_data), .C0 (nx4633)) ;
    AO21A1AI2_X0P5M_A12TS ix4598 (.Y (nx4597), .A0 (nx4592), .A1 (nx430), .B0 (
                          nx2098), .C0 (nx4628)) ;
    NAND4_X0P5A_A12TS ix2099 (.Y (nx2098), .A (nx4600), .B (nx4602), .C (nx4608)
                      , .D (nx4610)) ;
    OAI21_X0P5M_A12TS ix4601 (.Y (nx4600), .A0 (nx406), .A1 (nx4377), .B0 (
                      nx4436)) ;
    NOR2_X0P5A_A12TS ix4607 (.Y (nx4606), .A (nx948), .B (nx4310)) ;
    AOI22_X0P5M_A12TS ix4609 (.Y (nx4608), .A0 (nx4325), .A1 (nx4604), .B0 (
                      nx4398), .B1 (nx4606)) ;
    NOR3_X0P5A_A12TS ix4611 (.Y (nx4610), .A (nx2054), .B (nx544), .C (nx2042)
                     ) ;
    OAI22_X0P5M_A12TS ix2055 (.Y (nx2054), .A0 (nx484), .A1 (nx2046), .B0 (
                      nx4446), .B1 (nx4614)) ;
    NAND2_X0P5A_A12TS ix2047 (.Y (nx2046), .A (nx4444), .B (nx4310)) ;
    AO1B2_X0P5M_A12TS ix2043 (.Y (nx2042), .A0N (nx4621), .B0 (nx4356), .B1 (
                      nx2036)) ;
    AOI32_X0P5M_A12TS ix4622 (.Y (nx4621), .A0 (nx4317), .A1 (nx170), .A2 (
                      nx4308), .B0 (nx250), .B1 (nx318)) ;
    OAI21_X0P5M_A12TS ix319 (.Y (nx318), .A0 (nx234), .A1 (nx160), .B0 (nx306)
                      ) ;
    NAND2_X0P5A_A12TS ix307 (.Y (nx306), .A (nx4332), .B (nx4285)) ;
    OAI211_X0P5M_A12TS ix2037 (.Y (nx2036), .A0 (nx196), .A1 (nx4267), .B0 (
                       nx4626), .C0 (nx242)) ;
    NAND2_X0P5A_A12TS ix4627 (.Y (nx4626), .A (nx4348), .B (nx4273)) ;
    NAND2_X0P5A_A12TS ix4634 (.Y (nx4633), .A (psw_set_0), .B (wait_data)) ;
    DFFRPQ_X0P5M_A12TS reg_psw_set_1 (.Q (psw_set_1), .CK (wb_clk_i), .D (nx4147
                       ), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4148 (.Y (nx4147), .A0 (nx4637), .A1 (nx4390), .B0 (
                          wait_data), .C0 (nx4642)) ;
    AO21A1AI2_X0P5M_A12TS ix4638 (.Y (nx4637), .A0 (nx4377), .A1 (nx430), .B0 (
                          nx2120), .C0 (nx4275)) ;
    NAND2_X0P5A_A12TS ix4643 (.Y (nx4642), .A (psw_set_1), .B (wait_data)) ;
    DFFRPQ_X0P5M_A12TS reg_alu_op_0 (.Q (alu_op_0__dup_838), .CK (wb_clk_i), .D (
                       nx4047), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4650 (.Y (nx4649), .A0 (nx1408), .A1 (nx1388), .A2 (
                      nx1372), .B0 (nx4226)) ;
    OAI211_X0P5M_A12TS ix1409 (.Y (nx1408), .A0 (nx434), .A1 (nx4275), .B0 (
                       nx4653), .C0 (nx4657)) ;
    AOI32_X0P5M_A12TS ix4654 (.Y (nx4653), .A0 (nx756), .A1 (nx126), .A2 (nx4285
                      ), .B0 (nx804), .B1 (nx1214)) ;
    NOR2_X0P5A_A12TS ix805 (.Y (nx804), .A (nx4273), .B (nx84)) ;
    NOR2_X0P5A_A12TS ix1215 (.Y (nx1214), .A (nx4299), .B (nx196)) ;
    AOI22_X0P5M_A12TS ix4658 (.Y (nx4657), .A0 (nx756), .A1 (nx1396), .B0 (nx870
                      ), .B1 (nx1196)) ;
    NOR2_X0P5A_A12TS ix871 (.Y (nx870), .A (nx160), .B (nx234)) ;
    NOR2_X0P5A_A12TS ix1197 (.Y (nx1196), .A (nx84), .B (nx4560)) ;
    OAI22_X0P5M_A12TS ix1389 (.Y (nx1388), .A0 (nx4662), .A1 (nx4664), .B0 (
                      nx4188), .B1 (nx4667)) ;
    AOI32_X0P5M_A12TS ix4668 (.Y (nx4667), .A0 (nx756), .A1 (nx4429), .A2 (nx346
                      ), .B0 (nx126), .B1 (nx760)) ;
    OAI211_X0P5M_A12TS ix1373 (.Y (nx1372), .A0 (nx4297), .A1 (nx4670), .B0 (
                       nx4673), .C0 (nx4675)) ;
    AOI22_X0P5M_A12TS ix4671 (.Y (nx4670), .A0 (nx4285), .A1 (nx820), .B0 (
                      nx4308), .B1 (nx760)) ;
    NOR2_X0P5A_A12TS ix821 (.Y (nx820), .A (nx4267), .B (nx84)) ;
    NAND3_X0P5A_A12TS ix4676 (.Y (nx4675), .A (nx1356), .B (nx4267), .C (nx804)
                      ) ;
    NOR2_X0P5A_A12TS ix1357 (.Y (nx1356), .A (nx184), .B (nx4446)) ;
    DFFRPQ_X0P5M_A12TS reg_alu_op_1 (.Q (alu_op_1__dup_839), .CK (wb_clk_i), .D (
                       nx4057), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4058 (.Y (nx4057), .A0 (nx4683), .A1 (nx4696), .B0 (
                          wait_data), .C0 (nx4714)) ;
    AOI211_X0P5M_A12TS ix4684 (.Y (nx4683), .A0 (nx4685), .A1 (nx84), .B0 (
                       nx1484), .C0 (nx1472)) ;
    NOR2_X0P5A_A12TS ix4686 (.Y (nx4685), .A (nx4446), .B (nx290)) ;
    OAI21_X0P5M_A12TS ix1485 (.Y (nx1484), .A0 (nx4662), .A1 (nx4340), .B0 (
                      nx4688)) ;
    AOI32_X0P5M_A12TS ix4689 (.Y (nx4688), .A0 (nx870), .A1 (nx250), .A2 (nx756)
                      , .B0 (nx124), .B1 (nx784)) ;
    OAI22_X0P5M_A12TS ix1473 (.Y (nx1472), .A0 (nx4271), .A1 (nx4692), .B0 (
                      nx4560), .B1 (nx4694)) ;
    NAND2_X0P5A_A12TS ix4695 (.Y (nx4694), .A (nx804), .B (nx4424)) ;
    AOI221_X0P5M_A12TS ix4697 (.Y (nx4696), .A0 (nx834), .A1 (nx796), .B0 (
                       op1_cur_2), .B1 (nx1454), .C0 (nx1444)) ;
    NAND2_X0P5A_A12TS ix797 (.Y (nx796), .A (nx4699), .B (nx4278)) ;
    OAI21_X0P5M_A12TS ix4700 (.Y (nx4699), .A0 (op1_cur_0), .A1 (op1_cur_1), .B0 (
                      op1_cur_2)) ;
    NAND2_X0P5A_A12TS ix4705 (.Y (nx4704), .A (nx4310), .B (nx834)) ;
    OAI22_X0P5M_A12TS ix1445 (.Y (nx1444), .A0 (nx234), .A1 (nx4707), .B0 (
                      nx4710), .B1 (nx4712)) ;
    AOI22_X0P5M_A12TS ix4708 (.Y (nx4707), .A0 (op1_cur_1), .A1 (nx806), .B0 (
                      nx126), .B1 (nx820)) ;
    AOI32_X0P5M_A12TS ix4713 (.Y (nx4712), .A0 (nx870), .A1 (nx4278), .A2 (
                      nx4361), .B0 (nx194), .B1 (nx430)) ;
    NAND2_X0P5A_A12TS ix4715 (.Y (nx4714), .A (alu_op_1__dup_839), .B (wait_data
                      )) ;
    SDFFRPQ_X0P5M_A12TS reg_alu_op_2 (.Q (alu_op_2__dup_840), .CK (wb_clk_i), .D (
                        nx1556), .R (wb_rst_i), .SE (wait_data), .SI (
                        alu_op_2__dup_840)) ;
    NAND4B_X0P5M_A12TS ix1557 (.Y (nx1556), .AN (nx1484), .B (nx4721), .C (
                       nx4723), .D (nx4726)) ;
    AOI32_X0P5M_A12TS ix4722 (.Y (nx4721), .A0 (nx126), .A1 (nx4310), .A2 (nx834
                      ), .B0 (nx760), .B1 (nx1356)) ;
    AO21A1AI2_X0P5M_A12TS ix4724 (.Y (nx4723), .A0 (nx794), .A1 (nx4348), .B0 (
                          nx1540), .C0 (nx756)) ;
    AOI21_X0P5M_A12TS ix1541 (.Y (nx1540), .A0 (nx396), .A1 (nx4299), .B0 (nx196
                      )) ;
    AOI32_X0P5M_A12TS ix4727 (.Y (nx4726), .A0 (nx1510), .A1 (nx4308), .A2 (
                      nx806), .B0 (nx430), .B1 (nx1526)) ;
    OAI21_X0P5M_A12TS ix1511 (.Y (nx1510), .A0 (op1_cur_0), .A1 (nx126), .B0 (
                      nx4297)) ;
    DFFRPQ_X0P5M_A12TS reg_alu_op_3 (.Q (alu_op_3__dup_841), .CK (wb_clk_i), .D (
                       nx4077), .R (wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix4738 (.Y (nx4737), .A0 (nx1620), .A1 (nx1596), .B0 (
                       nx4628), .C0 (nx4226)) ;
    OAI221_X0P5M_A12TS ix1621 (.Y (nx1620), .A0 (nx4273), .A1 (nx4294), .B0 (
                       nx196), .B1 (nx4560), .C0 (nx4306)) ;
    OAI211_X0P5M_A12TS ix1597 (.Y (nx1596), .A0 (nx266), .A1 (nx4741), .B0 (
                       nx4743), .C0 (nx4745)) ;
    NAND2_X0P5A_A12TS ix4742 (.Y (nx4741), .A (nx184), .B (op1_cur_2)) ;
    NAND3_X0P5A_A12TS ix4744 (.Y (nx4743), .A (nx4285), .B (nx4267), .C (nx126)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix4746 (.Y (nx4745), .A0 (nx4348), .A1 (nx796), .B0 (
                          nx1214), .C0 (nx4273)) ;
    DFFRPQ_X0P5M_A12TS reg_src_sel3 (.Q (src_sel3), .CK (wb_clk_i), .D (nx4177)
                       , .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix4178 (.Y (nx4177), .A0N (nx4749), .B0 (src_sel3), .B1 (
                      wait_data)) ;
    AO21A1AI2_X0P5M_A12TS ix4750 (.Y (nx4749), .A0 (nx4628), .A1 (nx2272), .B0 (
                          nx1932), .C0 (nx4226)) ;
    NAND4_X0P5A_A12TS ix2273 (.Y (nx2272), .A (nx4507), .B (nx332), .C (nx4755)
                      , .D (nx4526)) ;
    AOI32_X0P5M_A12TS ix4756 (.Y (nx4755), .A0 (nx282), .A1 (op1_cur_1), .A2 (
                      nx4299), .B0 (nx4317), .B1 (nx4382)) ;
    OA21A1OI2_X0P5M_A12TS ix1933 (.Y (nx1932), .A0 (nx1242), .A1 (nx4446), .B0 (
                          nx1254), .C0 (nx1568)) ;
    DFFRPQ_X0P5M_A12TS reg_src_sel2_0 (.Q (src_sel2_0), .CK (wb_clk_i), .D (
                       nx4117), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix4118 (.Y (nx4117), .A0N (nx4761), .B0 (src_sel2_0), .B1 (
                      wait_data)) ;
    OAI31_X0P5M_A12TS ix4762 (.Y (nx4761), .A0 (nx1952), .A1 (nx1932), .A2 (
                      nx1920), .B0 (nx4226)) ;
    OA21A1OI2_X0P5M_A12TS ix1953 (.Y (nx1952), .A0 (nx264), .A1 (nx4446), .B0 (
                          nx4400), .C0 (nx1568)) ;
    AO21A1AI2_X0P5M_A12TS ix1921 (.Y (nx1920), .A0 (nx4766), .A1 (nx4771), .B0 (
                          nx1568), .C0 (nx4785)) ;
    AND4_X0P5M_A12TS ix4767 (.Y (nx4766), .A (nx968), .B (nx1312), .C (nx4617), 
                     .D (nx1068)) ;
    NAND2_X0P5A_A12TS ix969 (.Y (nx968), .A (nx4436), .B (nx4546)) ;
    NAND2_X0P5A_A12TS ix1313 (.Y (nx1312), .A (nx4317), .B (nx4377)) ;
    NAND2_X0P5A_A12TS ix1069 (.Y (nx1068), .A (nx4395), .B (nx4402)) ;
    AOI211_X0P5M_A12TS ix4772 (.Y (nx4771), .A0 (nx4773), .A1 (nx250), .B0 (
                       nx1898), .C0 (nx1872)) ;
    OAI21_X0P5M_A12TS ix1899 (.Y (nx1898), .A0 (nx532), .A1 (nx462), .B0 (nx4777
                      )) ;
    AOI22_X0P5M_A12TS ix4778 (.Y (nx4777), .A0 (nx4779), .A1 (nx250), .B0 (
                      nx4436), .B1 (nx4773)) ;
    NOR2_X0P5A_A12TS ix4780 (.Y (nx4779), .A (nx304), .B (nx266)) ;
    AOI22_X0P5M_A12TS ix1873 (.Y (nx1872), .A0 (nx1084), .A1 (nx488), .B0 (nx946
                      ), .B1 (nx1006)) ;
    NAND2_X0P5A_A12TS ix1085 (.Y (nx1084), .A (nx4285), .B (nx170)) ;
    NAND3_X0P5A_A12TS ix947 (.Y (nx946), .A (op1_cur_1), .B (nx4267), .C (nx4429
                      )) ;
    OAI31_X0P5M_A12TS ix4786 (.Y (nx4785), .A0 (nx406), .A1 (nx4773), .A2 (nx472
                      ), .B0 (nx1850)) ;
    NOR2_X0P5A_A12TS ix1851 (.Y (nx1850), .A (nx1568), .B (nx4446)) ;
    DFFRPQ_X0P5M_A12TS reg_src_sel2_1 (.Q (src_sel2_1), .CK (wb_clk_i), .D (
                       nx4127), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4128 (.Y (nx4127), .A0 (nx4791), .A1 (nx4630), .B0 (
                          wait_data), .C0 (nx4807)) ;
    OA21A1OI2_X0P5M_A12TS ix4792 (.Y (nx4791), .A0 (nx2010), .A1 (nx2002), .B0 (
                          nx4628), .C0 (nx1972)) ;
    NAND3_X0P5A_A12TS ix2011 (.Y (nx2010), .A (nx4794), .B (nx1312), .C (nx1292)
                      ) ;
    OAI21_X0P5M_A12TS ix4795 (.Y (nx4794), .A0 (nx4592), .A1 (nx4456), .B0 (
                      nx4436)) ;
    NAND3_X0P5A_A12TS ix2003 (.Y (nx2002), .A (nx4569), .B (nx4798), .C (nx4800)
                      ) ;
    NAND3_X0P5A_A12TS ix4799 (.Y (nx4798), .A (nx4571), .B (op1_cur_1), .C (
                      nx4429)) ;
    AOI32_X0P5M_A12TS ix4801 (.Y (nx4800), .A0 (nx4802), .A1 (nx4310), .A2 (
                      nx4325), .B0 (nx4436), .B1 (nx4420)) ;
    OA21A1OI2_X0P5M_A12TS ix1973 (.Y (nx1972), .A0 (nx196), .A1 (nx170), .B0 (
                          nx242), .C0 (nx4805)) ;
    NAND2_X0P5A_A12TS ix4808 (.Y (nx4807), .A (src_sel2_1), .B (wait_data)) ;
    SDFFRPQ_X0P5M_A12TS reg_src_sel1_0 (.Q (src_sel1_0), .CK (wb_clk_i), .D (
                        nx1766), .R (wb_rst_i), .SE (wait_data), .SI (src_sel1_0
                        )) ;
    NAND4B_X0P5M_A12TS ix1767 (.Y (nx1766), .AN (nx1730), .B (nx4812), .C (
                       nx4827), .D (nx4834)) ;
    OAI222_X0P5M_A12TS ix1731 (.Y (nx1730), .A0 (nx396), .A1 (nx4694), .B0 (
                       nx4271), .B1 (nx4664), .C0 (nx4460), .C1 (nx4704)) ;
    AOI211_X0P5M_A12TS ix4813 (.Y (nx4812), .A0 (nx804), .A1 (nx1214), .B0 (
                       nx1762), .C0 (nx1742)) ;
    AOI32_X0P5M_A12TS ix4820 (.Y (nx4819), .A0 (nx1748), .A1 (nx4429), .A2 (
                      nx806), .B0 (nx442), .B1 (nx82)) ;
    NOR2_X0P5A_A12TS ix1749 (.Y (nx1748), .A (nx4310), .B (op1_cur_1)) ;
    MXIT2_X0P5M_A12TS ix1743 (.Y (nx1742), .A (nx4823), .B (nx4825), .S0 (nx4299
                      )) ;
    NAND2_X0P5A_A12TS ix4824 (.Y (nx4823), .A (nx4308), .B (nx834)) ;
    NAND2_X0P5A_A12TS ix4826 (.Y (nx4825), .A (nx820), .B (nx4281)) ;
    AOI32_X0P5M_A12TS ix4828 (.Y (nx4827), .A0 (nx820), .A1 (nx124), .A2 (nx4285
                      ), .B0 (nx806), .B1 (nx1712)) ;
    OAI22_X0P5M_A12TS ix1713 (.Y (nx1712), .A0 (op1_cur_2), .A1 (nx4830), .B0 (
                      nx4188), .B1 (nx4832)) ;
    NAND2_X0P5A_A12TS ix4831 (.Y (nx4830), .A (nx4310), .B (op1_cur_0)) ;
    AOI21_X0P5M_A12TS ix4833 (.Y (nx4832), .A0 (op1_cur_1), .A1 (op1_cur_2), .B0 (
                      nx124)) ;
    NAND3_X0P5A_A12TS ix4835 (.Y (nx4834), .A (op1_cur_2), .B (nx4285), .C (
                      nx834)) ;
    DFFRPQ_X0P5M_A12TS reg_src_sel1_1 (.Q (src_sel1_1), .CK (wb_clk_i), .D (
                       nx4097), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix4098 (.Y (nx4097), .A0N (nx4838), .B0 (src_sel1_1), .B1 (
                      wait_data)) ;
    OAI31_X0P5M_A12TS ix4839 (.Y (nx4838), .A0 (nx1820), .A1 (nx1816), .A2 (
                      nx1802), .B0 (nx4226)) ;
    OAI222_X0P5M_A12TS ix1817 (.Y (nx1816), .A0 (nx4662), .A1 (nx4340), .B0 (
                       nx4823), .B1 (nx396), .C0 (nx194), .C1 (nx4844)) ;
    OAI211_X0P5M_A12TS ix1803 (.Y (nx1802), .A0 (nx4278), .A1 (nx4847), .B0 (
                       nx4849), .C0 (nx4853)) ;
    NAND2_X0P5A_A12TS ix4848 (.Y (nx4847), .A (nx4285), .B (nx834)) ;
    AOI222_X0P5M_A12TS ix4850 (.Y (nx4849), .A0 (nx1466), .A1 (nx796), .B0 (
                       nx430), .B1 (nx1002), .C0 (nx756), .C1 (nx1356)) ;
    NOR2_X0P5A_A12TS ix1003 (.Y (nx1002), .A (nx4310), .B (nx84)) ;
    AOI31_X0P5M_A12TS ix4854 (.Y (nx4853), .A0 (nx806), .A1 (nx126), .A2 (nx4348
                      ), .B0 (nx1780)) ;
    NOR3_X0P5A_A12TS ix1781 (.Y (nx1780), .A (nx4825), .B (nx304), .C (nx424)) ;
    SDFFRPQ_X0P5M_A12TS reg_src_sel1_2 (.Q (src_sel1_2), .CK (wb_clk_i), .D (
                        nx1842), .R (wb_rst_i), .SE (wait_data), .SI (src_sel1_2
                        )) ;
    OAI221_X0P5M_A12TS ix1843 (.Y (nx1842), .A0 (nx1254), .A1 (nx84), .B0 (nx442
                       ), .B1 (nx4817), .C0 (nx4858)) ;
    AO21A1AI2_X0P5M_A12TS ix4859 (.Y (nx4858), .A0 (nx4456), .A1 (nx250), .B0 (
                          nx4516), .C0 (nx4257)) ;
    SDFFRPQ_X0P5M_A12TS reg_wr_sfr_0 (.Q (wr_sfr_0__dup_836), .CK (wb_clk_i), .D (
                        nx1282), .R (wb_rst_i), .SE (wait_data), .SI (
                        wr_sfr_0__dup_836)) ;
    NAND4_X0P5A_A12TS ix1283 (.Y (nx1282), .A (nx4865), .B (nx4653), .C (nx4869)
                      , .D (nx4872)) ;
    AOI21_X0P5M_A12TS ix4866 (.Y (nx4865), .A0 (nx4390), .A1 (nx1272), .B0 (
                      nx1228)) ;
    AOI211_X0P5M_A12TS ix1273 (.Y (nx1272), .A0 (nx4354), .A1 (nx4390), .B0 (
                       nx4257), .C0 (nx82)) ;
    AOI21_X0P5M_A12TS ix1229 (.Y (nx1228), .A0 (nx148), .A1 (nx4299), .B0 (
                      nx4823)) ;
    AO21A1AI2_X0P5M_A12TS ix4870 (.Y (nx4869), .A0 (nx4188), .A1 (nx1196), .B0 (
                          nx1188), .C0 (nx4310)) ;
    NOR2_X0P5A_A12TS ix1189 (.Y (nx1188), .A (nx84), .B (nx4446)) ;
    AOI31_X0P5M_A12TS ix4873 (.Y (nx4872), .A0 (nx430), .A1 (nx184), .A2 (nx820)
                      , .B0 (nx1178)) ;
    NOR3_X0P5A_A12TS ix1179 (.Y (nx1178), .A (nx4875), .B (nx160), .C (nx4710)
                     ) ;
    AOI21_X0P5M_A12TS ix4876 (.Y (nx4875), .A0 (nx184), .A1 (nx126), .B0 (nx1168
                      )) ;
    NOR2_X0P5A_A12TS ix1169 (.Y (nx1168), .A (nx184), .B (nx4560)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_sfr_1 (.Q (wr_sfr_1__dup_837), .CK (wb_clk_i), .D (
                       nx4037), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix4038 (.Y (nx4037), .A0 (nx4883), .A1 (wait_data), .B0 (
                      nx4889)) ;
    AOI211_X0P5M_A12TS ix4884 (.Y (nx4883), .A0 (nx4546), .A1 (nx1188), .B0 (
                       nx1324), .C0 (nx1076)) ;
    AOI31_X0P5M_A12TS ix1325 (.Y (nx1324), .A0 (nx968), .A1 (nx1312), .A2 (
                      nx4574), .B0 (nx84)) ;
    OAI21_X0P5M_A12TS ix1077 (.Y (nx1076), .A0 (nx1068), .A1 (nx84), .B0 (nx4887
                      )) ;
    NAND3_X0P5A_A12TS ix4888 (.Y (nx4887), .A (nx4255), .B (nx442), .C (nx78)) ;
    NAND2_X0P5A_A12TS ix4890 (.Y (nx4889), .A (wr_sfr_1__dup_837), .B (wait_data
                      )) ;
    DFFRPQ_X0P5M_A12TS reg_wr (.Q (wr_dup_832), .CK (wb_clk_i), .D (nx3987), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix3988 (.Y (nx3987), .A0 (nx4896), .A1 (nx4907), .B0 (
                          wait_data), .C0 (nx4918)) ;
    NOR3_X0P5A_A12TS ix4897 (.Y (nx4896), .A (nx878), .B (nx860), .C (nx844)) ;
    OA21A1OI2_X0P5M_A12TS ix879 (.Y (nx878), .A0 (nx84), .A1 (nx4899), .B0 (
                          nx4901), .C0 (nx4832)) ;
    NAND2_X0P5A_A12TS ix4902 (.Y (nx4901), .A (nx4348), .B (nx756)) ;
    AO21A1AI2_X0P5M_A12TS ix861 (.Y (nx860), .A0 (nx4514), .A1 (nx200), .B0 (
                          nx224), .C0 (nx4887)) ;
    AO21A1AI2_X0P5M_A12TS ix845 (.Y (nx844), .A0 (nx272), .A1 (nx126), .B0 (
                          nx4825), .C0 (nx4905)) ;
    AO21A1AI2_X0P5M_A12TS ix4906 (.Y (nx4905), .A0 (nx4308), .A1 (nx820), .B0 (
                          nx834), .C0 (nx250)) ;
    AOI211_X0P5M_A12TS ix4908 (.Y (nx4907), .A0 (nx796), .A1 (nx810), .B0 (nx792
                       ), .C0 (nx780)) ;
    OAI22_X0P5M_A12TS ix811 (.Y (nx810), .A0 (nx196), .A1 (nx4271), .B0 (nx4188)
                      , .B1 (nx4910)) ;
    NAND2_X0P5A_A12TS ix4911 (.Y (nx4910), .A (nx160), .B (nx804)) ;
    NOR3_X0P5A_A12TS ix793 (.Y (nx792), .A (nx4901), .B (op1_cur_0), .C (
                     op1_cur_2)) ;
    OAI31_X0P5M_A12TS ix781 (.Y (nx780), .A0 (nx4914), .A1 (nx304), .A2 (nx4297)
                      , .B0 (nx4916)) ;
    AOI21_X0P5M_A12TS ix4915 (.Y (nx4914), .A0 (nx4267), .A1 (nx4275), .B0 (
                      nx756)) ;
    NAND4_X0P5A_A12TS ix4917 (.Y (nx4916), .A (nx194), .B (op1_cur_0), .C (
                      op1_cur_2), .D (nx760)) ;
    NAND2_X0P5A_A12TS ix4919 (.Y (nx4918), .A (wr_dup_832), .B (wait_data)) ;
    INV_X0P5B_A12TS ix343 (.Y (bit_addr), .A (nx4921)) ;
    AOI211_X0P5M_A12TS ix4922 (.Y (nx4921), .A0 (nx4257), .A1 (nx4538), .B0 (
                       nx328), .C0 (nx262)) ;
    OAI21_X0P5M_A12TS ix329 (.Y (nx328), .A0 (nx84), .A1 (nx4621), .B0 (nx4924)
                      ) ;
    OAI222_X0P5M_A12TS ix263 (.Y (nx262), .A0 (nx242), .A1 (nx4466), .B0 (nx200)
                       , .B1 (nx224), .C0 (nx84), .C1 (nx4451)) ;
    SDFFRPQ_X0P5M_A12TS reg_ram_wr_sel_0 (.Q (ram_wr_sel_0__dup_833), .CK (
                        wb_clk_i), .D (nx1046), .R (wb_rst_i), .SE (wait_data), 
                        .SI (ram_wr_sel_0__dup_833)) ;
    OAI211_X0P5M_A12TS ix1047 (.Y (nx1046), .A0 (nx84), .A1 (nx4933), .B0 (
                       nx4944), .C0 (nx4947)) ;
    AND4_X0P5M_A12TS ix4934 (.Y (nx4933), .A (nx4582), .B (nx4514), .C (nx4935)
                     , .D (nx4937)) ;
    AOI22_X0P5M_A12TS ix4936 (.Y (nx4935), .A0 (nx4317), .A1 (nx4592), .B0 (
                      nx4576), .B1 (nx4606)) ;
    AOI211_X0P5M_A12TS ix4938 (.Y (nx4937), .A0 (nx4317), .A1 (nx4546), .B0 (
                       nx930), .C0 (nx904)) ;
    OAI222_X0P5M_A12TS ix931 (.Y (nx930), .A0 (nx450), .A1 (nx4941), .B0 (nx174)
                       , .B1 (nx4294), .C0 (nx532), .C1 (nx364)) ;
    NAND2_X0P5A_A12TS ix451 (.Y (nx450), .A (nx4285), .B (nx4364)) ;
    NAND2_X0P5A_A12TS ix4942 (.Y (nx4941), .A (op1_cur_1), .B (nx4299)) ;
    OAI22_X0P5M_A12TS ix905 (.Y (nx904), .A0 (nx398), .A1 (nx4536), .B0 (nx532)
                      , .B1 (nx308)) ;
    AOI211_X0P5M_A12TS ix4945 (.Y (nx4944), .A0 (nx4779), .A1 (nx254), .B0 (
                       nx288), .C0 (nx860)) ;
    AOI21_X0P5M_A12TS ix289 (.Y (nx288), .A0 (nx4626), .A1 (nx264), .B0 (nx4466)
                      ) ;
    AOI32_X0P5M_A12TS ix4948 (.Y (nx4947), .A0 (nx1020), .A1 (nx184), .A2 (
                      nx4332), .B0 (nx1002), .B1 (nx1012)) ;
    NOR2_X0P5A_A12TS ix1021 (.Y (nx1020), .A (nx532), .B (nx84)) ;
    NOR2_X0P5A_A12TS ix1013 (.Y (nx1012), .A (nx1006), .B (nx948)) ;
    DFFRPQ_X0P5M_A12TS reg_ram_wr_sel_1 (.Q (ram_wr_sel_1__dup_834), .CK (
                       wb_clk_i), .D (nx4007), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4957 (.Y (nx4956), .A0 (nx1136), .A1 (nx1076), .A2 (
                      nx1066), .B0 (nx4226)) ;
    AOI31_X0P5M_A12TS ix1137 (.Y (nx1136), .A0 (nx4959), .A1 (nx4798), .A2 (
                      nx4961), .B0 (nx84)) ;
    AOI32_X0P5M_A12TS ix4962 (.Y (nx4961), .A0 (nx4402), .A1 (nx184), .A2 (nx170
                      ), .B0 (nx4576), .B1 (nx4395)) ;
    DFFRPQ_X0P5M_A12TS reg_ram_wr_sel_2 (.Q (ram_wr_sel_2__dup_835), .CK (
                       wb_clk_i), .D (nx4017), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4970 (.Y (nx4969), .A0 (nx4382), .A1 (nx1020), .B0 (
                          nx850), .C0 (nx4226)) ;
    OAI21_X0P5M_A12TS ix2439 (.Y (ram_rd_sel_0), .A0 (wait_data), .A1 (nx4973), 
                      .B0 (nx4994)) ;
    NOR3_X0P5A_A12TS ix461 (.Y (nx460), .A (nx150), .B (nx4273), .C (nx304)) ;
    NAND4_X0P5A_A12TS ix2415 (.Y (nx2414), .A (nx1256), .B (nx1068), .C (nx4977)
                      , .D (nx4983)) ;
    NOR3_X0P5A_A12TS ix4978 (.Y (nx4977), .A (nx1302), .B (nx4981), .C (nx4448)
                     ) ;
    OAI21_X0P5M_A12TS ix1303 (.Y (nx1302), .A0 (nx946), .A1 (nx492), .B0 (nx1292
                      )) ;
    NOR2_X0P5A_A12TS ix4982 (.Y (nx4981), .A (nx306), .B (nx398)) ;
    NOR3_X0P5A_A12TS ix4984 (.Y (nx4983), .A (nx2394), .B (nx2388), .C (nx2084)
                     ) ;
    NAND3_X0P5A_A12TS ix2395 (.Y (nx2394), .A (nx4935), .B (nx4415), .C (nx4798)
                      ) ;
    OAI31_X0P5M_A12TS ix2389 (.Y (nx2388), .A0 (nx4987), .A1 (nx194), .A2 (nx488
                      ), .B0 (nx4989)) ;
    OAI22_X0P5M_A12TS ix2085 (.Y (nx2084), .A0 (nx508), .A1 (nx952), .B0 (nx2046
                      ), .B1 (nx4987)) ;
    NAND2_X0P5A_A12TS ix4995 (.Y (nx4994), .A (wait_data), .B (ram_rd_sel_r_0)
                      ) ;
    DFFRPQ_X0P5M_A12TS reg_ram_rd_sel_r_0 (.Q (ram_rd_sel_r_0), .CK (wb_clk_i), 
                       .D (nx2426), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2427 (.Y (nx2426), .A0 (nx4482), .A1 (nx4478), .B0 (
                      nx4998)) ;
    AOI22_X0P5M_A12TS ix4999 (.Y (nx4998), .A0 (nx460), .A1 (nx4478), .B0 (
                      nx4275), .B1 (nx2414)) ;
    OAI21_X0P5M_A12TS ix2513 (.Y (ram_rd_sel_1), .A0 (wait_data), .A1 (nx5001), 
                      .B0 (nx5018)) ;
    AOI21_X0P5M_A12TS ix5004 (.Y (nx5003), .A0 (nx78), .A1 (nx658), .B0 (nx328)
                      ) ;
    AOI32_X0P5M_A12TS ix5007 (.Y (nx5006), .A0 (nx1002), .A1 (nx4325), .A2 (
                      nx4444), .B0 (nx1020), .B1 (nx2484)) ;
    NAND3_X0P5A_A12TS ix2485 (.Y (nx2484), .A (nx242), .B (nx1242), .C (nx4536)
                      ) ;
    OAI21_X0P5M_A12TS ix5010 (.Y (nx5009), .A0 (nx2462), .A1 (nx2452), .B0 (
                      nx4275)) ;
    NAND4_X0P5A_A12TS ix2463 (.Y (nx2462), .A (nx4415), .B (nx332), .C (nx5012)
                      , .D (nx4777)) ;
    NOR2_X0P5A_A12TS ix5013 (.Y (nx5012), .A (nx216), .B (nx1128)) ;
    OAI22_X0P5M_A12TS ix1129 (.Y (nx1128), .A0 (nx150), .A1 (nx274), .B0 (nx946)
                      , .B1 (nx516)) ;
    NAND3_X0P5A_A12TS ix2453 (.Y (nx2452), .A (nx4600), .B (nx4582), .C (nx5016)
                      ) ;
    AOI211_X0P5M_A12TS ix5017 (.Y (nx5016), .A0 (nx4317), .A1 (nx4592), .B0 (
                       nx930), .C0 (nx904)) ;
    NAND2_X0P5A_A12TS ix5019 (.Y (nx5018), .A (wait_data), .B (ram_rd_sel_r_1)
                      ) ;
    DFFRPQ_X0P5M_A12TS reg_ram_rd_sel_r_1 (.Q (ram_rd_sel_r_1), .CK (wb_clk_i), 
                       .D (nx2500), .R (wb_rst_i)) ;
    NAND4_X0P5A_A12TS ix2501 (.Y (nx2500), .A (nx5003), .B (comp_sel_0), .C (
                      nx5006), .D (nx5009)) ;
    OAI21_X0P5M_A12TS ix2545 (.Y (ram_rd_sel_2), .A0 (wait_data), .A1 (nx5023), 
                      .B0 (nx5029)) ;
    NAND2_X0P5A_A12TS ix5030 (.Y (nx5029), .A (wait_data), .B (ram_rd_sel_r_2)
                      ) ;
    DFFRPQ_X0P5M_A12TS reg_ram_rd_sel_r_2 (.Q (ram_rd_sel_r_2), .CK (wb_clk_i), 
                       .D (nx2532), .R (wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix2533 (.Y (nx2532), .A0 (nx84), .A1 (nx5033), .B0 (
                       comp_sel_0), .C0 (nx4390)) ;
    NOR3_X0P5A_A12TS ix5034 (.Y (nx5033), .A (nx5027), .B (nx4578), .C (nx4981)
                     ) ;
    INV_X0P5B_A12TS ix5024 (.Y (nx5023), .A (nx2532)) ;
    INV_X0P5B_A12TS ix5002 (.Y (nx5001), .A (nx2500)) ;
    INV_X0P5B_A12TS ix4974 (.Y (nx4973), .A (nx2426)) ;
    INV_X0P5B_A12TS ix4603 (.Y (nx4602), .A (nx2084)) ;
    INV_X0P5B_A12TS ix4605 (.Y (nx4604), .A (nx2046)) ;
    INV_X0P5B_A12TS ix4631 (.Y (nx4630), .A (nx1952)) ;
    INV_X0P5B_A12TS ix4806 (.Y (nx4805), .A (nx1850)) ;
    INV_X0P5B_A12TS ix4629 (.Y (nx4628), .A (nx1568)) ;
    INV_X0P5B_A12TS ix4551 (.Y (nx4550), .A (nx1540)) ;
    INV_X0P5B_A12TS ix1467 (.Y (nx1466), .A (nx4694)) ;
    INV_X0P5B_A12TS ix1397 (.Y (nx1396), .A (nx4340)) ;
    INV_X0P5B_A12TS ix1293 (.Y (nx1292), .A (nx4578)) ;
    INV_X0P5B_A12TS ix4818 (.Y (nx4817), .A (nx1272)) ;
    INV_X0P5B_A12TS ix5028 (.Y (nx5027), .A (nx1256)) ;
    INV_X0P5B_A12TS ix4693 (.Y (nx4692), .A (nx1214)) ;
    INV_X0P5B_A12TS ix4845 (.Y (nx4844), .A (nx1196)) ;
    INV_X0P5B_A12TS ix4665 (.Y (nx4664), .A (nx1168)) ;
    INV_X0P5B_A12TS ix4960 (.Y (nx4959), .A (nx1128)) ;
    INV_X0P5B_A12TS ix1067 (.Y (nx1066), .A (nx4858)) ;
    INV_X0P5B_A12TS ix1007 (.Y (nx1006), .A (nx4325)) ;
    INV_X0P5B_A12TS ix953 (.Y (nx952), .A (nx4606)) ;
    INV_X0P5B_A12TS ix4803 (.Y (nx4802), .A (nx948)) ;
    INV_X0P5B_A12TS ix4577 (.Y (nx4576), .A (nx946)) ;
    INV_X0P5B_A12TS ix915 (.Y (nx914), .A (nx4941)) ;
    INV_X0P5B_A12TS ix4900 (.Y (nx4899), .A (nx870)) ;
    INV_X0P5B_A12TS ix851 (.Y (nx850), .A (nx4887)) ;
    INV_X0P5B_A12TS ix4663 (.Y (nx4662), .A (nx834)) ;
    INV_X0P5B_A12TS ix808 (.Y (nx806), .A (nx4910)) ;
    INV_X0P5B_A12TS ix4711 (.Y (nx4710), .A (nx804)) ;
    INV_X0P5B_A12TS ix4339 (.Y (nx4338), .A (nx796)) ;
    INV_X0P5B_A12TS ix795 (.Y (nx794), .A (nx4699)) ;
    INV_X0P5B_A12TS ix785 (.Y (nx784), .A (nx4901)) ;
    INV_X0P5B_A12TS ix757 (.Y (nx756), .A (nx4271)) ;
    INV_X0P5B_A12TS ix659 (.Y (nx658), .A (nx4482)) ;
    INV_X0P5B_A12TS ix583 (.Y (nx582), .A (nx4526)) ;
    INV_X0P5B_A12TS ix4423 (.Y (nx4422), .A (nx564)) ;
    INV_X0P5B_A12TS ix545 (.Y (nx544), .A (nx4434)) ;
    INV_X0P5B_A12TS ix4437 (.Y (nx4436), .A (nx532)) ;
    INV_X0P5B_A12TS ix4618 (.Y (nx4617), .A (nx530)) ;
    INV_X0P5B_A12TS ix4405 (.Y (nx4404), .A (nx516)) ;
    INV_X0P5B_A12TS ix509 (.Y (nx508), .A (nx4402)) ;
    INV_X0P5B_A12TS ix4260 (.Y (nx4259), .A (nx506)) ;
    INV_X0P5B_A12TS ix493 (.Y (nx492), .A (nx4395)) ;
    INV_X0P5B_A12TS ix485 (.Y (nx484), .A (nx4398)) ;
    INV_X0P5B_A12TS ix473 (.Y (nx472), .A (nx4536)) ;
    INV_X0P5B_A12TS ix463 (.Y (nx462), .A (nx4779)) ;
    INV_X0P5B_A12TS ix4774 (.Y (nx4773), .A (nx450)) ;
    INV_X0P5B_A12TS ix4391 (.Y (nx4390), .A (nx442)) ;
    INV_X0P5B_A12TS ix435 (.Y (nx434), .A (nx4685)) ;
    INV_X0P5B_A12TS ix431 (.Y (nx430), .A (nx4446)) ;
    INV_X0P5B_A12TS ix4430 (.Y (nx4429), .A (nx424)) ;
    INV_X0P5B_A12TS ix4615 (.Y (nx4614), .A (nx406)) ;
    INV_X0P5B_A12TS ix401 (.Y (nx400), .A (nx4981)) ;
    INV_X0P5B_A12TS ix399 (.Y (nx398), .A (nx4356)) ;
    INV_X0P5B_A12TS ix4515 (.Y (nx4514), .A (nx376)) ;
    INV_X0P5B_A12TS ix4472 (.Y (nx4471), .A (nx368)) ;
    INV_X0P5B_A12TS ix365 (.Y (nx364), .A (nx4420)) ;
    INV_X0P5B_A12TS ix4517 (.Y (nx4516), .A (nx352)) ;
    INV_X0P5B_A12TS ix347 (.Y (nx346), .A (nx4281)) ;
    INV_X0P5B_A12TS ix333 (.Y (nx332), .A (nx4538)) ;
    INV_X0P5B_A12TS ix309 (.Y (nx308), .A (nx4382)) ;
    INV_X0P5B_A12TS ix305 (.Y (nx304), .A (nx4285)) ;
    INV_X0P5B_A12TS ix4591 (.Y (nx4590), .A (nx290)) ;
    INV_X0P5B_A12TS ix4925 (.Y (nx4924), .A (nx288)) ;
    INV_X0P5B_A12TS ix283 (.Y (nx282), .A (nx4626)) ;
    INV_X0P5B_A12TS ix277 (.Y (nx276), .A (nx4592)) ;
    INV_X0P5B_A12TS ix275 (.Y (nx274), .A (nx4546)) ;
    INV_X0P5B_A12TS ix273 (.Y (nx272), .A (nx4348)) ;
    INV_X0P5B_A12TS ix265 (.Y (nx264), .A (nx4377)) ;
    INV_X0P5B_A12TS ix255 (.Y (nx254), .A (nx4466)) ;
    INV_X0P5B_A12TS ix4461 (.Y (nx4460), .A (nx250)) ;
    INV_X0P5B_A12TS ix4440 (.Y (nx4439), .A (nx242)) ;
    INV_X0P5B_A12TS ix4309 (.Y (nx4308), .A (nx234)) ;
    INV_X0P5B_A12TS ix225 (.Y (nx224), .A (nx4478)) ;
    INV_X0P5B_A12TS ix4452 (.Y (nx4451), .A (nx216)) ;
    INV_X0P5B_A12TS ix199 (.Y (nx198), .A (nx4456)) ;
    INV_X0P5B_A12TS ix4425 (.Y (nx4424), .A (nx196)) ;
    INV_X0P5B_A12TS ix195 (.Y (nx194), .A (nx4310)) ;
    INV_X0P5B_A12TS ix185 (.Y (nx184), .A (nx4188)) ;
    INV_X0P5B_A12TS ix4433 (.Y (nx4432), .A (nx174)) ;
    INV_X0P5B_A12TS ix171 (.Y (nx170), .A (nx4273)) ;
    INV_X0P5B_A12TS ix161 (.Y (nx160), .A (nx4267)) ;
    INV_X0P5B_A12TS ix4318 (.Y (nx4317), .A (nx150)) ;
    INV_X0P5B_A12TS ix149 (.Y (nx148), .A (nx4361)) ;
    INV_X0P5B_A12TS ix127 (.Y (nx126), .A (nx4299)) ;
    INV_X0P5B_A12TS ix125 (.Y (nx124), .A (nx4278)) ;
    INV_X0P5B_A12TS ix4491 (.Y (nx4490), .A (nx98)) ;
    INV_X0P5B_A12TS ix4276 (.Y (nx4275), .A (nx84)) ;
    INV_X0P5B_A12TS ix83 (.Y (nx82), .A (nx4255)) ;
    INV_X0P5B_A12TS ix79 (.Y (nx78), .A (nx4257)) ;
    INV_X0P5B_A12TS ix4192 (.Y (NOT_nx10), .A (nx10)) ;
    INV_X0P5B_A12TS ix137 (.Y (op1_cur_1), .A (nx4372)) ;
    NAND4B_X0P5M_A12TS ix4217 (.Y (nx4216), .AN (op1_n_4), .B (op1_n_2), .C (
                       nx24), .D (op1_n_7)) ;
    AO22_X0P5M_A12TS ix147 (.Y (op1_cur_0), .A0 (op1_n_0), .A1 (nx110), .B0 (
                     op_0), .B1 (nx102)) ;
    AO22_X0P5M_A12TS ix115 (.Y (op1_cur_2), .A0 (op1_n_2), .A1 (nx110), .B0 (
                     op_2), .B1 (nx102)) ;
    AND2_X0P5M_A12TS ix4282 (.Y (nx4281), .A (op1_cur_0), .B (nx4372)) ;
    OR2_X0P5M_A12TS ix507 (.Y (nx506), .A (nx4372), .B (nx4267)) ;
    NAND4B_X0P5M_A12TS ix1241 (.Y (nx1240), .AN (nx1080), .B (nx4299), .C (
                       op1_cur_1), .D (nx4267)) ;
    AO1B2_X0P5M_A12TS ix377 (.Y (nx376), .A0N (nx352), .B0 (nx4456), .B1 (nx250)
                      ) ;
    NAND4B_X0P5M_A12TS ix4487 (.Y (nx4486), .AN (op1_n_0), .B (op1_n_1), .C (
                       nx4214), .D (nx4302)) ;
    NAND4B_X0P5M_A12TS ix4489 (.Y (nx4488), .AN (op1_n_6), .B (op1_n_5), .C (
                       nx4288), .D (nx4490)) ;
    NAND3B_X0P5M_A12TS ix4493 (.Y (nx4492), .AN (op_3), .B (nx608), .C (op_5)) ;
    NAND4B_X0P5M_A12TS ix4499 (.Y (nx4498), .AN (nx656), .B (nx4390), .C (nx570)
                       , .D (nx4478)) ;
    NAND2B_X0P7M_A12TS ix4561 (.Y (nx4560), .AN (nx4297), .B (op1_cur_0)) ;
    OA211_X0P5M_A12TS ix4583 (.Y (nx4582), .A0 (nx242), .A1 (nx4460), .B0 (
                      nx4794), .C0 (nx968)) ;
    NAND4B_X0P5M_A12TS ix2121 (.Y (nx2120), .AN (nx2054), .B (nx4600), .C (
                       nx4602), .D (nx4608)) ;
    AO1B2_X0P5M_A12TS ix4048 (.Y (nx4047), .A0N (nx4649), .B0 (alu_op_0__dup_838
                      ), .B1 (wait_data)) ;
    NAND3B_X0P5M_A12TS ix4674 (.Y (nx4673), .AN (nx4560), .B (nx4310), .C (nx820
                       )) ;
    NOR2B_X0P7M_A12TS ix1503 (.Y (alu_op_1), .AN (alu_op_1__dup_839), .B (
                      wait_data)) ;
    AO1B2_X0P5M_A12TS ix1455 (.Y (nx1454), .A0N (nx4704), .B0 (nx4348), .B1 (
                      nx760)) ;
    NOR2B_X0P7M_A12TS ix1565 (.Y (alu_op_2), .AN (alu_op_2__dup_840), .B (
                      wait_data)) ;
    AO22_X0P5M_A12TS ix1527 (.Y (nx1526), .A0 (nx4348), .A1 (nx820), .B0 (nx4382
                     ), .B1 (nx84)) ;
    AO1B2_X0P5M_A12TS ix4078 (.Y (nx4077), .A0N (nx4737), .B0 (alu_op_3__dup_841
                      ), .B1 (wait_data)) ;
    NAND3B_X0P5M_A12TS ix1763 (.Y (nx1762), .AN (nx1188), .B (nx4817), .C (
                       nx4819)) ;
    NAND3B_X0P5M_A12TS ix1821 (.Y (nx1820), .AN (nx1228), .B (nx4817), .C (
                       nx4819)) ;
    NOR2B_X0P7M_A12TS ix1291 (.Y (wr_sfr_0), .AN (wr_sfr_0__dup_836), .B (
                      wait_data)) ;
    NOR2B_X0P7M_A12TS ix1341 (.Y (wr_sfr_1), .AN (wr_sfr_1__dup_837), .B (
                      wait_data)) ;
    NOR2B_X0P7M_A12TS ix893 (.Y (wr), .AN (wr_dup_832), .B (wait_data)) ;
    NOR2B_X0P7M_A12TS ix1055 (.Y (ram_wr_sel_0), .AN (ram_wr_sel_0__dup_833), .B (
                      wait_data)) ;
    AO1B2_X0P5M_A12TS ix4008 (.Y (nx4007), .A0N (nx4956), .B0 (
                      ram_wr_sel_1__dup_834), .B1 (wait_data)) ;
    AO1B2_X0P5M_A12TS ix4018 (.Y (nx4017), .A0N (nx4969), .B0 (
                      ram_wr_sel_2__dup_835), .B1 (wait_data)) ;
    OR2_X0P5M_A12TS ix4988 (.Y (nx4987), .A (nx4372), .B (nx424)) ;
    OR3_X0P5M_A12TS ix4990 (.Y (nx4989), .A (nx946), .B (nx4188), .C (nx4273)) ;
    NOR2B_X0P7M_A12TS ix1419 (.Y (alu_op_0), .AN (alu_op_0__dup_838), .B (
                      wait_data)) ;
    NOR2B_X0P7M_A12TS ix1635 (.Y (alu_op_3), .AN (alu_op_3__dup_841), .B (
                      wait_data)) ;
    NOR2B_X0P7M_A12TS ix1149 (.Y (ram_wr_sel_1), .AN (ram_wr_sel_1__dup_834), .B (
                      wait_data)) ;
    NOR2B_X0P7M_A12TS ix1163 (.Y (ram_wr_sel_2), .AN (ram_wr_sel_2__dup_835), .B (
                      wait_data)) ;
    INV_X0P5B_A12TS ix1496 (.Y (nx1495), .A (alu_op_1)) ;
    NOR2_X0P5A_A12TS ix173 (.Y (enable_mul), .A (nx1501), .B (nx12)) ;
    NAND2_X0P5A_A12TS ix1502 (.Y (nx1501), .A (alu_op_1), .B (alu_op_0)) ;
    INV_X0P5B_A12TS ix1506 (.Y (nx1505), .A (alu_op_2)) ;
    OAI21_X0P5M_A12TS ix89 (.Y (sub_result_0), .A0 (alu_cy), .A1 (nx1509), .B0 (
                      nx80)) ;
    AOI21_X0P5M_A12TS ix1510 (.Y (nx1509), .A0 (src1_0), .A1 (nx1511), .B0 (
                      nx1513)) ;
    NAND2_X0P5A_A12TS ix1512 (.Y (nx1511), .A (src2_0), .B (src1_0)) ;
    NOR2B_X0P7M_A12TS ix1514 (.Y (nx1513), .AN (src2_0), .B (src1_0)) ;
    NAND2_X0P5A_A12TS ix81 (.Y (nx80), .A (nx1509), .B (alu_cy)) ;
    XOR2_X0P5M_A12TS ix842 (.Y (sub_result_1), .A (nx80), .B (nx1519)) ;
    XOR2_X0P5M_A12TS ix1520 (.Y (nx1519), .A (nx1521), .B (nx1513)) ;
    OAI21_X0P5M_A12TS ix1522 (.Y (nx1521), .A0 (src1_1), .A1 (src2_1), .B0 (
                      nx1523)) ;
    NAND2_X0P5A_A12TS ix1524 (.Y (nx1523), .A (src2_1), .B (src1_1)) ;
    XOR2_X0P5M_A12TS ix465 (.Y (sub_result_2), .A (nx298), .B (nx1539)) ;
    INV_X0P5B_A12TS ix1534 (.Y (nx1533), .A (src1_0)) ;
    INV_X0P5B_A12TS ix1538 (.Y (nx1537), .A (alu_cy)) ;
    XNOR2_X0P5M_A12TS ix1540 (.Y (nx1539), .A (nx1541), .B (nx454)) ;
    OAI21_X0P5M_A12TS ix1542 (.Y (nx1541), .A0 (src1_2), .A1 (src2_2), .B0 (
                      nx1543)) ;
    NAND2_X0P5A_A12TS ix1544 (.Y (nx1543), .A (src2_2), .B (src1_2)) ;
    CGENI_X1M_A12TS ix455 (.CON (nx454), .A (nx1547), .B (nx1513), .CI (src2_1)
                    ) ;
    INV_X0P5B_A12TS ix1548 (.Y (nx1547), .A (src1_1)) ;
    XOR2_X0P5M_A12TS ix587 (.Y (sub_result_3), .A (nx458), .B (nx1557)) ;
    XOR2_X0P5M_A12TS ix1558 (.Y (nx1557), .A (nx1559), .B (nx1563)) ;
    OAI21_X0P5M_A12TS ix1560 (.Y (nx1559), .A0 (src1_3), .A1 (src2_3), .B0 (
                      nx1561)) ;
    NAND2_X0P5A_A12TS ix1562 (.Y (nx1561), .A (src2_3), .B (src1_3)) ;
    CGENI_X1M_A12TS ix1564 (.CON (nx1563), .A (src1_2), .B (nx454), .CI (nx1565)
                    ) ;
    INV_X0P5B_A12TS ix1566 (.Y (nx1565), .A (src2_2)) ;
    XNOR2_X0P5M_A12TS ix721 (.Y (sub_result_4), .A (nx1569), .B (nx1581)) ;
    XOR2_X0P5M_A12TS ix1570 (.Y (nx1569), .A (nx580), .B (nx710)) ;
    CGENI_X1M_A12TS ix843 (.CON (nx710), .A (nx1579), .B (nx1563), .CI (src2_3)
                    ) ;
    INV_X0P5B_A12TS ix1580 (.Y (nx1579), .A (src1_3)) ;
    AOI21_X0P5M_A12TS ix1582 (.Y (nx1581), .A0 (src1_4), .A1 (nx1583), .B0 (
                      nx1585)) ;
    NAND2_X0P5A_A12TS ix1584 (.Y (nx1583), .A (src2_4), .B (src1_4)) ;
    NOR2B_X0P7M_A12TS ix1586 (.Y (nx1585), .AN (src2_4), .B (src1_4)) ;
    XOR2_X0P5M_A12TS ix844 (.Y (sub_result_5), .A (nx714), .B (nx1591)) ;
    NAND2_X0P5A_A12TS ix715 (.Y (nx714), .A (nx1581), .B (nx1569)) ;
    XOR2_X0P5M_A12TS ix1592 (.Y (nx1591), .A (nx1593), .B (nx1585)) ;
    OAI21_X0P5M_A12TS ix1594 (.Y (nx1593), .A0 (src1_5), .A1 (src2_5), .B0 (
                      nx1595)) ;
    NAND2_X0P5A_A12TS ix1596 (.Y (nx1595), .A (src2_5), .B (src1_5)) ;
    XOR2_X0P5M_A12TS ix985 (.Y (sub_result_6), .A (nx836), .B (nx1603)) ;
    XNOR2_X0P5M_A12TS ix1604 (.Y (nx1603), .A (nx1605), .B (nx996)) ;
    OAI21_X0P5M_A12TS ix1606 (.Y (nx1605), .A0 (src1_6), .A1 (src2_6), .B0 (
                      nx1607)) ;
    NAND2_X0P5A_A12TS ix1608 (.Y (nx1607), .A (src2_6), .B (src1_6)) ;
    CGENI_X1M_A12TS ix975 (.CON (nx996), .A (nx1611), .B (nx1585), .CI (src2_5)
                    ) ;
    INV_X0P5B_A12TS ix1612 (.Y (nx1611), .A (src1_5)) ;
    XNOR2_X0P5M_A12TS ix846 (.Y (sub_result_7), .A (nx1615), .B (nx1627)) ;
    XNOR2_X0P5M_A12TS ix1616 (.Y (nx1615), .A (nx997), .B (nx1623)) ;
    CGENI_X1M_A12TS ix1624 (.CON (nx1623), .A (src1_6), .B (nx996), .CI (nx1625)
                    ) ;
    INV_X0P5B_A12TS ix1626 (.Y (nx1625), .A (src2_6)) ;
    OAI21_X0P5M_A12TS ix1628 (.Y (nx1627), .A0 (src1_7), .A1 (src2_7), .B0 (
                      nx1629)) ;
    NAND2_X0P5A_A12TS ix1630 (.Y (nx1629), .A (src2_7), .B (src1_7)) ;
    OAI211_X0P5M_A12TS ix1665 (.Y (desOv), .A0 (nx1633), .A1 (nx1639), .B0 (
                       nx1645), .C0 (nx1693)) ;
    XOR2_X0P5M_A12TS ix1634 (.Y (nx1633), .A (nx1615), .B (nx1614)) ;
    CGENI_X1M_A12TS ix1615 (.CON (nx1614), .A (nx1637), .B (src2_7), .CI (nx1615
                    )) ;
    INV_X0P5B_A12TS ix1638 (.Y (nx1637), .A (src1_7)) ;
    NAND2_X0P5A_A12TS ix1640 (.Y (nx1639), .A (nx1641), .B (nx1643)) ;
    NOR2_X0P5A_A12TS ix1642 (.Y (nx1641), .A (alu_op_0), .B (nx1495)) ;
    NOR2_X0P5A_A12TS ix1644 (.Y (nx1643), .A (alu_op_2), .B (alu_op_3)) ;
    AOI22_X0P5M_A12TS ix1646 (.Y (nx1645), .A0 (mulOv), .A1 (enable_mul), .B0 (
                      nx1658), .B1 (nx50)) ;
    XNOR2_X0P5M_A12TS ix1659 (.Y (nx1658), .A (nx1172), .B (nx1651)) ;
    OAI21_X0P5M_A12TS ix1173 (.Y (nx1172), .A0 (nx1651), .A1 (nx1689), .B0 (
                      nx1629)) ;
    XOR2_X0P5M_A12TS ix1652 (.Y (nx1651), .A (nx1653), .B (nx882)) ;
    CGENI_X1M_A12TS ix1654 (.CON (nx1653), .A (nx868), .B (src1_6), .CI (src2_6)
                    ) ;
    OAI21_X0P5M_A12TS ix869 (.Y (nx868), .A0 (nx1583), .A1 (nx1657), .B0 (nx1595
                      )) ;
    NOR2_X0P5A_A12TS ix1658 (.Y (nx1657), .A (src1_5), .B (src2_5)) ;
    NOR2_X0P5A_A12TS ix883 (.Y (nx882), .A (nx1661), .B (nx1663)) ;
    XOR2_X0P5M_A12TS ix1662 (.Y (nx1661), .A (nx868), .B (nx1605)) ;
    NOR2_X0P5A_A12TS ix643 (.Y (nx642), .A (nx1668), .B (nx1581)) ;
    XNOR2_X0P5M_A12TS ix1669 (.Y (nx1668), .A (nx622), .B (nx514)) ;
    OAI21_X0P5M_A12TS ix623 (.Y (nx622), .A0 (nx1671), .A1 (nx1676), .B0 (nx1561
                      )) ;
    CGENI_X1M_A12TS ix1672 (.CON (nx1671), .A (nx350), .B (src1_2), .CI (src2_2)
                    ) ;
    OAI21_X0P5M_A12TS ix351 (.Y (nx350), .A0 (nx1511), .A1 (nx1674), .B0 (nx1523
                      )) ;
    NOR2_X0P5A_A12TS ix1675 (.Y (nx1674), .A (src1_1), .B (src2_1)) ;
    NOR2_X0P5A_A12TS ix1677 (.Y (nx1676), .A (src1_3), .B (src2_3)) ;
    NOR2_X0P5A_A12TS ix515 (.Y (nx514), .A (nx1679), .B (nx1681)) ;
    XNOR2_X0P5M_A12TS ix1680 (.Y (nx1679), .A (nx1671), .B (nx1559)) ;
    NOR2_X0P5A_A12TS ix847 (.Y (nx973), .A (nx1685), .B (nx1687)) ;
    XNOR2_X0P5M_A12TS ix1686 (.Y (nx1685), .A (nx1511), .B (nx1521)) ;
    NOR2_X0P5A_A12TS ix1690 (.Y (nx1689), .A (src1_7), .B (src2_7)) ;
    NOR2_X0P5A_A12TS ix51 (.Y (nx50), .A (nx2), .B (nx12)) ;
    NAND2_X0P5A_A12TS ix848 (.Y (nx2), .A (alu_op_0), .B (nx1495)) ;
    NAND2_X0P5A_A12TS ix1694 (.Y (nx1693), .A (divOv), .B (enable_div)) ;
    OAI21_X0P5M_A12TS ix1647 (.Y (desAc), .A0 (nx1668), .A1 (nx1696), .B0 (
                      nx1700)) ;
    AOI22_X0P5M_A12TS ix1701 (.Y (nx1700), .A0 (srcAc), .A1 (nx22), .B0 (nx1569)
                      , .B1 (nx94)) ;
    NAND4_X0P5A_A12TS ix849 (.Y (desCy), .A (nx1706), .B (nx1718), .C (nx1001), 
                      .D (nx1733)) ;
    AOI211_X0P5M_A12TS ix1707 (.Y (nx1706), .A0 (src1_7), .A1 (nx971), .B0 (
                       nx1630), .C0 (nx1618)) ;
    NOR2_X0P5A_A12TS ix850 (.Y (nx971), .A (nx1501), .B (nx970)) ;
    NAND2_X0P5A_A12TS ix852 (.Y (nx970), .A (nx1505), .B (alu_op_3)) ;
    OAI22_X0P5M_A12TS ix1631 (.Y (nx1630), .A0 (alu_cy), .A1 (nx1711), .B0 (
                      nx1714), .B1 (nx1696)) ;
    NAND2_X0P5A_A12TS ix1712 (.Y (nx1711), .A (nx1641), .B (nx6)) ;
    NOR2_X0P5A_A12TS ix7 (.Y (nx6), .A (alu_op_3), .B (nx1505)) ;
    NOR2_X0P5A_A12TS ix1619 (.Y (nx1618), .A (nx1614), .B (nx1639)) ;
    OAI31_X0P5M_A12TS ix1719 (.Y (nx1718), .A0 (nx22), .A1 (nx252), .A2 (nx1598)
                      , .B0 (alu_cy)) ;
    NOR2_X0P5A_A12TS ix253 (.Y (nx252), .A (nx970), .B (nx2)) ;
    OAI221_X0P5M_A12TS ix1599 (.Y (nx1598), .A0 (nx970), .A1 (nx60), .B0 (nx1722
                       ), .B1 (nx1724), .C0 (nx1727)) ;
    INV_X0P5B_A12TS ix1723 (.Y (nx1722), .A (bit_out)) ;
    NAND3_X0P5A_A12TS ix1728 (.Y (nx1727), .A (nx1722), .B (alu_op_3), .C (nx18)
                      ) ;
    NOR2_X0P5A_A12TS ix19 (.Y (nx18), .A (alu_op_1), .B (alu_op_0)) ;
    AO21A1AI2_X0P5M_A12TS ix853 (.Y (nx1001), .A0 (nx1537), .A1 (nx222), .B0 (
                          nx252), .C0 (bit_out)) ;
    OA21A1OI2_X0P5M_A12TS ix1734 (.Y (nx1733), .A0 (nx1546), .A1 (nx326), .B0 (
                          nx969), .C0 (nx1000)) ;
    XNOR3_X0P5M_A12TS ix1547 (.Y (nx1546), .A (nx1736), .B (alu_cy), .C (nx1032)
                      ) ;
    OAI21_X0P5M_A12TS ix1737 (.Y (nx1736), .A0 (src1_6), .A1 (src1_5), .B0 (
                      src1_7)) ;
    OAI31_X0P5M_A12TS ix1740 (.Y (nx1739), .A0 (src1_6), .A1 (src1_5), .A2 (
                      src1_7), .B0 (nx1736)) ;
    NAND2_X0P5A_A12TS ix1744 (.Y (nx1743), .A (src1_4), .B (nx326)) ;
    NOR2_X0P5A_A12TS ix1747 (.Y (nx1746), .A (src1_2), .B (src1_1)) ;
    OAI31_X0P5M_A12TS ix854 (.Y (nx1000), .A0 (nx60), .A1 (bit_out), .A2 (nx970)
                      , .B0 (nx1750)) ;
    NAND3_X0P5A_A12TS ix1751 (.Y (nx1750), .A (nx972), .B (src1_0), .C (nx1698)
                      ) ;
    NAND3_X0P5A_A12TS ix181 (.Y (des_acc_0), .A (nx1754), .B (nx1770), .C (
                      nx1773)) ;
    AOI21_X0P5M_A12TS ix1755 (.Y (nx1754), .A0 (mulsrc1_0), .A1 (enable_mul), .B0 (
                      nx168)) ;
    OAI21_X0P5M_A12TS ix169 (.Y (nx168), .A0 (alu_op_0), .A1 (nx1757), .B0 (
                      nx1760)) ;
    AOI32_X0P5M_A12TS ix1758 (.Y (nx1757), .A0 (nx1533), .A1 (alu_op_1), .A2 (
                      alu_op_2), .B0 (nx40), .B1 (nx128)) ;
    NOR2_X0P5A_A12TS ix129 (.Y (nx128), .A (alu_op_1), .B (nx970)) ;
    AO21A1AI2_X0P5M_A12TS ix1761 (.Y (nx1760), .A0 (src1_0), .A1 (nx128), .B0 (
                          nx162), .C0 (alu_op_0)) ;
    OAI21_X0P5M_A12TS ix163 (.Y (nx162), .A0 (nx1511), .A1 (nx1763), .B0 (nx1765
                      )) ;
    NAND2_X0P5A_A12TS ix1764 (.Y (nx1763), .A (alu_op_1), .B (nx6)) ;
    OAI21_X0P5M_A12TS ix1766 (.Y (nx1765), .A0 (nx136), .A1 (nx128), .B0 (src2_0
                      )) ;
    NOR2_X0P5A_A12TS ix855 (.Y (nx136), .A (nx1495), .B (nx1768)) ;
    NAND2_X0P5A_A12TS ix1769 (.Y (nx1768), .A (alu_op_3), .B (alu_op_2)) ;
    AOI22_X0P5M_A12TS ix1771 (.Y (nx1770), .A0 (src1_1), .A1 (nx114), .B0 (
                      divsrc1_0), .B1 (enable_div)) ;
    NOR2_X0P5A_A12TS ix856 (.Y (nx114), .A (alu_op_1), .B (nx1768)) ;
    AOI221_X0P5M_A12TS ix1774 (.Y (nx1773), .A0 (alu_cy), .A1 (nx971), .B0 (
                       sub_result_0), .B1 (nx94), .C0 (nx76)) ;
    AO21A1AI2_X0P5M_A12TS ix77 (.Y (nx76), .A0 (nx1776), .A1 (nx1778), .B0 (
                          nx1533), .C0 (nx1003)) ;
    NAND2_X0P5A_A12TS ix1777 (.Y (nx1776), .A (nx1643), .B (nx18)) ;
    NAND2_X0P5A_A12TS ix1779 (.Y (nx1778), .A (nx1698), .B (nx6)) ;
    AOI31_X0P5M_A12TS ix857 (.Y (nx1003), .A0 (nx1641), .A1 (src1_7), .A2 (
                      nx1782), .B0 (nx56)) ;
    AOI211_X0P5M_A12TS ix57 (.Y (nx56), .A0 (nx1509), .A1 (nx1537), .B0 (nx44), 
                       .C0 (nx1696)) ;
    NOR2_X0P5A_A12TS ix45 (.Y (nx44), .A (nx1537), .B (nx1509)) ;
    NAND4_X0P5A_A12TS ix858 (.Y (des_acc_1), .A (nx1787), .B (nx1793), .C (
                      nx1795), .D (nx1800)) ;
    AOI22_X0P5M_A12TS ix1788 (.Y (nx1787), .A0 (mulsrc1_1), .A1 (enable_mul), .B0 (
                      nx980), .B1 (nx338)) ;
    XNOR2_X0P5M_A12TS ix859 (.Y (nx980), .A (src1_1), .B (nx1790)) ;
    NOR2_X0P5A_A12TS ix1791 (.Y (nx1790), .A (nx326), .B (srcAc)) ;
    NOR3_X0P5A_A12TS ix339 (.Y (nx338), .A (nx1505), .B (alu_op_3), .C (nx2)) ;
    AOI22_X0P5M_A12TS ix1794 (.Y (nx1793), .A0 (src1_2), .A1 (nx114), .B0 (
                      divsrc1_1), .B1 (enable_div)) ;
    AOI22_X0P5M_A12TS ix1796 (.Y (nx1795), .A0 (src1_0), .A1 (nx978), .B0 (
                      sub_result_1), .B1 (nx94)) ;
    NOR2_X0P5A_A12TS ix860 (.Y (nx978), .A (nx1495), .B (nx1798)) ;
    NAND2_X0P5A_A12TS ix1799 (.Y (nx1798), .A (nx1505), .B (alu_op_3)) ;
    AOI21_X0P5M_A12TS ix1801 (.Y (nx1800), .A0 (des1_1), .A1 (nx977), .B0 (nx974
                      )) ;
    NAND2_X0P5A_A12TS ix271 (.Y (des1_1), .A (nx1803), .B (nx1811)) ;
    AOI222_X0P5M_A12TS ix1804 (.Y (nx1803), .A0 (nx182), .A1 (nx252), .B0 (
                       src2_1), .B1 (nx244), .C0 (nx258), .C1 (nx976)) ;
    NOR2_X0P5A_A12TS ix245 (.Y (nx244), .A (nx1501), .B (nx1768)) ;
    XNOR2_X0P5M_A12TS ix259 (.Y (nx258), .A (src1_0), .B (nx1808)) ;
    XNOR2_X0P5M_A12TS ix1809 (.Y (nx1808), .A (src1_1), .B (alu_cy)) ;
    AOI221_X0P5M_A12TS ix1812 (.Y (nx1811), .A0 (nx188), .A1 (nx222), .B0 (
                       src1_1), .B1 (nx975), .C0 (nx240)) ;
    OAI22_X0P5M_A12TS ix862 (.Y (nx975), .A0 (alu_op_2), .A1 (nx1501), .B0 (
                      nx128), .B1 (nx1815)) ;
    OAI22_X0P5M_A12TS ix241 (.Y (nx240), .A0 (nx1523), .A1 (nx1724), .B0 (src1_1
                      ), .B1 (nx1711)) ;
    OAI21_X0P5M_A12TS ix863 (.Y (nx977), .A0 (alu_op_0), .A1 (nx12), .B0 (nx1819
                      )) ;
    AOI21_X0P5M_A12TS ix1820 (.Y (nx1819), .A0 (alu_op_2), .A1 (alu_op_1), .B0 (
                      nx278)) ;
    NOR2_X0P5A_A12TS ix279 (.Y (nx278), .A (alu_op_1), .B (nx1798)) ;
    AOI211_X0P5M_A12TS ix864 (.Y (nx974), .A0 (nx1687), .A1 (nx1685), .B0 (nx973
                       ), .C0 (nx1696)) ;
    NAND4_X0P5A_A12TS ix487 (.Y (des_acc_2), .A (nx1824), .B (nx1826), .C (
                      nx1828), .D (nx1849)) ;
    AOI22_X0P5M_A12TS ix1825 (.Y (nx1824), .A0 (mulsrc1_2), .A1 (enable_mul), .B0 (
                      divsrc1_2), .B1 (enable_div)) ;
    AOI22_X0P5M_A12TS ix1827 (.Y (nx1826), .A0 (src1_3), .A1 (nx114), .B0 (
                      src1_1), .B1 (nx978)) ;
    AOI22_X0P5M_A12TS ix1829 (.Y (nx1828), .A0 (des1_2), .A1 (nx985), .B0 (
                      sub_result_2), .B1 (nx94)) ;
    NAND2_X0P5A_A12TS ix423 (.Y (des1_2), .A (nx1831), .B (nx1839)) ;
    AOI222_X0P5M_A12TS ix1832 (.Y (nx1831), .A0 (nx981), .A1 (nx252), .B0 (
                       src2_2), .B1 (nx244), .C0 (nx414), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix415 (.Y (nx414), .A (nx1835), .B (nx1837)) ;
    CGENI_X1M_A12TS ix1836 (.CON (nx1835), .A (src1_0), .B (src1_1), .CI (alu_cy
                    )) ;
    XNOR2_X0P5M_A12TS ix1838 (.Y (nx1837), .A (alu_cy), .B (src1_2)) ;
    AOI221_X0P5M_A12TS ix1840 (.Y (nx1839), .A0 (nx358), .A1 (nx222), .B0 (
                       src1_2), .B1 (nx975), .C0 (nx984)) ;
    NOR2_X0P5A_A12TS ix865 (.Y (nx1004), .A (src1_2), .B (src2_2)) ;
    OAI22_X0P5M_A12TS ix866 (.Y (nx984), .A0 (nx1543), .A1 (nx1724), .B0 (src1_2
                      ), .B1 (nx1711)) ;
    NAND2B_X0P7M_A12TS ix867 (.Y (nx985), .AN (nx440), .B (nx1819)) ;
    OAI21_X0P5M_A12TS ix441 (.Y (nx440), .A0 (alu_op_0), .A1 (nx12), .B0 (nx1847
                      )) ;
    AOI31_X0P5M_A12TS ix1850 (.Y (nx1849), .A0 (nx983), .A1 (nx979), .A2 (nx338)
                      , .B0 (nx370)) ;
    OAI21_X0P5M_A12TS ix1855 (.Y (nx1854), .A0 (src1_2), .A1 (src1_1), .B0 (
                      src1_3)) ;
    AOI211_X0P5M_A12TS ix371 (.Y (nx370), .A0 (nx1859), .A1 (nx1862), .B0 (nx982
                       ), .C0 (nx1696)) ;
    XOR2_X0P5M_A12TS ix1863 (.Y (nx1862), .A (nx350), .B (nx1541)) ;
    NOR2_X0P5A_A12TS ix868 (.Y (nx982), .A (nx1862), .B (nx1859)) ;
    NAND4_X0P5A_A12TS ix870 (.Y (des_acc_3), .A (nx1866), .B (nx1868), .C (
                      nx1870), .D (nx1887)) ;
    AOI22_X0P5M_A12TS ix1867 (.Y (nx1866), .A0 (mulsrc1_3), .A1 (enable_mul), .B0 (
                      divsrc1_3), .B1 (enable_div)) ;
    AOI22_X0P5M_A12TS ix1869 (.Y (nx1868), .A0 (src1_4), .A1 (nx114), .B0 (
                      src1_2), .B1 (nx978)) ;
    AOI22_X0P5M_A12TS ix1871 (.Y (nx1870), .A0 (des1_3), .A1 (nx989), .B0 (
                      sub_result_3), .B1 (nx94)) ;
    NAND2_X0P5A_A12TS ix563 (.Y (des1_3), .A (nx1873), .B (nx1882)) ;
    AOI222_X0P5M_A12TS ix1874 (.Y (nx1873), .A0 (nx502), .A1 (nx252), .B0 (
                       src2_3), .B1 (nx244), .C0 (nx988), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix872 (.Y (nx988), .A (nx1877), .B (nx1880)) ;
    CGENI_X1M_A12TS ix1878 (.CON (nx1877), .A (nx410), .B (alu_cy), .CI (src1_2)
                    ) ;
    XNOR2_X0P5M_A12TS ix1881 (.Y (nx1880), .A (alu_cy), .B (src1_3)) ;
    AOI221_X0P5M_A12TS ix1883 (.Y (nx1882), .A0 (nx987), .A1 (nx222), .B0 (
                       src1_3), .B1 (nx975), .C0 (nx536)) ;
    OAI22_X0P5M_A12TS ix537 (.Y (nx536), .A0 (nx1561), .A1 (nx1724), .B0 (src1_3
                      ), .B1 (nx1711)) ;
    NAND2B_X0P7M_A12TS ix873 (.Y (nx989), .AN (nx440), .B (nx1819)) ;
    AOI31_X0P5M_A12TS ix1888 (.Y (nx1887), .A0 (nx1854), .A1 (srcAc), .A2 (nx986
                      ), .B0 (nx520)) ;
    AOI21_X0P5M_A12TS ix874 (.Y (nx986), .A0 (nx1746), .A1 (nx1579), .B0 (nx1890
                      )) ;
    AOI211_X0P5M_A12TS ix521 (.Y (nx520), .A0 (nx1681), .A1 (nx1679), .B0 (nx514
                       ), .C0 (nx1696)) ;
    NAND4_X0P5A_A12TS ix743 (.Y (des_acc_4), .A (nx1894), .B (nx1896), .C (
                      nx1005), .D (nx1926)) ;
    AOI22_X0P5M_A12TS ix1895 (.Y (nx1894), .A0 (mulsrc1_4), .A1 (enable_mul), .B0 (
                      divsrc1_4), .B1 (enable_div)) ;
    AOI22_X0P5M_A12TS ix1897 (.Y (nx1896), .A0 (src1_5), .A1 (nx114), .B0 (
                      src1_3), .B1 (nx978)) ;
    AOI22_X0P5M_A12TS ix875 (.Y (nx1005), .A0 (des1_4), .A1 (nx977), .B0 (
                      sub_result_4), .B1 (nx94)) ;
    OAI211_X1M_A12TS ix699 (.Y (des1_4), .A0 (nx1581), .A1 (nx1901), .B0 (nx1903
                     ), .C0 (nx1914)) ;
    NAND2_X0P5A_A12TS ix1902 (.Y (nx1901), .A (nx1782), .B (nx18)) ;
    AOI21_X0P5M_A12TS ix1904 (.Y (nx1903), .A0 (nx684), .A1 (nx976), .B0 (nx694)
                      ) ;
    XOR2_X0P5M_A12TS ix685 (.Y (nx684), .A (nx1906), .B (nx1911)) ;
    CGENI_X1M_A12TS ix1907 (.CON (nx1906), .A (nx550), .B (alu_cy), .CI (src1_3)
                    ) ;
    XNOR2_X0P5M_A12TS ix1912 (.Y (nx1911), .A (src1_4), .B (alu_cy)) ;
    OAI22_X0P5M_A12TS ix695 (.Y (nx694), .A0 (nx1583), .A1 (nx1724), .B0 (src1_4
                      ), .B1 (nx1711)) ;
    OA21A1OI2_X0P5M_A12TS ix1915 (.Y (nx1914), .A0 (nx664), .A1 (nx252), .B0 (
                          src2_4), .C0 (nx662)) ;
    AOI21_X0P5M_A12TS ix663 (.Y (nx662), .A0 (nx1007), .A1 (nx1922), .B0 (nx1924
                      )) ;
    AOI21_X0P5M_A12TS ix876 (.Y (nx1007), .A0 (nx1537), .A1 (nx244), .B0 (nx975)
                      ) ;
    INV_X0P5B_A12TS ix1925 (.Y (nx1924), .A (src1_4)) ;
    AOI31_X0P5M_A12TS ix1927 (.Y (nx1926), .A0 (nx610), .A1 (nx1743), .A2 (nx338
                      ), .B0 (nx648)) ;
    NAND2B_X0P7M_A12TS ix611 (.Y (nx610), .AN (src1_4), .B (nx1854)) ;
    AOI211_X0P5M_A12TS ix649 (.Y (nx648), .A0 (nx1581), .A1 (nx1668), .B0 (nx642
                       ), .C0 (nx1696)) ;
    NAND4_X0P5A_A12TS ix877 (.Y (des_acc_5), .A (nx1931), .B (nx1933), .C (
                      nx1935), .D (nx1958)) ;
    AOI22_X0P5M_A12TS ix1932 (.Y (nx1931), .A0 (mulsrc1_5), .A1 (enable_mul), .B0 (
                      divsrc1_5), .B1 (enable_div)) ;
    AOI22_X0P5M_A12TS ix1934 (.Y (nx1933), .A0 (src1_6), .A1 (nx114), .B0 (
                      src1_4), .B1 (nx978)) ;
    AOI22_X0P5M_A12TS ix1936 (.Y (nx1935), .A0 (des1_5), .A1 (nx977), .B0 (
                      sub_result_5), .B1 (nx94)) ;
    OAI211_X1M_A12TS ix831 (.Y (des1_5), .A0 (nx1938), .A1 (nx1945), .B0 (nx1947
                     ), .C0 (nx1950)) ;
    XNOR2_X0P5M_A12TS ix1939 (.Y (nx1938), .A (nx1940), .B (nx1943)) ;
    CGENI_X1M_A12TS ix1941 (.CON (nx1940), .A (nx680), .B (src1_4), .CI (alu_cy)
                    ) ;
    XNOR2_X0P5M_A12TS ix1944 (.Y (nx1943), .A (src1_5), .B (alu_cy)) ;
    NAND2_X0P5A_A12TS ix1946 (.Y (nx1945), .A (nx972), .B (nx1641)) ;
    AOI22_X0P5M_A12TS ix1948 (.Y (nx1947), .A0 (nx744), .A1 (nx252), .B0 (src2_5
                      ), .B1 (nx664)) ;
    AOI221_X0P5M_A12TS ix1951 (.Y (nx1950), .A0 (nx750), .A1 (nx222), .B0 (
                       src1_5), .B1 (nx990), .C0 (nx993)) ;
    OAI22_X0P5M_A12TS ix878 (.Y (nx993), .A0 (nx1595), .A1 (nx1724), .B0 (src1_5
                      ), .B1 (nx1711)) ;
    AOI21_X0P5M_A12TS ix1959 (.Y (nx1958), .A0 (nx338), .A1 (nx786), .B0 (nx762)
                      ) ;
    XNOR2_X0P5M_A12TS ix787 (.Y (nx786), .A (nx776), .B (nx992)) ;
    OAI21_X0P5M_A12TS ix777 (.Y (nx776), .A0 (src1_5), .A1 (nx768), .B0 (nx1963)
                      ) ;
    NOR2_X0P5A_A12TS ix769 (.Y (nx768), .A (src1_5), .B (nx1743)) ;
    NAND3_X0P5A_A12TS ix880 (.Y (nx992), .A (nx1854), .B (nx1537), .C (nx1736)
                      ) ;
    AOI211_X0P5M_A12TS ix763 (.Y (nx762), .A0 (nx1968), .A1 (nx1970), .B0 (nx991
                       ), .C0 (nx1696)) ;
    XNOR2_X0P5M_A12TS ix1971 (.Y (nx1970), .A (nx1583), .B (nx1593)) ;
    NOR2_X0P5A_A12TS ix881 (.Y (nx991), .A (nx1970), .B (nx1968)) ;
    NAND4_X0P5A_A12TS ix882 (.Y (des_acc_6), .A (nx1974), .B (nx1976), .C (
                      nx1978), .D (nx1997)) ;
    AOI22_X0P5M_A12TS ix1975 (.Y (nx1974), .A0 (mulsrc1_6), .A1 (enable_mul), .B0 (
                      divsrc1_6), .B1 (enable_div)) ;
    AOI22_X0P5M_A12TS ix1977 (.Y (nx1976), .A0 (src1_7), .A1 (nx114), .B0 (
                      src1_5), .B1 (nx978)) ;
    AOI22_X0P5M_A12TS ix1979 (.Y (nx1978), .A0 (des1_6), .A1 (nx977), .B0 (
                      sub_result_6), .B1 (nx94)) ;
    OAI211_X1M_A12TS ix963 (.Y (des1_6), .A0 (nx1981), .A1 (nx1945), .B0 (nx1988
                     ), .C0 (nx1991)) ;
    XNOR2_X0P5M_A12TS ix1982 (.Y (nx1981), .A (nx1983), .B (nx1986)) ;
    CGENI_X1M_A12TS ix1984 (.CON (nx1983), .A (nx814), .B (src1_5), .CI (alu_cy)
                    ) ;
    XNOR2_X0P5M_A12TS ix1987 (.Y (nx1986), .A (src1_6), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix1989 (.Y (nx1988), .A0 (nx994), .A1 (nx252), .B0 (src2_6
                      ), .B1 (nx664)) ;
    AOI221_X0P5M_A12TS ix1992 (.Y (nx1991), .A0 (nx876), .A1 (nx222), .B0 (
                       src1_6), .B1 (nx990), .C0 (nx936)) ;
    NOR2_X0P5A_A12TS ix1995 (.Y (nx1994), .A (src1_6), .B (src2_6)) ;
    OAI22_X0P5M_A12TS ix937 (.Y (nx936), .A0 (nx1607), .A1 (nx1724), .B0 (src1_6
                      ), .B1 (nx1711)) ;
    OA21A1OI2_X0P5M_A12TS ix1998 (.Y (nx1997), .A0 (nx916), .A1 (nx900), .B0 (
                          nx338), .C0 (nx888)) ;
    AOI211_X0P5M_A12TS ix917 (.Y (nx916), .A0 (nx2000), .A1 (nx1008), .B0 (
                       nx2006), .C0 (nx910)) ;
    AOI21_X0P5M_A12TS ix884 (.Y (nx1008), .A0 (src1_5), .A1 (src1_6), .B0 (
                      nx2004)) ;
    NOR2_X0P5A_A12TS ix2005 (.Y (nx2004), .A (src1_6), .B (src1_5)) ;
    NOR3_X0P5A_A12TS ix911 (.Y (nx910), .A (src1_5), .B (src1_6), .C (nx1743)) ;
    AND4_X0P5M_A12TS ix901 (.Y (nx900), .A (nx1854), .B (src1_6), .C (nx1537), .D (
                     nx1736)) ;
    AOI211_X0P5M_A12TS ix889 (.Y (nx888), .A0 (nx1663), .A1 (nx1661), .B0 (nx882
                       ), .C0 (nx1696)) ;
    NAND4_X0P5A_A12TS ix1161 (.Y (des_acc_7), .A (nx2013), .B (nx2016), .C (
                      nx2033), .D (nx2035)) ;
    NAND2_X0P5A_A12TS ix2014 (.Y (nx2013), .A (nx1152), .B (nx50)) ;
    XOR2_X0P5M_A12TS ix1153 (.Y (nx1152), .A (nx1651), .B (nx1627)) ;
    MXIT2_X0P5M_A12TS ix2017 (.Y (nx2016), .A (nx1118), .B (nx1140), .S0 (
                      alu_op_0)) ;
    OAI222_X0P5M_A12TS ix1119 (.Y (nx1118), .A0 (src1_7), .A1 (nx1763), .B0 (
                       nx1627), .B1 (nx2019), .C0 (nx2021), .C1 (nx2028)) ;
    XNOR2_X0P5M_A12TS ix2022 (.Y (nx2021), .A (nx2023), .B (nx2026)) ;
    CGENI_X1M_A12TS ix2024 (.CON (nx2023), .A (nx995), .B (src1_6), .CI (alu_cy)
                    ) ;
    XNOR2_X0P5M_A12TS ix2027 (.Y (nx2026), .A (src1_7), .B (alu_cy)) ;
    OAI222_X0P5M_A12TS ix1141 (.Y (nx1140), .A0 (nx1629), .A1 (nx1763), .B0 (
                       nx2028), .B1 (nx2031), .C0 (nx1689), .C1 (nx2019)) ;
    MXIT2_X0P5M_A12TS ix2032 (.Y (nx2031), .A (src1_7), .B (src2_7), .S0 (alu_cy
                      )) ;
    AOI22_X0P5M_A12TS ix2034 (.Y (nx2033), .A0 (mulsrc1_7), .A1 (enable_mul), .B0 (
                      divsrc1_7), .B1 (enable_div)) ;
    AOI221_X0P5M_A12TS ix2036 (.Y (nx2035), .A0 (src1_7), .A1 (nx22), .B0 (
                       sub_result_7), .B1 (nx94), .C0 (nx1052)) ;
    OAI21_X0P5M_A12TS ix1053 (.Y (nx1052), .A0 (nx1768), .A1 (nx2038), .B0 (
                      nx2040)) ;
    AOI22_X0P5M_A12TS ix2039 (.Y (nx2038), .A0 (src1_0), .A1 (nx18), .B0 (alu_cy
                      ), .B1 (nx1698)) ;
    AOI31_X0P5M_A12TS ix2041 (.Y (nx2040), .A0 (nx1782), .A1 (alu_op_1), .A2 (
                      src1_6), .B0 (nx1048)) ;
    AOI21_X0P5M_A12TS ix1049 (.Y (nx1048), .A0 (nx2043), .A1 (nx2045), .B0 (
                      nx1778)) ;
    NAND4_X0P5A_A12TS ix2044 (.Y (nx2043), .A (nx1854), .B (nx1537), .C (src1_7)
                      , .D (nx2004)) ;
    OAI211_X0P5M_A12TS ix2046 (.Y (nx2045), .A0 (nx910), .A1 (nx1028), .B0 (
                       nx992), .C0 (nx2048)) ;
    INV_X0P5B_A12TS ix1029 (.Y (nx1028), .A (nx1739)) ;
    NAND4_X0P5A_A12TS ix1221 (.Y (des2_0), .A (nx2051), .B (nx2061), .C (nx2063)
                      , .D (nx2066)) ;
    AOI222_X0P5M_A12TS ix2052 (.Y (nx2051), .A0 (mulsrc2_0), .A1 (enable_mul), .B0 (
                       src1_0), .B1 (nx244), .C0 (nx1212), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix1213 (.Y (nx1212), .A (nx1009), .B (nx2059)) ;
    CGENI_X1M_A12TS ix885 (.CON (nx1009), .A (nx1104), .B (src1_7), .CI (alu_cy)
                    ) ;
    XNOR2_X0P5M_A12TS ix2060 (.Y (nx2059), .A (src2_0), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2062 (.Y (nx2061), .A0 (divsrc2_0), .A1 (enable_div), .B0 (
                      src2_0), .B1 (nx22)) ;
    NAND2_X0P5A_A12TS ix2064 (.Y (nx2063), .A (src1_4), .B (nx1184)) ;
    NOR2_X0P5A_A12TS ix1185 (.Y (nx1184), .A (nx1501), .B (nx1798)) ;
    OAI211_X0P5M_A12TS ix2067 (.Y (nx2066), .A0 (nx1172), .A1 (src3_0), .B0 (
                       nx2068), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2069 (.Y (nx2068), .A (src3_0), .B (nx1172)) ;
    NAND4_X0P5A_A12TS ix1267 (.Y (des2_1), .A (nx2071), .B (nx2079), .C (nx2081)
                      , .D (nx2083)) ;
    AOI222_X0P5M_A12TS ix2072 (.Y (nx2071), .A0 (mulsrc2_1), .A1 (enable_mul), .B0 (
                       src1_1), .B1 (nx244), .C0 (nx1258), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix1259 (.Y (nx1258), .A (nx2074), .B (nx2077)) ;
    CGENI_X1M_A12TS ix2075 (.CON (nx2074), .A (nx1208), .B (src2_0), .CI (alu_cy
                    )) ;
    XNOR2_X0P5M_A12TS ix2078 (.Y (nx2077), .A (src2_1), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2080 (.Y (nx2079), .A0 (divsrc2_1), .A1 (enable_div), .B0 (
                      src2_1), .B1 (nx22)) ;
    NAND2_X0P5A_A12TS ix2082 (.Y (nx2081), .A (src1_5), .B (nx1184)) ;
    OAI211_X0P5M_A12TS ix2084 (.Y (nx2083), .A0 (nx1176), .A1 (src3_1), .B0 (
                       nx2086), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2087 (.Y (nx2086), .A (src3_1), .B (nx1176)) ;
    NAND4_X0P5A_A12TS ix886 (.Y (des2_2), .A (nx2089), .B (nx2099), .C (nx2101)
                      , .D (nx2103)) ;
    AOI222_X0P5M_A12TS ix2090 (.Y (nx2089), .A0 (mulsrc2_2), .A1 (enable_mul), .B0 (
                       src1_2), .B1 (nx244), .C0 (nx1304), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix1305 (.Y (nx1304), .A (nx2092), .B (nx2097)) ;
    CGENI_X1M_A12TS ix2093 (.CON (nx2092), .A (nx998), .B (src2_1), .CI (alu_cy)
                    ) ;
    XNOR2_X0P5M_A12TS ix2098 (.Y (nx2097), .A (src2_2), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2100 (.Y (nx2099), .A0 (divsrc2_2), .A1 (enable_div), .B0 (
                      src2_2), .B1 (nx22)) ;
    NAND2_X0P5A_A12TS ix2102 (.Y (nx2101), .A (src1_6), .B (nx1184)) ;
    OAI211_X0P5M_A12TS ix2104 (.Y (nx2103), .A0 (nx1224), .A1 (src3_2), .B0 (
                       nx2108), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2109 (.Y (nx2108), .A (src3_2), .B (nx1224)) ;
    NAND4_X0P5A_A12TS ix1359 (.Y (des2_3), .A (nx2111), .B (nx2121), .C (nx2123)
                      , .D (nx2125)) ;
    AOI222_X0P5M_A12TS ix2112 (.Y (nx2111), .A0 (mulsrc2_3), .A1 (enable_mul), .B0 (
                       src1_3), .B1 (nx244), .C0 (nx1350), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix1351 (.Y (nx1350), .A (nx2114), .B (nx2119)) ;
    CGENI_X1M_A12TS ix2115 (.CON (nx2114), .A (nx1300), .B (src2_2), .CI (alu_cy
                    )) ;
    XNOR2_X0P5M_A12TS ix2120 (.Y (nx2119), .A (src2_3), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2122 (.Y (nx2121), .A0 (divsrc2_3), .A1 (enable_div), .B0 (
                      src2_3), .B1 (nx22)) ;
    NAND2_X0P5A_A12TS ix2124 (.Y (nx2123), .A (src1_7), .B (nx1184)) ;
    OAI211_X0P5M_A12TS ix2126 (.Y (nx2125), .A0 (nx1270), .A1 (src3_3), .B0 (
                       nx2130), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2131 (.Y (nx2130), .A (src3_3), .B (nx1270)) ;
    NAND4_X0P5A_A12TS ix1411 (.Y (des2_4), .A (nx2133), .B (nx2142), .C (nx2144)
                      , .D (nx2146)) ;
    AOI222_X0P5M_A12TS ix2134 (.Y (nx2133), .A0 (mulsrc2_4), .A1 (enable_mul), .B0 (
                       src2_4), .B1 (nx1386), .C0 (nx1402), .C1 (nx976)) ;
    OAI21_X0P5M_A12TS ix1387 (.Y (nx1386), .A0 (alu_cy), .A1 (nx1917), .B0 (
                      nx1776)) ;
    XOR2_X0P5M_A12TS ix1406 (.Y (nx1402), .A (nx2137), .B (nx2140)) ;
    CGENI_X1M_A12TS ix2138 (.CON (nx2137), .A (nx1346), .B (src2_3), .CI (alu_cy
                    )) ;
    XNOR2_X0P5M_A12TS ix2141 (.Y (nx2140), .A (src2_4), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2143 (.Y (nx2142), .A0 (divsrc2_4), .A1 (enable_div), .B0 (
                      src1_4), .B1 (nx664)) ;
    NAND2_X0P5A_A12TS ix2145 (.Y (nx2144), .A (src1_0), .B (nx971)) ;
    OAI211_X0P5M_A12TS ix2147 (.Y (nx2146), .A0 (nx1316), .A1 (src3_4), .B0 (
                       nx2151), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2152 (.Y (nx2151), .A (src3_4), .B (nx1316)) ;
    NAND4_X0P5A_A12TS ix1457 (.Y (des2_5), .A (nx2154), .B (nx2164), .C (nx2166)
                      , .D (nx2168)) ;
    AOI222_X0P5M_A12TS ix2155 (.Y (nx2154), .A0 (mulsrc2_5), .A1 (enable_mul), .B0 (
                       src2_5), .B1 (nx1386), .C0 (nx1448), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix1449 (.Y (nx1448), .A (nx2157), .B (nx2162)) ;
    CGENI_X1M_A12TS ix2158 (.CON (nx2157), .A (nx1398), .B (src2_4), .CI (alu_cy
                    )) ;
    XNOR2_X0P5M_A12TS ix2163 (.Y (nx2162), .A (src2_5), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2165 (.Y (nx2164), .A0 (divsrc2_5), .A1 (enable_div), .B0 (
                      src1_5), .B1 (nx664)) ;
    NAND2_X0P5A_A12TS ix2167 (.Y (nx2166), .A (src1_1), .B (nx971)) ;
    OAI211_X0P5M_A12TS ix2169 (.Y (nx2168), .A0 (nx1362), .A1 (src3_5), .B0 (
                       nx2173), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2174 (.Y (nx2173), .A (src3_5), .B (nx1362)) ;
    NAND4_X0P5A_A12TS ix887 (.Y (des2_6), .A (nx2176), .B (nx2186), .C (nx1010)
                      , .D (nx2190)) ;
    AOI222_X0P5M_A12TS ix2177 (.Y (nx2176), .A0 (mulsrc2_6), .A1 (enable_mul), .B0 (
                       src2_6), .B1 (nx1386), .C0 (nx1494), .C1 (nx976)) ;
    XOR2_X0P5M_A12TS ix1495 (.Y (nx1494), .A (nx2179), .B (nx2184)) ;
    CGENI_X1M_A12TS ix2180 (.CON (nx2179), .A (nx999), .B (src2_5), .CI (alu_cy)
                    ) ;
    XNOR2_X0P5M_A12TS ix2185 (.Y (nx2184), .A (src2_6), .B (alu_cy)) ;
    AOI22_X0P5M_A12TS ix2187 (.Y (nx2186), .A0 (divsrc2_6), .A1 (enable_div), .B0 (
                      src1_6), .B1 (nx664)) ;
    NAND2_X0P5A_A12TS ix888 (.Y (nx1010), .A (src1_2), .B (nx971)) ;
    OAI211_X0P5M_A12TS ix2191 (.Y (nx2190), .A0 (nx1414), .A1 (src3_6), .B0 (
                       nx2195), .C0 (nx50)) ;
    NAND2_X0P5A_A12TS ix2196 (.Y (nx2195), .A (src3_6), .B (nx1414)) ;
    NAND3_X0P5A_A12TS ix1543 (.Y (des2_7), .A (nx2198), .B (nx2207), .C (nx2209)
                      ) ;
    AOI222_X0P5M_A12TS ix2199 (.Y (nx2198), .A0 (src2_7), .A1 (nx1386), .B0 (
                       nx1520), .B1 (nx50), .C0 (nx1534), .C1 (nx976)) ;
    XNOR2_X0P5M_A12TS ix1521 (.Y (nx1520), .A (src3_7), .B (nx2195)) ;
    XNOR3_X0P5M_A12TS ix1535 (.Y (nx1534), .A (nx2202), .B (src2_7), .C (alu_cy)
                      ) ;
    CGENI_X1M_A12TS ix2203 (.CON (nx2202), .A (nx1490), .B (src2_6), .CI (alu_cy
                    )) ;
    AOI22_X0P5M_A12TS ix2208 (.Y (nx2207), .A0 (mulsrc2_7), .A1 (enable_mul), .B0 (
                      src1_7), .B1 (nx664)) ;
    AOI22_X0P5M_A12TS ix2210 (.Y (nx2209), .A0 (divsrc2_7), .A1 (enable_div), .B0 (
                      src1_3), .B1 (nx971)) ;
    AO1B2_X0P5M_A12TS ix890 (.Y (des1_7), .A0N (nx2016), .B0 (src1_7), .B1 (
                      nx975)) ;
    INV_X0P5B_A12TS ix1491 (.Y (nx1490), .A (nx2179)) ;
    INV_X0P5B_A12TS ix891 (.Y (nx999), .A (nx2157)) ;
    INV_X0P5B_A12TS ix1415 (.Y (nx1414), .A (nx2173)) ;
    INV_X0P5B_A12TS ix1399 (.Y (nx1398), .A (nx2137)) ;
    INV_X0P5B_A12TS ix1363 (.Y (nx1362), .A (nx2151)) ;
    INV_X0P5B_A12TS ix1347 (.Y (nx1346), .A (nx2114)) ;
    INV_X0P5B_A12TS ix1317 (.Y (nx1316), .A (nx2130)) ;
    INV_X0P5B_A12TS ix1301 (.Y (nx1300), .A (nx2092)) ;
    INV_X0P5B_A12TS ix1271 (.Y (nx1270), .A (nx2108)) ;
    INV_X0P5B_A12TS ix892 (.Y (nx998), .A (nx2074)) ;
    INV_X0P5B_A12TS ix1225 (.Y (nx1224), .A (nx2086)) ;
    INV_X0P5B_A12TS ix1209 (.Y (nx1208), .A (nx1009)) ;
    INV_X0P5B_A12TS ix1177 (.Y (nx1176), .A (nx2068)) ;
    INV_X0P5B_A12TS ix1715 (.Y (nx1714), .A (nx1172)) ;
    INV_X0P5B_A12TS ix1105 (.Y (nx1104), .A (nx2023)) ;
    INV_X0P5B_A12TS ix2049 (.Y (nx2048), .A (nx1032)) ;
    INV_X0P5B_A12TS ix894 (.Y (nx995), .A (nx1983)) ;
    INV_X0P5B_A12TS ix895 (.Y (nx876), .A (nx1605)) ;
    INV_X0P5B_A12TS ix896 (.Y (nx994), .A (nx1994)) ;
    INV_X0P5B_A12TS ix815 (.Y (nx814), .A (nx1940)) ;
    INV_X0P5B_A12TS ix2007 (.Y (nx2006), .A (nx992)) ;
    INV_X0P5B_A12TS ix2001 (.Y (nx2000), .A (nx768)) ;
    INV_X0P5B_A12TS ix1664 (.Y (nx1663), .A (nx991)) ;
    INV_X0P5B_A12TS ix751 (.Y (nx750), .A (nx1593)) ;
    INV_X0P5B_A12TS ix745 (.Y (nx744), .A (nx1657)) ;
    INV_X0P5B_A12TS ix681 (.Y (nx680), .A (nx1906)) ;
    INV_X0P5B_A12TS ix897 (.Y (nx990), .A (nx1007)) ;
    INV_X0P5B_A12TS ix1969 (.Y (nx1968), .A (nx642)) ;
    INV_X0P5B_A12TS ix551 (.Y (nx550), .A (nx1877)) ;
    INV_X0P5B_A12TS ix898 (.Y (nx987), .A (nx1559)) ;
    INV_X0P5B_A12TS ix503 (.Y (nx502), .A (nx1676)) ;
    INV_X0P5B_A12TS ix411 (.Y (nx410), .A (nx1835)) ;
    INV_X0P5B_A12TS ix1682 (.Y (nx1681), .A (nx982)) ;
    INV_X0P5B_A12TS ix359 (.Y (nx358), .A (nx1541)) ;
    INV_X0P5B_A12TS ix899 (.Y (nx981), .A (nx1004)) ;
    INV_X0P5B_A12TS ix1891 (.Y (nx1890), .A (nx338)) ;
    INV_X0P5B_A12TS ix900 (.Y (nx979), .A (nx1790)) ;
    INV_X0P5B_A12TS ix327 (.Y (nx326), .A (nx1854)) ;
    INV_X0P5B_A12TS ix902 (.Y (nx976), .A (nx1945)) ;
    INV_X0P5B_A12TS ix1923 (.Y (nx1922), .A (nx252)) ;
    INV_X0P5B_A12TS ix1918 (.Y (nx1917), .A (nx244)) ;
    INV_X0P5B_A12TS ix223 (.Y (nx222), .A (nx1901)) ;
    INV_X0P5B_A12TS ix1860 (.Y (nx1859), .A (nx973)) ;
    INV_X0P5B_A12TS ix189 (.Y (nx188), .A (nx1521)) ;
    INV_X0P5B_A12TS ix183 (.Y (nx182), .A (nx1674)) ;
    INV_X0P5B_A12TS ix2029 (.Y (nx2028), .A (nx136)) ;
    INV_X0P5B_A12TS ix2020 (.Y (nx2019), .A (nx128)) ;
    INV_X0P5B_A12TS ix903 (.Y (nx972), .A (nx1768)) ;
    INV_X0P5B_A12TS ix95 (.Y (nx94), .A (nx1639)) ;
    INV_X0P5B_A12TS ix1783 (.Y (nx1782), .A (nx970)) ;
    INV_X0P5B_A12TS ix61 (.Y (nx60), .A (nx1641)) ;
    INV_X0P5B_A12TS ix1697 (.Y (nx1696), .A (nx50)) ;
    INV_X0P5B_A12TS ix1688 (.Y (nx1687), .A (nx44)) ;
    INV_X0P5B_A12TS ix41 (.Y (nx40), .A (nx1509)) ;
    INV_X0P5B_A12TS ix23 (.Y (nx22), .A (nx1776)) ;
    INV_X0P5B_A12TS ix13 (.Y (nx12), .A (nx1643)) ;
    INV_X0P5B_A12TS ix904 (.Y (nx969), .A (nx1778)) ;
    INV_X0P5B_A12TS ix1699 (.Y (nx1698), .A (nx2)) ;
    AND2_X0P5M_A12TS ix119 (.Y (enable_div), .A (nx6), .B (nx18)) ;
    NAND2B_X0P7M_A12TS ix299 (.Y (nx298), .AN (nx80), .B (nx1519)) ;
    NAND2B_X0P7M_A12TS ix459 (.Y (nx458), .AN (nx298), .B (nx1539)) ;
    NAND2B_X0P7M_A12TS ix581 (.Y (nx580), .AN (nx458), .B (nx1557)) ;
    NAND2B_X0P7M_A12TS ix837 (.Y (nx836), .AN (nx714), .B (nx1591)) ;
    NAND2B_X0P7M_A12TS ix979 (.Y (nx997), .AN (nx836), .B (nx1603)) ;
    NAND2B_X0P7M_A12TS ix1725 (.Y (nx1724), .AN (nx1501), .B (nx6)) ;
    NOR2B_X0P7M_A12TS ix1033 (.Y (nx1032), .AN (nx910), .B (nx1739)) ;
    AND2_X0P5M_A12TS ix1816 (.Y (nx1815), .A (nx970), .B (alu_op_1)) ;
    NAND4B_X0P5M_A12TS ix1848 (.Y (nx1847), .AN (alu_op_3), .B (alu_op_0), .C (
                       nx1790), .D (alu_op_2)) ;
    AO21_X0P5M_A12TS ix906 (.Y (nx983), .A0 (src1_1), .A1 (src1_2), .B0 (nx1746)
                     ) ;
    AND2_X0P5M_A12TS ix907 (.Y (nx664), .A (alu_cy), .B (nx244)) ;
    NAND2B_X0P7M_A12TS ix1964 (.Y (nx1963), .AN (nx1743), .B (src1_5)) ;
    AO21_X0P5M_A12TS ix1165 (.Y (des1_0), .A0 (src1_0), .A1 (nx975), .B0 (nx168)
                     ) ;
    NOR2_X0P5A_A12TS ix340 (.Y (nx339), .A (nx341), .B (wr_addr_7)) ;
    INV_X0P5B_A12TS ix342 (.Y (nx341), .A (bit_addr_r)) ;
    DFFRPQ_X0P5M_A12TS reg_bit_addr_r (.Q (bit_addr_r), .CK (wb_clk_i), .D (
                       bit_addr), .R (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix352 (.Y (nx351), .A (nx353), .B (rd_addr_7)) ;
    INV_X0P5B_A12TS ix354 (.Y (nx353), .A (bit_addr)) ;
    NAND4_X0P5A_A12TS ix360 (.Y (NOT_rd_en), .A (nx1055), .B (nx395), .C (nx401)
                      , .D (nx1056)) ;
    NOR3_X0P5A_A12TS ix1011 (.Y (nx1055), .A (nx363), .B (nx88), .C (nx106)) ;
    NAND3_X0P5A_A12TS ix364 (.Y (nx363), .A (nx365), .B (wr_dup_1054), .C (nx373
                      )) ;
    AOI22_X0P5M_A12TS ix368 (.Y (nx367), .A0 (nx353), .A1 (rd_addr_1), .B0 (
                      rd_addr_4), .B1 (nx351)) ;
    INV_X0P5B_A12TS ix1012 (.Y (wr_addr_m_1), .A (nx371)) ;
    AOI22_X0P5M_A12TS ix372 (.Y (nx371), .A0 (wr_addr_1), .A1 (nx341), .B0 (
                      wr_addr_4), .B1 (nx339)) ;
    AOI22_X0P5M_A12TS ix376 (.Y (nx375), .A0 (nx353), .A1 (rd_addr_0), .B0 (
                      rd_addr_3), .B1 (nx351)) ;
    INV_X0P5B_A12TS ix1014 (.Y (wr_addr_m_0), .A (nx379)) ;
    AOI22_X0P5M_A12TS ix380 (.Y (nx379), .A0 (wr_addr_0), .A1 (nx341), .B0 (
                      wr_addr_3), .B1 (nx339)) ;
    AOI22_X0P5M_A12TS ix384 (.Y (nx383), .A0 (nx353), .A1 (rd_addr_2), .B0 (
                      rd_addr_5), .B1 (nx351)) ;
    INV_X0P5B_A12TS ix17 (.Y (wr_addr_m_2), .A (nx387)) ;
    AOI22_X0P5M_A12TS ix388 (.Y (nx387), .A0 (wr_addr_2), .A1 (nx341), .B0 (
                      wr_addr_5), .B1 (nx339)) ;
    XNOR2_X0P5M_A12TS ix107 (.Y (nx106), .A (nx391), .B (wr_addr_m_3)) ;
    MXIT2_X0P5M_A12TS ix392 (.Y (nx391), .A (rd_addr_3), .B (rd_addr_6), .S0 (
                      nx351)) ;
    MXT2_X0P5M_A12TS ix105 (.Y (wr_addr_m_3), .A (wr_addr_3), .B (wr_addr_6), .S0 (
                     nx339)) ;
    XOR2_X0P5M_A12TS ix396 (.Y (nx395), .A (nx397), .B (wr_addr_m_4)) ;
    NAND2_X0P5A_A12TS ix398 (.Y (nx397), .A (rd_addr_4), .B (nx20)) ;
    XOR2_X0P5M_A12TS ix402 (.Y (nx401), .A (nx403), .B (wr_addr_m_5)) ;
    NOR2_X0P5A_A12TS ix404 (.Y (nx403), .A (nx351), .B (rd_addr_5)) ;
    OR2_X0P5M_A12TS ix1015 (.Y (wr_addr_m_5), .A (nx339), .B (wr_addr_5)) ;
    NOR2_X0P5A_A12TS ix1016 (.Y (nx1056), .A (nx142), .B (nx144)) ;
    XNOR2_X0P5M_A12TS ix143 (.Y (nx142), .A (nx409), .B (wr_addr_m_6)) ;
    NAND2_X0P5A_A12TS ix410 (.Y (nx409), .A (rd_addr_6), .B (nx20)) ;
    XOR2_X0P5M_A12TS ix145 (.Y (nx144), .A (rd_addr_7), .B (wr_addr_7)) ;
    OAI211_X0P5M_A12TS ix317 (.Y (wr_data_m_0), .A0 (nx302), .A1 (nx423), .B0 (
                       nx427), .C0 (nx447)) ;
    DFFRPQ_X0P5M_A12TS reg_bit_select_1 (.Q (bit_select_1), .CK (wb_clk_i), .D (
                       rd_addr_1), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_bit_select_2 (.Q (bit_select_2), .CK (wb_clk_i), .D (
                       rd_addr_2), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix424 (.Y (nx423), .A (desCy), .B (nx192)) ;
    NOR2_X0P5A_A12TS ix193 (.Y (nx192), .A (bit_select_0), .B (nx341)) ;
    DFFRPQ_X0P5M_A12TS reg_bit_select_0 (.Q (bit_select_0), .CK (wb_clk_i), .D (
                       rd_addr_0), .R (wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix428 (.Y (nx427), .A0 (nx302), .A1 (bit_select_0), .B0 (
                       ram_data_0), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix325 (.Y (ram_data_0), .A (rd_data_m_0), .B (wr_data_r_0)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_0 (.Q (wr_data_r_0), .CK (wb_clk_i), .D (
                       wr_data_m_0), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_rd_en_r (.Q (rd_en_r), .CK (wb_clk_i), .D (nx154), .R (
                       wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix448 (.Y (nx447), .A (des1_0), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix1017 (.Y (wr_data_m_1), .A0 (nx302), .A1 (nx451), .B0 (
                       nx453), .C0 (nx1059)) ;
    NAND3_X0P5A_A12TS ix452 (.Y (nx451), .A (desCy), .B (bit_select_0), .C (
                      bit_addr_r)) ;
    OAI211_X0P5M_A12TS ix454 (.Y (nx453), .A0 (nx302), .A1 (nx455), .B0 (
                       ram_data_1), .C0 (bit_addr_r)) ;
    INV_X0P5B_A12TS ix456 (.Y (nx455), .A (bit_select_0)) ;
    MXT2_X0P5M_A12TS ix1018 (.Y (ram_data_1), .A (rd_data_m_1), .B (wr_data_r_1)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_1 (.Q (wr_data_r_1), .CK (wb_clk_i), .D (
                       wr_data_m_1), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix462 (.Y (nx1059), .A (des1_1), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix281 (.Y (wr_data_m_2), .A0 (nx1058), .A1 (nx423), .B0 (
                       nx467), .C0 (nx471)) ;
    OAI211_X0P5M_A12TS ix468 (.Y (nx467), .A0 (nx1058), .A1 (bit_select_0), .B0 (
                       ram_data_2), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix1019 (.Y (ram_data_2), .A (rd_data_m_2), .B (wr_data_r_2)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_2 (.Q (wr_data_r_2), .CK (wb_clk_i), .D (
                       wr_data_m_2), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix472 (.Y (nx471), .A (des1_2), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix1020 (.Y (wr_data_m_3), .A0 (nx1058), .A1 (nx451), .B0 (
                       nx475), .C0 (nx481)) ;
    OAI211_X0P5M_A12TS ix476 (.Y (nx475), .A0 (nx1058), .A1 (nx455), .B0 (
                       ram_data_3), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix439 (.Y (ram_data_3), .A (rd_data_m_3), .B (wr_data_r_3)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_3 (.Q (wr_data_r_3), .CK (wb_clk_i), .D (
                       wr_data_m_3), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix482 (.Y (nx481), .A (des1_3), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix1022 (.Y (wr_data_m_4), .A0 (nx226), .A1 (nx423), .B0 (
                       nx487), .C0 (nx491)) ;
    OAI211_X0P5M_A12TS ix488 (.Y (nx487), .A0 (nx226), .A1 (bit_select_0), .B0 (
                       ram_data_4), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix249 (.Y (ram_data_4), .A (rd_data_m_4), .B (wr_data_r_4)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_4 (.Q (wr_data_r_4), .CK (wb_clk_i), .D (
                       wr_data_m_4), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix492 (.Y (nx491), .A (des1_4), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix395 (.Y (wr_data_m_5), .A0 (nx226), .A1 (nx451), .B0 (
                       nx1060), .C0 (nx498)) ;
    OAI211_X0P5M_A12TS ix1023 (.Y (nx1060), .A0 (nx226), .A1 (nx455), .B0 (
                       ram_data_5), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix403 (.Y (ram_data_5), .A (rd_data_m_5), .B (wr_data_r_5)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_5 (.Q (wr_data_r_5), .CK (wb_clk_i), .D (
                       wr_data_m_5), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix499 (.Y (nx498), .A (des1_5), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix203 (.Y (wr_data_m_6), .A0 (nx1057), .A1 (nx423), .B0 (
                       nx1061), .C0 (nx1062)) ;
    NAND2_X0P5A_A12TS ix1024 (.Y (nx1057), .A (bit_select_1), .B (bit_select_2)
                      ) ;
    OAI211_X0P5M_A12TS ix1025 (.Y (nx1061), .A0 (nx1057), .A1 (bit_select_0), .B0 (
                       ram_data_6), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix211 (.Y (ram_data_6), .A (rd_data_m_6), .B (wr_data_r_6)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_6 (.Q (wr_data_r_6), .CK (wb_clk_i), .D (
                       wr_data_m_6), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix1026 (.Y (nx1062), .A (des1_6), .B (nx341)) ;
    OAI211_X0P5M_A12TS ix361 (.Y (wr_data_m_7), .A0 (nx1057), .A1 (nx451), .B0 (
                       nx509), .C0 (nx513)) ;
    OAI211_X0P5M_A12TS ix510 (.Y (nx509), .A0 (nx1057), .A1 (nx455), .B0 (
                       ram_data_7), .C0 (bit_addr_r)) ;
    MXT2_X0P5M_A12TS ix1027 (.Y (ram_data_7), .A (rd_data_m_7), .B (wr_data_r_7)
                     , .S0 (rd_en_r)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_data_r_7 (.Q (wr_data_r_7), .CK (wb_clk_i), .D (
                       wr_data_m_7), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix514 (.Y (nx513), .A (des1_7), .B (nx341)) ;
    AO21A1AI2_X0P5M_A12TS ix1028 (.Y (bit_data), .A0 (nx531), .A1 (nx537), .B0 (
                          bit_select_0), .C0 (nx543)) ;
    AOI22_X0P5M_A12TS ix532 (.Y (nx531), .A0 (ram_data_0), .A1 (nx533), .B0 (
                      ram_data_2), .B1 (nx535)) ;
    NOR2_X0P5A_A12TS ix534 (.Y (nx533), .A (bit_select_1), .B (bit_select_2)) ;
    AOI22_X0P5M_A12TS ix538 (.Y (nx537), .A0 (ram_data_4), .A1 (nx539), .B0 (
                      ram_data_6), .B1 (nx541)) ;
    AO1B2_X0P5M_A12TS ix544 (.Y (nx543), .A0N (bit_select_0), .B0 (nx545), .B1 (
                      nx547)) ;
    AOI22_X0P5M_A12TS ix546 (.Y (nx545), .A0 (ram_data_1), .A1 (nx533), .B0 (
                      ram_data_3), .B1 (nx535)) ;
    AOI22_X0P5M_A12TS ix548 (.Y (nx547), .A0 (ram_data_5), .A1 (nx539), .B0 (
                      ram_data_7), .B1 (nx541)) ;
    INV_X0P5B_A12TS ix303 (.Y (nx302), .A (nx533)) ;
    INV_X0P5B_A12TS ix1030 (.Y (nx1058), .A (nx535)) ;
    INV_X0P5B_A12TS ix227 (.Y (nx226), .A (nx539)) ;
    INV_X0P5B_A12TS ix542 (.Y (nx541), .A (nx1057)) ;
    INV_X0P5B_A12TS ix155 (.Y (nx154), .A (NOT_rd_en)) ;
    INV_X0P5B_A12TS ix21 (.Y (nx20), .A (nx351)) ;
    INV_X2M_A12TS ix117 (.Y (rd_addr_m_4), .A (nx397)) ;
    INV_X0P5B_A12TS ix139 (.Y (rd_addr_m_6), .A (nx409)) ;
    INV_X11M_A12TS ix71 (.Y (rd_addr_m_0), .A (nx375)) ;
    INV_X13M_A12TS ix1031 (.Y (rd_addr_m_1), .A (nx367)) ;
    INV_X4M_A12TS ix31 (.Y (rd_addr_m_2), .A (nx383)) ;
    INV_X4M_A12TS ix97 (.Y (rd_addr_m_3), .A (nx391)) ;
    INV_X1M_A12TS ix1032 (.Y (rd_addr_m_5), .A (nx403)) ;
    NOR2B_X0P7M_A12TS ix1034 (.Y (wr_addr_m_4), .AN (wr_addr_4), .B (nx339)) ;
    NOR2B_X0P7M_A12TS ix141 (.Y (wr_addr_m_6), .AN (wr_addr_6), .B (nx339)) ;
    XNOR2_X0P5M_A12TS ix366 (.Y (nx365), .A (nx367), .B (nx371)) ;
    XNOR2_X0P5M_A12TS ix374 (.Y (nx373), .A (nx375), .B (nx379)) ;
    XOR2_X0P5M_A12TS ix1035 (.Y (nx88), .A (nx383), .B (nx387)) ;
    NOR2B_X0P7M_A12TS ix536 (.Y (nx535), .AN (bit_select_1), .B (bit_select_2)
                      ) ;
    NOR2B_X0P7M_A12TS ix540 (.Y (nx539), .AN (bit_select_2), .B (bit_select_1)
                      ) ;
    MXT2_X0P5M_A12TS ix453 (.Y (src3_0), .A (dptr_hi_0), .B (pc_8), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix1064 (.Y (src3_1), .A (dptr_hi_1), .B (pc_9), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix469 (.Y (src3_2), .A (dptr_hi_2), .B (pc_10), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix477 (.Y (src3_3), .A (dptr_hi_3), .B (pc_11), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix1065 (.Y (src3_4), .A (dptr_hi_4), .B (pc_12), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix1066 (.Y (src3_5), .A (dptr_hi_5), .B (pc_13), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix501 (.Y (src3_6), .A (dptr_hi_6), .B (pc_14), .S0 (
                     src_sel3)) ;
    MXT2_X0P5M_A12TS ix1068 (.Y (src3_7), .A (dptr_hi_7), .B (pc_15), .S0 (
                     src_sel3)) ;
    AO1B2_X0P5M_A12TS ix1070 (.Y (src2_0), .A0N (nx526), .B0 (ram_out_0), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix527 (.Y (nx526), .A0 (acc_0), .A1 (nx1145), .B0 (op2_r_0
                      ), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_0 (.Q (op2_r_0), .CK (wb_clk_i), .D (op2_n_0), 
                       .R (wb_rst_i)) ;
    AND2_X0P5M_A12TS ix1071 (.Y (nx1146), .A (src_sel2_0), .B (src_sel2_1)) ;
    NOR2_X0P5A_A12TS ix1072 (.Y (nx1144), .A (src_sel2_0), .B (src_sel2_1)) ;
    AO1B2_X0P5M_A12TS ix39 (.Y (src2_1), .A0N (nx1153), .B0 (ram_out_1), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix1073 (.Y (nx1153), .A0 (acc_1), .A1 (nx1145), .B0 (
                      op2_r_1), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_1 (.Q (op2_r_1), .CK (wb_clk_i), .D (op2_n_1), 
                       .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix53 (.Y (src2_2), .A0N (nx1154), .B0 (ram_out_2), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix1074 (.Y (nx1154), .A0 (acc_2), .A1 (nx1145), .B0 (
                      op2_r_2), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_2 (.Q (op2_r_2), .CK (wb_clk_i), .D (op2_n_2), 
                       .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix67 (.Y (src2_3), .A0N (nx1155), .B0 (ram_out_3), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix1075 (.Y (nx1155), .A0 (acc_3), .A1 (nx1145), .B0 (
                      op2_r_3), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_3 (.Q (op2_r_3), .CK (wb_clk_i), .D (op2_n_3), 
                       .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix1076 (.Y (src2_4), .A0N (nx1156), .B0 (ram_out_4), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix1078 (.Y (nx1156), .A0 (acc_4), .A1 (nx1145), .B0 (
                      op2_r_4), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_4 (.Q (op2_r_4), .CK (wb_clk_i), .D (op2_n_4), 
                       .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix1079 (.Y (src2_5), .A0N (nx551), .B0 (ram_out_5), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix552 (.Y (nx551), .A0 (acc_5), .A1 (nx1145), .B0 (op2_r_5
                      ), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_5 (.Q (op2_r_5), .CK (wb_clk_i), .D (op2_n_5), 
                       .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix109 (.Y (src2_6), .A0N (nx555), .B0 (ram_out_6), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix556 (.Y (nx555), .A0 (acc_6), .A1 (nx1145), .B0 (op2_r_6
                      ), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_6 (.Q (op2_r_6), .CK (wb_clk_i), .D (op2_n_6), 
                       .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix123 (.Y (src2_7), .A0N (nx559), .B0 (ram_out_7), .B1 (
                      nx1144)) ;
    AOI22_X0P5M_A12TS ix560 (.Y (nx559), .A0 (acc_7), .A1 (nx1145), .B0 (op2_r_7
                      ), .B1 (nx1146)) ;
    DFFRPQ_X0P5M_A12TS reg_op2_r_7 (.Q (op2_r_7), .CK (wb_clk_i), .D (op2_n_7), 
                       .R (wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix1080 (.Y (src1_0), .A (nx563), .B (nx572), .C (nx578)) ;
    AOI222_X0P5M_A12TS ix564 (.Y (nx563), .A0 (ram_out_0), .A1 (nx1150), .B0 (
                       op2_r_0), .B1 (nx1151), .C0 (pc_8), .C1 (nx176)) ;
    NOR3_X0P5A_A12TS ix1082 (.Y (nx1150), .A (src_sel1_0), .B (src_sel1_2), .C (
                     src_sel1_1)) ;
    NOR3_X0P5A_A12TS ix1083 (.Y (nx1151), .A (nx567), .B (src_sel1_2), .C (
                     src_sel1_1)) ;
    INV_X0P5B_A12TS ix568 (.Y (nx567), .A (src_sel1_0)) ;
    NOR3_X0P5A_A12TS ix177 (.Y (nx176), .A (src_sel1_0), .B (nx1157), .C (
                     src_sel1_1)) ;
    INV_X0P5B_A12TS ix1084 (.Y (nx1157), .A (src_sel1_2)) ;
    AOI22_X0P5M_A12TS ix573 (.Y (nx572), .A0 (acc_0), .A1 (nx1149), .B0 (pc_0), 
                      .B1 (nx1148)) ;
    NOR3_X0P5A_A12TS ix1086 (.Y (nx1149), .A (nx567), .B (src_sel1_2), .C (nx575
                     )) ;
    INV_X0P5B_A12TS ix576 (.Y (nx575), .A (src_sel1_1)) ;
    NOR3_X0P5A_A12TS ix1087 (.Y (nx1148), .A (nx567), .B (nx1157), .C (
                     src_sel1_1)) ;
    AOI22_X0P5M_A12TS ix579 (.Y (nx578), .A0 (op1_r_0), .A1 (nx1147), .B0 (
                      op3_r_0), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_0 (.Q (op1_r_0), .CK (wb_clk_i), .D (op1_n_0), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_0 (.Q (op3_r_0), .CK (wb_clk_i), .D (op3_n_0), 
                       .R (wb_rst_i)) ;
    NOR3_X0P5A_A12TS ix135 (.Y (nx134), .A (src_sel1_0), .B (src_sel1_2), .C (
                     nx575)) ;
    NAND3_X1M_A12TS ix1088 (.Y (src1_1), .A (nx585), .B (nx587), .C (nx589)) ;
    AOI222_X0P5M_A12TS ix586 (.Y (nx585), .A0 (ram_out_1), .A1 (nx1150), .B0 (
                       op2_r_1), .B1 (nx1151), .C0 (pc_9), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix588 (.Y (nx587), .A0 (acc_1), .A1 (nx1149), .B0 (pc_1), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix590 (.Y (nx589), .A0 (op1_r_1), .A1 (nx1147), .B0 (
                      op3_r_1), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_1 (.Q (op1_r_1), .CK (wb_clk_i), .D (op1_n_1), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_1 (.Q (op3_r_1), .CK (wb_clk_i), .D (op3_n_1), 
                       .R (wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix1089 (.Y (src1_2), .A (nx594), .B (nx596), .C (nx598)) ;
    AOI222_X0P5M_A12TS ix595 (.Y (nx594), .A0 (ram_out_2), .A1 (nx1150), .B0 (
                       op2_r_2), .B1 (nx1151), .C0 (pc_10), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix597 (.Y (nx596), .A0 (acc_2), .A1 (nx1149), .B0 (pc_2), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix599 (.Y (nx598), .A0 (op1_r_2), .A1 (nx1147), .B0 (
                      op3_r_2), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_2 (.Q (op1_r_2), .CK (wb_clk_i), .D (op1_n_2), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_2 (.Q (op3_r_2), .CK (wb_clk_i), .D (op3_n_2), 
                       .R (wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix1090 (.Y (src1_3), .A (nx603), .B (nx605), .C (nx607)) ;
    AOI222_X0P5M_A12TS ix604 (.Y (nx603), .A0 (ram_out_3), .A1 (nx1150), .B0 (
                       op2_r_3), .B1 (nx1151), .C0 (pc_11), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix606 (.Y (nx605), .A0 (acc_3), .A1 (nx1149), .B0 (pc_3), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix608 (.Y (nx607), .A0 (op1_r_3), .A1 (nx1147), .B0 (
                      op3_r_3), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_3 (.Q (op1_r_3), .CK (wb_clk_i), .D (op1_n_3), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_3 (.Q (op3_r_3), .CK (wb_clk_i), .D (op3_n_3), 
                       .R (wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix1091 (.Y (src1_4), .A (nx612), .B (nx614), .C (nx616)) ;
    AOI222_X0P5M_A12TS ix613 (.Y (nx612), .A0 (ram_out_4), .A1 (nx1150), .B0 (
                       op2_r_4), .B1 (nx1151), .C0 (pc_12), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix615 (.Y (nx614), .A0 (acc_4), .A1 (nx1149), .B0 (pc_4), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix617 (.Y (nx616), .A0 (op1_r_4), .A1 (nx1147), .B0 (
                      op3_r_4), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_4 (.Q (op1_r_4), .CK (wb_clk_i), .D (op1_n_4), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_4 (.Q (op3_r_4), .CK (wb_clk_i), .D (op3_n_4), 
                       .R (wb_rst_i)) ;
    NAND3_X1M_A12TS ix1092 (.Y (src1_5), .A (nx621), .B (nx623), .C (nx625)) ;
    AOI222_X0P5M_A12TS ix622 (.Y (nx621), .A0 (ram_out_5), .A1 (nx1150), .B0 (
                       op2_r_5), .B1 (nx1151), .C0 (pc_13), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix624 (.Y (nx623), .A0 (acc_5), .A1 (nx1149), .B0 (pc_5), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix626 (.Y (nx625), .A0 (op1_r_5), .A1 (nx1147), .B0 (
                      op3_r_5), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_5 (.Q (op1_r_5), .CK (wb_clk_i), .D (op1_n_5), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_5 (.Q (op3_r_5), .CK (wb_clk_i), .D (op3_n_5), 
                       .R (wb_rst_i)) ;
    NAND3_X1M_A12TS ix1093 (.Y (src1_6), .A (nx630), .B (nx632), .C (nx634)) ;
    AOI222_X0P5M_A12TS ix631 (.Y (nx630), .A0 (ram_out_6), .A1 (nx1150), .B0 (
                       op2_r_6), .B1 (nx1151), .C0 (pc_14), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix633 (.Y (nx632), .A0 (acc_6), .A1 (nx1149), .B0 (pc_6), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix635 (.Y (nx634), .A0 (op1_r_6), .A1 (nx1147), .B0 (
                      op3_r_6), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_6 (.Q (op1_r_6), .CK (wb_clk_i), .D (op1_n_6), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_6 (.Q (op3_r_6), .CK (wb_clk_i), .D (op3_n_6), 
                       .R (wb_rst_i)) ;
    NAND3_X1M_A12TS ix445 (.Y (src1_7), .A (nx639), .B (nx641), .C (nx643)) ;
    AOI222_X0P5M_A12TS ix640 (.Y (nx639), .A0 (ram_out_7), .A1 (nx1150), .B0 (
                       op2_r_7), .B1 (nx1151), .C0 (pc_15), .C1 (nx176)) ;
    AOI22_X0P5M_A12TS ix642 (.Y (nx641), .A0 (acc_7), .A1 (nx1149), .B0 (pc_7), 
                      .B1 (nx1148)) ;
    AOI22_X0P5M_A12TS ix644 (.Y (nx643), .A0 (op1_r_7), .A1 (nx1147), .B0 (
                      op3_r_7), .B1 (nx134)) ;
    DFFRPQ_X0P5M_A12TS reg_op1_r_7 (.Q (op1_r_7), .CK (wb_clk_i), .D (op1_n_7), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_op3_r_7 (.Q (op3_r_7), .CK (wb_clk_i), .D (op3_n_7), 
                       .R (wb_rst_i)) ;
    NOR2B_X0P7M_A12TS ix1094 (.Y (nx1145), .AN (src_sel2_0), .B (src_sel2_1)) ;
    AND3_X0P5M_A12TS ix1095 (.Y (nx1147), .A (src_sel1_0), .B (src_sel1_2), .C (
                     src_sel1_1)) ;
    AO21A1AI2_X0P5M_A12TS ix1158 (.Y (eq), .A0 (nx111), .A1 (nx119), .B0 (
                          comp_sel_1), .C0 (nx125)) ;
    NAND4_X0P5A_A12TS ix112 (.Y (nx111), .A (nx1177), .B (nx46), .C (nx54), .D (
                      nx1179)) ;
    NOR3_X0P5A_A12TS ix1159 (.Y (nx1177), .A (sub_result_6), .B (nx1180), .C (
                     sub_result_7)) ;
    INV_X0P5B_A12TS ix1160 (.Y (nx1180), .A (comp_sel_0)) ;
    NOR2_X0P5A_A12TS ix47 (.Y (nx46), .A (sub_result_5), .B (sub_result_4)) ;
    NOR2_X0P5A_A12TS ix55 (.Y (nx54), .A (sub_result_3), .B (sub_result_2)) ;
    NOR2_X0P5A_A12TS ix1162 (.Y (nx1179), .A (sub_result_1), .B (sub_result_0)
                     ) ;
    NAND4_X0P5A_A12TS ix120 (.Y (nx119), .A (nx8), .B (nx14), .C (nx1175), .D (
                      nx28)) ;
    NOR3_X0P5A_A12TS ix9 (.Y (nx8), .A (acc_6), .B (comp_sel_0), .C (acc_7)) ;
    NOR2_X0P5A_A12TS ix15 (.Y (nx14), .A (acc_5), .B (acc_4)) ;
    NOR2_X0P5A_A12TS ix1164 (.Y (nx1175), .A (acc_3), .B (acc_2)) ;
    NOR2_X0P5A_A12TS ix29 (.Y (nx28), .A (acc_1), .B (acc_0)) ;
    AO21A1AI2_X0P5M_A12TS ix126 (.Y (nx125), .A0 (bit_out), .A1 (comp_sel_0), .B0 (
                          nx74), .C0 (comp_sel_1)) ;
    NOR2B_X0P7M_A12TS ix78 (.Y (nx74), .AN (cy), .B (comp_sel_0)) ;
    AO21B_X2M_A12TS ix1181 (.Y (alu_cy), .B0N (nx43), .A0 (bit_out), .A1 (
                    cy_sel_1)) ;
    OAI21_X0P5M_A12TS ix44 (.Y (nx43), .A0 (cy_sel_1), .A1 (cy), .B0 (cy_sel_0)
                      ) ;
    NAND4_X0P5A_A12TS ix1184 (.Y (ri_0), .A (nx1992), .B (nx1241), .C (nx1244), 
                      .D (nx1245)) ;
    AOI22_X0P5M_A12TS ix1993 (.Y (nx1992), .A0 (des1_0), .A1 (nx1235), .B0 (
                      buff_4__0), .B1 (nx212)) ;
    INV_X0P5B_A12TS ix1186 (.Y (nx1235), .A (nx1995)) ;
    OR6_X0P5M_A12TS ix1996 (.Y (nx1995), .A (wr_addr_5), .B (wr_addr_7), .C (
                    wr_addr_6), .D (wr_addr_2), .E (wr_addr_1), .F (nx1238)) ;
    DFFRPQ_X0P5M_A12TS reg_wr_bit_r (.Q (wr_bit_r), .CK (wb_clk_i), .D (bit_addr
                       ), .R (wb_rst_i)) ;
    XNOR2_X0P5M_A12TS ix2002 (.Y (nx2001), .A (op1_cur_0), .B (wr_addr_0)) ;
    XNOR2_X0P5M_A12TS ix2004 (.Y (nx2003), .A (bank_sel_0), .B (wr_addr_3)) ;
    XNOR2_X0P5M_A12TS ix2006 (.Y (nx2005), .A (bank_sel_1), .B (wr_addr_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__0 (.Q (buff_4__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__0)
                        ) ;
    NAND3_X0P5A_A12TS ix2009 (.Y (NOT_nx202), .A (nx118), .B (nx2015), .C (
                      nx2017)) ;
    NAND2B_X0P7M_A12TS ix1187 (.Y (nx1239), .AN (wr_bit_r), .B (wr)) ;
    INV_X0P5B_A12TS ix2016 (.Y (nx2015), .A (wr_addr_0)) ;
    INV_X0P5B_A12TS ix2018 (.Y (nx2017), .A (wr_addr_3)) ;
    NOR3_X0P5A_A12TS ix213 (.Y (nx212), .A (nx2020), .B (nx2024), .C (op1_cur_0)
                     ) ;
    INV_X0P5B_A12TS ix2025 (.Y (nx2024), .A (bank_sel_1)) ;
    AOI22_X0P5M_A12TS ix1188 (.Y (nx1241), .A0 (buff_5__0), .A1 (nx190), .B0 (
                      buff_6__0), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__0 (.Q (buff_5__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__0)
                        ) ;
    NAND3_X0P5A_A12TS ix2030 (.Y (NOT_nx182), .A (nx118), .B (wr_addr_0), .C (
                      nx2017)) ;
    NOR3_X0P5A_A12TS ix191 (.Y (nx190), .A (nx2020), .B (nx2024), .C (nx2032)) ;
    INV_X0P5B_A12TS ix2033 (.Y (nx2032), .A (op1_cur_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__0 (.Q (buff_6__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__0)
                        ) ;
    NAND3_X0P5A_A12TS ix1190 (.Y (NOT_nx164), .A (nx118), .B (nx2015), .C (
                      wr_addr_3)) ;
    NOR3_X0P5A_A12TS ix1191 (.Y (nx1237), .A (nx1243), .B (nx2024), .C (
                     op1_cur_0)) ;
    NAND2_X0P5A_A12TS ix1192 (.Y (nx1243), .A (bank_sel_0), .B (nx1995)) ;
    AOI22_X0P5M_A12TS ix1193 (.Y (nx1244), .A0 (buff_0__0), .A1 (nx152), .B0 (
                      buff_7__0), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__0 (.Q (buff_0__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__0)
                        ) ;
    NAND3_X0P5A_A12TS ix1194 (.Y (NOT_nx140), .A (nx1234), .B (nx2015), .C (
                      nx2017)) ;
    NOR2_X0P5A_A12TS ix1195 (.Y (nx1234), .A (wr_addr_4), .B (nx1239)) ;
    NOR3_X0P5A_A12TS ix153 (.Y (nx152), .A (nx2020), .B (bank_sel_1), .C (
                     op1_cur_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__0 (.Q (buff_7__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__0)
                        ) ;
    NAND3_X0P5A_A12TS ix1196 (.Y (NOT_nx122), .A (nx118), .B (wr_addr_0), .C (
                      wr_addr_3)) ;
    NOR3_X0P5A_A12TS ix131 (.Y (nx130), .A (nx1243), .B (nx2024), .C (nx2032)) ;
    AOI222_X0P5M_A12TS ix1198 (.Y (nx1245), .A0 (buff_1__0), .A1 (nx1236), .B0 (
                       buff_2__0), .B1 (nx86), .C0 (buff_3__0), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__0 (.Q (buff_1__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__0)
                        ) ;
    NAND3_X0P5A_A12TS ix1199 (.Y (NOT_nx94), .A (nx1234), .B (wr_addr_0), .C (
                      nx2017)) ;
    NOR3_X0P5A_A12TS ix1200 (.Y (nx1236), .A (nx2020), .B (bank_sel_1), .C (
                     nx2032)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__0 (.Q (buff_2__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__0)
                        ) ;
    NAND3_X0P5A_A12TS ix2059 (.Y (NOT_nx74), .A (nx1234), .B (nx2015), .C (
                      wr_addr_3)) ;
    NOR3_X0P5A_A12TS ix87 (.Y (nx86), .A (nx1243), .B (bank_sel_1), .C (
                     op1_cur_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__0 (.Q (buff_3__0), .CK (wb_clk_i), .D (
                        des1_0), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__0)
                        ) ;
    NAND3_X0P5A_A12TS ix2063 (.Y (NOT_nx14), .A (nx1234), .B (wr_addr_0), .C (
                      wr_addr_3)) ;
    NOR3_X0P5A_A12TS ix1201 (.Y (nx66), .A (nx1243), .B (bank_sel_1), .C (nx2032
                     )) ;
    NAND4_X0P5A_A12TS ix1202 (.Y (ri_1), .A (nx1246), .B (nx2069), .C (nx2073), 
                      .D (nx1247)) ;
    AOI22_X0P5M_A12TS ix1203 (.Y (nx1246), .A0 (des1_1), .A1 (nx1235), .B0 (
                      buff_4__1), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__1 (.Q (buff_4__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__1)
                        ) ;
    AOI22_X0P5M_A12TS ix2070 (.Y (nx2069), .A0 (buff_5__1), .A1 (nx190), .B0 (
                      buff_6__1), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__1 (.Q (buff_5__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__1)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__1 (.Q (buff_6__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__1)
                        ) ;
    AOI22_X0P5M_A12TS ix2074 (.Y (nx2073), .A0 (buff_0__1), .A1 (nx152), .B0 (
                      buff_7__1), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__1 (.Q (buff_0__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__1)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__1 (.Q (buff_7__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__1)
                        ) ;
    AOI222_X0P5M_A12TS ix1204 (.Y (nx1247), .A0 (buff_1__1), .A1 (nx1236), .B0 (
                       buff_2__1), .B1 (nx86), .C0 (buff_3__1), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__1 (.Q (buff_1__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__1)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__1 (.Q (buff_2__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__1)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__1 (.Q (buff_3__1), .CK (wb_clk_i), .D (
                        des1_1), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__1)
                        ) ;
    NAND4_X0P5A_A12TS ix355 (.Y (ri_2), .A (nx1248), .B (nx1249), .C (nx2090), .D (
                      nx2094)) ;
    AOI22_X0P5M_A12TS ix1205 (.Y (nx1248), .A0 (des1_2), .A1 (nx1235), .B0 (
                      buff_4__2), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__2 (.Q (buff_4__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__2)
                        ) ;
    AOI22_X0P5M_A12TS ix1206 (.Y (nx1249), .A0 (buff_5__2), .A1 (nx190), .B0 (
                      buff_6__2), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__2 (.Q (buff_5__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__2)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__2 (.Q (buff_6__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__2)
                        ) ;
    AOI22_X0P5M_A12TS ix2091 (.Y (nx2090), .A0 (buff_0__2), .A1 (nx152), .B0 (
                      buff_7__2), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__2 (.Q (buff_0__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__2)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__2 (.Q (buff_7__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__2)
                        ) ;
    AOI222_X0P5M_A12TS ix2095 (.Y (nx2094), .A0 (buff_1__2), .A1 (nx1236), .B0 (
                       buff_2__2), .B1 (nx86), .C0 (buff_3__2), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__2 (.Q (buff_1__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__2)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__2 (.Q (buff_2__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__2)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__2 (.Q (buff_3__2), .CK (wb_clk_i), .D (
                        des1_2), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__2)
                        ) ;
    NAND4_X0P5A_A12TS ix1207 (.Y (ri_3), .A (nx2100), .B (nx1250), .C (nx2107), 
                      .D (nx1251)) ;
    AOI22_X0P5M_A12TS ix2101 (.Y (nx2100), .A0 (des1_3), .A1 (nx1235), .B0 (
                      buff_4__3), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__3 (.Q (buff_4__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__3)
                        ) ;
    AOI22_X0P5M_A12TS ix1208 (.Y (nx1250), .A0 (buff_5__3), .A1 (nx190), .B0 (
                      buff_6__3), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__3 (.Q (buff_5__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__3)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__3 (.Q (buff_6__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__3)
                        ) ;
    AOI22_X0P5M_A12TS ix2108 (.Y (nx2107), .A0 (buff_0__3), .A1 (nx152), .B0 (
                      buff_7__3), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__3 (.Q (buff_0__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__3)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__3 (.Q (buff_7__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__3)
                        ) ;
    AOI222_X0P5M_A12TS ix1210 (.Y (nx1251), .A0 (buff_1__3), .A1 (nx1236), .B0 (
                       buff_2__3), .B1 (nx86), .C0 (buff_3__3), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__3 (.Q (buff_1__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__3)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__3 (.Q (buff_2__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__3)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__3 (.Q (buff_3__3), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__3)
                        ) ;
    NAND4_X0P5A_A12TS ix1211 (.Y (ri_4), .A (nx2117), .B (nx1253), .C (nx2124), 
                      .D (nx2128)) ;
    AOI22_X0P5M_A12TS ix2118 (.Y (nx2117), .A0 (des1_4), .A1 (nx1235), .B0 (
                      buff_4__4), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__4 (.Q (buff_4__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__4)
                        ) ;
    AOI22_X0P5M_A12TS ix1212 (.Y (nx1253), .A0 (buff_5__4), .A1 (nx190), .B0 (
                      buff_6__4), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__4 (.Q (buff_5__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__4)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__4 (.Q (buff_6__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__4)
                        ) ;
    AOI22_X0P5M_A12TS ix2125 (.Y (nx2124), .A0 (buff_0__4), .A1 (nx152), .B0 (
                      buff_7__4), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__4 (.Q (buff_0__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__4)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__4 (.Q (buff_7__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__4)
                        ) ;
    AOI222_X0P5M_A12TS ix2129 (.Y (nx2128), .A0 (buff_1__4), .A1 (nx1236), .B0 (
                       buff_2__4), .B1 (nx86), .C0 (buff_3__4), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__4 (.Q (buff_1__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__4)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__4 (.Q (buff_2__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__4)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__4 (.Q (buff_3__4), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__4)
                        ) ;
    NAND4_X0P5A_A12TS ix553 (.Y (ri_5), .A (nx2134), .B (nx1255), .C (nx2141), .D (
                      nx2145)) ;
    AOI22_X0P5M_A12TS ix2135 (.Y (nx2134), .A0 (des1_5), .A1 (nx1235), .B0 (
                      buff_4__5), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__5 (.Q (buff_4__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__5)
                        ) ;
    AOI22_X0P5M_A12TS ix1214 (.Y (nx1255), .A0 (buff_5__5), .A1 (nx190), .B0 (
                      buff_6__5), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__5 (.Q (buff_5__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__5)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__5 (.Q (buff_6__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__5)
                        ) ;
    AOI22_X0P5M_A12TS ix2142 (.Y (nx2141), .A0 (buff_0__5), .A1 (nx152), .B0 (
                      buff_7__5), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__5 (.Q (buff_0__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__5)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__5 (.Q (buff_7__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__5)
                        ) ;
    AOI222_X0P5M_A12TS ix2146 (.Y (nx2145), .A0 (buff_1__5), .A1 (nx1236), .B0 (
                       buff_2__5), .B1 (nx86), .C0 (buff_3__5), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__5 (.Q (buff_1__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__5)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__5 (.Q (buff_2__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__5)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__5 (.Q (buff_3__5), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__5)
                        ) ;
    NAND4_X0P5A_A12TS ix619 (.Y (ri_6), .A (nx1257), .B (nx1259), .C (nx2158), .D (
                      nx1260)) ;
    AOI22_X0P5M_A12TS ix1216 (.Y (nx1257), .A0 (des1_6), .A1 (nx1235), .B0 (
                      buff_4__6), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__6 (.Q (buff_4__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__6)
                        ) ;
    AOI22_X0P5M_A12TS ix1217 (.Y (nx1259), .A0 (buff_5__6), .A1 (nx190), .B0 (
                      buff_6__6), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__6 (.Q (buff_5__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__6)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__6 (.Q (buff_6__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__6)
                        ) ;
    AOI22_X0P5M_A12TS ix2159 (.Y (nx2158), .A0 (buff_0__6), .A1 (nx152), .B0 (
                      buff_7__6), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__6 (.Q (buff_0__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__6)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__6 (.Q (buff_7__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__6)
                        ) ;
    AOI222_X0P5M_A12TS ix1218 (.Y (nx1260), .A0 (buff_1__6), .A1 (nx1236), .B0 (
                       buff_2__6), .B1 (nx86), .C0 (buff_3__6), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__6 (.Q (buff_1__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__6)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__6 (.Q (buff_2__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__6)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__6 (.Q (buff_3__6), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__6)
                        ) ;
    NAND4_X0P5A_A12TS ix1219 (.Y (ri_7), .A (nx1261), .B (nx2171), .C (nx2175), 
                      .D (nx1262)) ;
    AOI22_X0P5M_A12TS ix1220 (.Y (nx1261), .A0 (des1_7), .A1 (nx1235), .B0 (
                      buff_4__7), .B1 (nx212)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_4__7 (.Q (buff_4__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx202), .SI (buff_4__7)
                        ) ;
    AOI22_X0P5M_A12TS ix2172 (.Y (nx2171), .A0 (buff_5__7), .A1 (nx190), .B0 (
                      buff_6__7), .B1 (nx1237)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_5__7 (.Q (buff_5__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx182), .SI (buff_5__7)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_6__7 (.Q (buff_6__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx164), .SI (buff_6__7)
                        ) ;
    AOI22_X0P5M_A12TS ix2176 (.Y (nx2175), .A0 (buff_0__7), .A1 (nx152), .B0 (
                      buff_7__7), .B1 (nx130)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_0__7 (.Q (buff_0__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx140), .SI (buff_0__7)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_7__7 (.Q (buff_7__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx122), .SI (buff_7__7)
                        ) ;
    AOI222_X0P5M_A12TS ix1222 (.Y (nx1262), .A0 (buff_1__7), .A1 (nx1236), .B0 (
                       buff_2__7), .B1 (nx86), .C0 (buff_3__7), .C1 (nx66)) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_1__7 (.Q (buff_1__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx94), .SI (buff_1__7)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_2__7 (.Q (buff_2__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx74), .SI (buff_2__7)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_buff_3__7 (.Q (buff_3__7), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx14), .SI (buff_3__7)
                        ) ;
    NAND4B_X0P5M_A12TS ix1223 (.Y (nx1238), .AN (nx1239), .B (nx2001), .C (
                       nx2003), .D (nx2005)) ;
    NOR2B_X0P7M_A12TS ix1224 (.Y (nx118), .AN (wr_addr_4), .B (nx1239)) ;
    NAND2B_X0P7M_A12TS ix2021 (.Y (nx2020), .AN (bank_sel_0), .B (nx1995)) ;
    NOR2_X0P5A_A12TS ix1613 (.Y (wr_ind), .A (ram_wr_sel_2), .B (nx7505)) ;
    INV_X0P5B_A12TS ix7506 (.Y (nx7505), .A (ram_wr_sel_1)) ;
    DFFRPQ_X0P5M_A12TS reg_dmem_wait (.Q (wbd_stb_o), .CK (wb_clk_i), .D (
                       NOT_dack_i), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix7509 (.Y (NOT_dack_i), .A (wbd_ack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_reti (.Q (reti), .CK (wb_clk_i), .D (nx3968), .R (
                       wb_rst_i)) ;
    NOR3_X0P5A_A12TS ix3969 (.Y (nx3968), .A (nx7512), .B (nx8106), .C (nx8108)
                     ) ;
    NAND3_X0P5A_A12TS ix7513 (.Y (nx7512), .A (nx1478), .B (rd), .C (nx7867)) ;
    OAI211_X0P5M_A12TS ix1263 (.Y (nx1478), .A0 (nx7515), .A1 (nx7778), .B0 (
                       nx7780), .C0 (nx8083)) ;
    MXIT2_X0P5M_A12TS ix7516 (.Y (nx7515), .A (idat_cur_1), .B (idat_cur_9), .S0 (
                      op_pos_0)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_1 (.Q (idat_cur_1), .CK (wb_clk_i), .D (
                       nx5914), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5915 (.Y (nx5914), .A0 (nx7519), .A1 (NOT_nx5673), .B0 (
                      nx8075)) ;
    AOI32_X0P5M_A12TS ix7520 (.Y (nx7519), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[1]), .B1 (nx7521)) ;
    NAND2_X1M_A12TS ix7522 (.Y (nx7521), .A (ea_int), .B (ea_in)) ;
    OAI21_X3M_A12TS ix7524 (.Y (NOT_nx5673), .A0 (nx5672), .A1 (pc_wr_r2), .B0 (
                    nx26)) ;
    NAND2_X0P5A_A12TS ix1375 (.Y (nx5672), .A (nx7526), .B (nx7603)) ;
    AO21A1AI2_X0P5M_A12TS ix7527 (.Y (nx7526), .A0 (op_pos_1), .A1 (op_pos_0), .B0 (
                          op_pos_2), .C0 (rd)) ;
    DFFRPQ_X0P5M_A12TS reg_op_pos_1 (.Q (op_pos_1), .CK (wb_clk_i), .D (nx6424)
                       , .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix6425 (.Y (nx6424), .A0 (pc_wr_r2), .A1 (nx7539), .A2 (
                      NOT_rd), .B0 (nx8073)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_wr_r2 (.Q (pc_wr_r2), .CK (wb_clk_i), .D (pc_wr_r)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_wr_r (.Q (pc_wr_r), .CK (wb_clk_i), .D (nx36), .R (
                       wb_rst_i)) ;
    INV_X0P5B_A12TS ix7534 (.Y (nx7533), .A (pc_wr_sel_2)) ;
    INV_X0P5B_A12TS ix7538 (.Y (nx7537), .A (pc_wr_dup_1371)) ;
    XNOR2_X0P5M_A12TS ix7540 (.Y (nx7539), .A (nx7541), .B (nx8071)) ;
    NAND2_X0P5A_A12TS ix7542 (.Y (nx7541), .A (op_pos_0), .B (nx5677)) ;
    DFFRPQ_X0P5M_A12TS reg_op_pos_0 (.Q (op_pos_0), .CK (wb_clk_i), .D (nx6504)
                       , .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix6505 (.Y (nx6504), .A (nx7545), .B (nx7591), .S0 (nx8069
                      )) ;
    OAI211_X0P5M_A12TS ix7546 (.Y (nx7545), .A0 (nx5677), .A1 (op_pos_0), .B0 (
                       nx7603), .C0 (nx7541)) ;
    OAI211_X0P5M_A12TS ix1323 (.Y (nx5677), .A0 (op1_n_7), .A1 (nx8035), .B0 (
                       nx8056), .C0 (nx8037)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_7 (.Q (cdata_7), .CK (wb_clk_i), .D (nx6494), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6495 (.Y (nx6494), .A0 (nx7553), .A1 (nx7555), .B0 (
                      nx7570)) ;
    AOI32_X0P5M_A12TS ix7554 (.Y (nx7553), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[7]), .B1 (nx7521)) ;
    INV_X0P5B_A12TS ix7556 (.Y (nx7555), .A (istb_t)) ;
    DFFRPQ_X0P5M_A12TS reg_istb_t (.Q (istb_t), .CK (wb_clk_i), .D (nx5824), .R (
                       wb_rst_i)) ;
    INV_X0P5B_A12TS ix7560 (.Y (nx7559), .A (imem_wait)) ;
    DFFRPQ_X0P5M_A12TS reg_imem_wait (.Q (imem_wait), .CK (wb_clk_i), .D (nx5814
                       ), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix5815 (.Y (nx5814), .A0 (nx7559), .A1 (nx1469), .A2 (
                      wbi_ack_i), .B0 (NOT_nx226)) ;
    NAND3_X0P5A_A12TS ix7565 (.Y (NOT_nx226), .A (nx7566), .B (mem_act_2), .C (
                      nx7568)) ;
    INV_X0P5B_A12TS ix7567 (.Y (nx7566), .A (mem_act_1)) ;
    INV_X0P5B_A12TS ix7569 (.Y (nx7568), .A (mem_act_0)) ;
    NAND2_X0P5A_A12TS ix7571 (.Y (nx7570), .A (cdata_7), .B (nx7555)) ;
    NAND2_X0P5A_A12TS ix7573 (.Y (nx7572), .A (cdone), .B (nx7575)) ;
    DFFRPQ_X0P5M_A12TS reg_cdone (.Q (cdone), .CK (wb_clk_i), .D (istb_t), .R (
                       wb_rst_i)) ;
    INV_X0P5B_A12TS ix7576 (.Y (nx7575), .A (dack_ir)) ;
    DFFRPQ_X0P5M_A12TS reg_dack_ir (.Q (dack_ir), .CK (wb_clk_i), .D (wbd_ack_i)
                       , .R (wb_rst_i)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_7 (.Q (ddat_ir_7), .CK (wb_clk_i), .D (
                        wbd_dat_i[7]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_7)) ;
    AOI211_X0P5M_A12TS ix7582 (.Y (nx7581), .A0 (idat_old_15), .A1 (nx5675), .B0 (
                       nx1166), .C0 (nx1114)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_15 (.Q (idat_old_15), .CK (wb_clk_i), .D (
                        idat_cur_15), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_15)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_15 (.Q (idat_cur_15), .CK (wb_clk_i), .D (
                       nx5694), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5695 (.Y (nx5694), .A0 (nx7586), .A1 (NOT_nx5673), .B0 (
                      nx7588)) ;
    AOI32_X0P5M_A12TS ix7587 (.Y (nx7586), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[15]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7589 (.Y (nx7588), .A (idat_cur_15), .B (NOT_nx5673)) ;
    NOR2_X0P5A_A12TS ix1264 (.Y (nx5675), .A (nx7591), .B (nx7593)) ;
    INV_X0P5B_A12TS ix7592 (.Y (nx7591), .A (op_pos_0)) ;
    NAND2_X0P5A_A12TS ix7594 (.Y (nx7593), .A (nx7595), .B (nx164)) ;
    INV_X0P5B_A12TS ix7596 (.Y (nx7595), .A (op_pos_1)) ;
    NOR2_X0P5A_A12TS ix165 (.Y (nx164), .A (op_pos_2), .B (nx1473)) ;
    DFFRPQ_X0P5M_A12TS reg_op_pos_2 (.Q (op_pos_2), .CK (wb_clk_i), .D (nx6514)
                       , .R (wb_rst_i)) ;
    OAI221_X0P5M_A12TS ix6515 (.Y (nx6514), .A0 (nx7600), .A1 (nx1470), .B0 (
                       nx7607), .B1 (NOT_rd), .C0 (nx7603)) ;
    INV_X0P5B_A12TS ix7601 (.Y (nx7600), .A (op_pos_2)) ;
    INV_X0P5B_A12TS ix7604 (.Y (nx7603), .A (pc_wr_r2)) ;
    INV_X0P5B_A12TS ix7606 (.Y (NOT_rd), .A (rd)) ;
    AOI32_X0P5M_A12TS ix7608 (.Y (nx7607), .A0 (nx1340), .A1 (nx1070), .A2 (
                      nx392), .B0 (nx1354), .B1 (nx7610)) ;
    NOR2_X0P5A_A12TS ix1266 (.Y (nx1340), .A (nx7541), .B (nx7610)) ;
    NAND2_X0P5A_A12TS ix7611 (.Y (nx7610), .A (rd), .B (nx5672)) ;
    AOI211_X0P5M_A12TS ix7614 (.Y (nx7613), .A0 (nx416), .A1 (nx1492), .B0 (
                       nx7905), .C0 (nx1042)) ;
    NOR2_X0P5A_A12TS ix417 (.Y (nx416), .A (op1_n_3), .B (op1_n_1)) ;
    OAI222_X0P5M_A12TS ix1268 (.Y (op1_n_3), .A0 (nx7617), .A1 (nx7572), .B0 (
                       nx7625), .B1 (nx7575), .C0 (nx7628), .C1 (nx7687)) ;
    INV_X0P5B_A12TS ix7618 (.Y (nx7617), .A (cdata_3)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_3 (.Q (cdata_3), .CK (wb_clk_i), .D (nx5834), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5835 (.Y (nx5834), .A0 (nx7621), .A1 (nx7555), .B0 (
                      nx7623)) ;
    AOI32_X0P5M_A12TS ix7622 (.Y (nx7621), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[3]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7624 (.Y (nx7623), .A (cdata_3), .B (nx7555)) ;
    INV_X0P5B_A12TS ix7626 (.Y (nx7625), .A (ddat_ir_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_3 (.Q (ddat_ir_3), .CK (wb_clk_i), .D (
                        wbd_dat_i[3]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_3)) ;
    AOI211_X0P5M_A12TS ix7629 (.Y (nx7628), .A0 (idat_old_11), .A1 (nx5675), .B0 (
                       nx1477), .C0 (nx1474)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_11 (.Q (idat_old_11), .CK (wb_clk_i), .D (
                        idat_cur_11), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_11)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_11 (.Q (idat_cur_11), .CK (wb_clk_i), .D (
                       nx5724), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5725 (.Y (nx5724), .A0 (nx7633), .A1 (NOT_nx5673), .B0 (
                      nx7635)) ;
    AOI32_X0P5M_A12TS ix7634 (.Y (nx7633), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[11]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7636 (.Y (nx7635), .A (idat_cur_11), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix1269 (.Y (nx1477), .A0 (nx7638), .A1 (nx7654), .B0 (
                      nx7656), .B1 (nx7663)) ;
    MXIT2_X0P5M_A12TS ix7639 (.Y (nx7638), .A (idat_old_19), .B (idat_old_27), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_19 (.Q (idat_old_19), .CK (wb_clk_i), .D (
                        idat_cur_19), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_19)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_19 (.Q (idat_cur_19), .CK (wb_clk_i), .D (
                       nx5774), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5775 (.Y (nx5774), .A0 (nx7643), .A1 (NOT_nx5673), .B0 (
                      nx7645)) ;
    AOI32_X0P5M_A12TS ix7644 (.Y (nx7643), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[19]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7646 (.Y (nx7645), .A (idat_cur_19), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_27 (.Q (idat_old_27), .CK (wb_clk_i), .D (
                        idat_cur_27), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_27)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_27 (.Q (idat_cur_27), .CK (wb_clk_i), .D (
                       nx5794), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5795 (.Y (nx5794), .A0 (nx7650), .A1 (NOT_nx5673), .B0 (
                      nx7652)) ;
    AOI32_X0P5M_A12TS ix7651 (.Y (nx7650), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[27]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7653 (.Y (nx7652), .A (idat_cur_27), .B (NOT_nx5673)) ;
    NAND2_X0P5A_A12TS ix7655 (.Y (nx7654), .A (op_pos_1), .B (nx164)) ;
    INV_X0P5B_A12TS ix7657 (.Y (nx7656), .A (idat_old_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_3 (.Q (idat_old_3), .CK (wb_clk_i), .D (
                        idat_cur_3), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_3)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_3 (.Q (idat_cur_3), .CK (wb_clk_i), .D (
                       nx5744), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5745 (.Y (nx5744), .A0 (nx7621), .A1 (NOT_nx5673), .B0 (
                      nx7661)) ;
    NAND2_X0P5A_A12TS ix7662 (.Y (nx7661), .A (idat_cur_3), .B (NOT_nx5673)) ;
    NAND2_X0P5A_A12TS ix7664 (.Y (nx7663), .A (nx7665), .B (nx164)) ;
    NOR2_X0P5A_A12TS ix7666 (.Y (nx7665), .A (op_pos_0), .B (op_pos_1)) ;
    OAI22_X0P5M_A12TS ix1270 (.Y (nx1474), .A0 (nx7668), .A1 (nx7670), .B0 (
                      nx7683), .B1 (nx7685)) ;
    INV_X0P5B_A12TS ix7669 (.Y (nx7668), .A (idat_cur_11)) ;
    NAND2_X0P5A_A12TS ix7671 (.Y (nx7670), .A (op_pos_1), .B (nx138)) ;
    NOR2_X0P5A_A12TS ix1272 (.Y (nx138), .A (nx7600), .B (nx1473)) ;
    NOR2_X0P5A_A12TS ix1274 (.Y (nx1473), .A (nx7674), .B (nx7679)) ;
    INV_X0P5B_A12TS ix7675 (.Y (nx7674), .A (int_ack_t)) ;
    DFFRPQ_X0P5M_A12TS reg_int_ack_t (.Q (int_ack_t), .CK (wb_clk_i), .D (nx5754
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5755 (.Y (nx5754), .A0 (nx7674), .A1 (nx1471), .B0 (
                      NOT_intr)) ;
    OAI31_X0P5M_A12TS ix1275 (.Y (nx1471), .A0 (nx7679), .A1 (NOT_rd), .A2 (
                      pc_wr_r2), .B0 (NOT_intr)) ;
    NOR2_X0P5A_A12TS ix7680 (.Y (nx7679), .A (nx1469), .B (wbi_ack_i)) ;
    INV_X0P5B_A12TS ix7682 (.Y (NOT_intr), .A (intr)) ;
    MXIT2_X0P5M_A12TS ix7684 (.Y (nx7683), .A (idat_cur_3), .B (idat_cur_11), .S0 (
                      op_pos_0)) ;
    NAND2_X0P5A_A12TS ix7686 (.Y (nx7685), .A (nx7595), .B (nx138)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_1 (.Q (ddat_ir_1), .CK (wb_clk_i), .D (
                        wbd_dat_i[1]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_1)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_1 (.Q (cdata_1), .CK (wb_clk_i), .D (nx5934), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5935 (.Y (nx5934), .A0 (nx7519), .A1 (nx7555), .B0 (
                      nx7699)) ;
    NAND2_X0P5A_A12TS ix7700 (.Y (nx7699), .A (cdata_1), .B (nx7555)) ;
    NOR2_X0P5A_A12TS ix261 (.Y (nx260), .A (cdone), .B (dack_ir)) ;
    OAI21_X0P5M_A12TS ix1061 (.Y (nx1492), .A0 (op1_n_7), .A1 (nx7704), .B0 (
                      nx7751)) ;
    AOI222_X0P5M_A12TS ix7705 (.Y (nx7704), .A0 (cdata_5), .A1 (nx270), .B0 (
                       ddat_ir_5), .B1 (dack_ir), .C0 (nx1480), .C1 (nx260)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_5 (.Q (cdata_5), .CK (wb_clk_i), .D (nx6034), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6035 (.Y (nx6034), .A0 (nx7708), .A1 (nx7555), .B0 (
                      nx7710)) ;
    AOI32_X0P5M_A12TS ix7709 (.Y (nx7708), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[5]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7711 (.Y (nx7710), .A (cdata_5), .B (nx7555)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_5 (.Q (ddat_ir_5), .CK (wb_clk_i), .D (
                        wbd_dat_i[5]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_5)) ;
    MXIT2_X0P5M_A12TS ix7715 (.Y (nx7714), .A (idat_old_21), .B (idat_old_29), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_21 (.Q (idat_old_21), .CK (wb_clk_i), .D (
                        idat_cur_21), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_21)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_21 (.Q (idat_cur_21), .CK (wb_clk_i), .D (
                       nx5994), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5995 (.Y (nx5994), .A0 (nx7719), .A1 (NOT_nx5673), .B0 (
                      nx7721)) ;
    AOI32_X0P5M_A12TS ix7720 (.Y (nx7719), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[21]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7722 (.Y (nx7721), .A (idat_cur_21), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_29 (.Q (idat_old_29), .CK (wb_clk_i), .D (
                        idat_cur_29), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_29)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_29 (.Q (idat_cur_29), .CK (wb_clk_i), .D (
                       nx6014), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6015 (.Y (nx6014), .A0 (nx7726), .A1 (NOT_nx5673), .B0 (
                      nx7728)) ;
    AOI32_X0P5M_A12TS ix7727 (.Y (nx7726), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[29]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7729 (.Y (nx7728), .A (idat_cur_29), .B (NOT_nx5673)) ;
    INV_X0P5B_A12TS ix7731 (.Y (nx7730), .A (idat_old_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_5 (.Q (idat_old_5), .CK (wb_clk_i), .D (
                        idat_cur_5), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_5)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_5 (.Q (idat_cur_5), .CK (wb_clk_i), .D (
                       nx5974), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5975 (.Y (nx5974), .A0 (nx7708), .A1 (NOT_nx5673), .B0 (
                      nx7735)) ;
    NAND2_X0P5A_A12TS ix7736 (.Y (nx7735), .A (idat_cur_5), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_13 (.Q (idat_old_13), .CK (wb_clk_i), .D (
                        idat_cur_13), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_13)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_13 (.Q (idat_cur_13), .CK (wb_clk_i), .D (
                       nx5954), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5955 (.Y (nx5954), .A0 (nx7742), .A1 (NOT_nx5673), .B0 (
                      nx7744)) ;
    AOI32_X0P5M_A12TS ix7743 (.Y (nx7742), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[13]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7745 (.Y (nx7744), .A (idat_cur_13), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix467 (.Y (nx466), .A0 (nx7747), .A1 (nx7670), .B0 (nx7749
                      ), .B1 (nx7685)) ;
    INV_X0P5B_A12TS ix7748 (.Y (nx7747), .A (idat_cur_13)) ;
    MXIT2_X0P5M_A12TS ix7750 (.Y (nx7749), .A (idat_cur_5), .B (idat_cur_13), .S0 (
                      op_pos_0)) ;
    AO21A1AI2_X0P5M_A12TS ix7752 (.Y (nx7751), .A0 (op1_n_4), .A1 (nx7808), .B0 (
                          op1_n_0), .C0 (nx7704)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_4 (.Q (ddat_ir_4), .CK (wb_clk_i), .D (
                        wbd_dat_i[4]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_4)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_4 (.Q (cdata_4), .CK (wb_clk_i), .D (nx6214), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6215 (.Y (nx6214), .A0 (nx7761), .A1 (nx7555), .B0 (
                      nx7763)) ;
    AOI32_X0P5M_A12TS ix7762 (.Y (nx7761), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[4]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7764 (.Y (nx7763), .A (cdata_4), .B (nx7555)) ;
    OAI211_X0P5M_A12TS ix1276 (.Y (nx1485), .A0 (nx7766), .A1 (nx7778), .B0 (
                       nx7780), .C0 (nx7785)) ;
    MXIT2_X0P5M_A12TS ix7767 (.Y (nx7766), .A (idat_cur_4), .B (idat_cur_12), .S0 (
                      op_pos_0)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_4 (.Q (idat_cur_4), .CK (wb_clk_i), .D (
                       nx6194), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6195 (.Y (nx6194), .A0 (nx7761), .A1 (NOT_nx5673), .B0 (
                      nx7770)) ;
    NAND2_X0P5A_A12TS ix7771 (.Y (nx7770), .A (idat_cur_4), .B (NOT_nx5673)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_12 (.Q (idat_cur_12), .CK (wb_clk_i), .D (
                       nx6134), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6135 (.Y (nx6134), .A0 (nx7774), .A1 (NOT_nx5673), .B0 (
                      nx7776)) ;
    AOI32_X0P5M_A12TS ix7775 (.Y (nx7774), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[12]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7777 (.Y (nx7776), .A (idat_cur_12), .B (NOT_nx5673)) ;
    NAND2_X0P5A_A12TS ix7779 (.Y (nx7778), .A (op_pos_2), .B (nx7595)) ;
    AOI31_X0P5M_A12TS ix7786 (.Y (nx7785), .A0 (op_pos_1), .A1 (idat_cur_12), .A2 (
                      op_pos_2), .B0 (nx1483)) ;
    OA21A1OI2_X0P5M_A12TS ix1277 (.Y (nx1483), .A0 (nx7595), .A1 (nx7788), .B0 (
                          nx7804), .C0 (op_pos_2)) ;
    MXIT2_X0P5M_A12TS ix7789 (.Y (nx7788), .A (idat_old_20), .B (idat_old_28), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_20 (.Q (idat_old_20), .CK (wb_clk_i), .D (
                        idat_cur_20), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_20)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_20 (.Q (idat_cur_20), .CK (wb_clk_i), .D (
                       nx6144), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6145 (.Y (nx6144), .A0 (nx7793), .A1 (NOT_nx5673), .B0 (
                      nx7795)) ;
    AOI32_X0P5M_A12TS ix7794 (.Y (nx7793), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[20]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7796 (.Y (nx7795), .A (idat_cur_20), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_28 (.Q (idat_old_28), .CK (wb_clk_i), .D (
                        idat_cur_28), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_28)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_28 (.Q (idat_cur_28), .CK (wb_clk_i), .D (
                       nx6164), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6165 (.Y (nx6164), .A0 (nx7800), .A1 (NOT_nx5673), .B0 (
                      nx7802)) ;
    AOI32_X0P5M_A12TS ix7801 (.Y (nx7800), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[28]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7803 (.Y (nx7802), .A (idat_cur_28), .B (NOT_nx5673)) ;
    AOI32_X0P5M_A12TS ix7805 (.Y (nx7804), .A0 (op_pos_0), .A1 (idat_old_12), .A2 (
                      nx7595), .B0 (idat_old_4), .B1 (nx7665)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_12 (.Q (idat_old_12), .CK (wb_clk_i), .D (
                        idat_cur_12), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_12)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_4 (.Q (idat_old_4), .CK (wb_clk_i), .D (
                        idat_cur_4), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_4)) ;
    AOI222_X0P5M_A12TS ix7809 (.Y (nx7808), .A0 (cdata_2), .A1 (nx270), .B0 (
                       ddat_ir_2), .B1 (dack_ir), .C0 (nx1489), .C1 (nx260)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_2 (.Q (cdata_2), .CK (wb_clk_i), .D (nx6414), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6415 (.Y (nx6414), .A0 (nx7812), .A1 (nx7555), .B0 (
                      nx7814)) ;
    AOI32_X0P5M_A12TS ix7813 (.Y (nx7812), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[2]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7815 (.Y (nx7814), .A (cdata_2), .B (nx7555)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_2 (.Q (ddat_ir_2), .CK (wb_clk_i), .D (
                        wbd_dat_i[2]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_2)) ;
    MXIT2_X0P5M_A12TS ix7819 (.Y (nx7818), .A (idat_old_18), .B (idat_old_26), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_18 (.Q (idat_old_18), .CK (wb_clk_i), .D (
                        idat_cur_18), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_18)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_18 (.Q (idat_cur_18), .CK (wb_clk_i), .D (
                       nx6374), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6375 (.Y (nx6374), .A0 (nx7823), .A1 (NOT_nx5673), .B0 (
                      nx7825)) ;
    AOI32_X0P5M_A12TS ix7824 (.Y (nx7823), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[18]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7826 (.Y (nx7825), .A (idat_cur_18), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_26 (.Q (idat_old_26), .CK (wb_clk_i), .D (
                        idat_cur_26), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_26)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_26 (.Q (idat_cur_26), .CK (wb_clk_i), .D (
                       nx6394), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6395 (.Y (nx6394), .A0 (nx7830), .A1 (NOT_nx5673), .B0 (
                      nx7832)) ;
    AOI32_X0P5M_A12TS ix7831 (.Y (nx7830), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[26]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7833 (.Y (nx7832), .A (idat_cur_26), .B (NOT_nx5673)) ;
    INV_X0P5B_A12TS ix7835 (.Y (nx7834), .A (idat_old_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_2 (.Q (idat_old_2), .CK (wb_clk_i), .D (
                        idat_cur_2), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_2)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_2 (.Q (idat_cur_2), .CK (wb_clk_i), .D (
                       nx6354), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6355 (.Y (nx6354), .A0 (nx7812), .A1 (NOT_nx5673), .B0 (
                      nx7839)) ;
    NAND2_X0P5A_A12TS ix7840 (.Y (nx7839), .A (idat_cur_2), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_10 (.Q (idat_old_10), .CK (wb_clk_i), .D (
                        idat_cur_10), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_10)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_10 (.Q (idat_cur_10), .CK (wb_clk_i), .D (
                       nx6334), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6335 (.Y (nx6334), .A0 (nx7846), .A1 (NOT_nx5673), .B0 (
                      nx7848)) ;
    AOI32_X0P5M_A12TS ix7847 (.Y (nx7846), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[10]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7849 (.Y (nx7848), .A (idat_cur_10), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix1278 (.Y (nx1487), .A0 (nx7851), .A1 (nx7670), .B0 (
                      nx7853), .B1 (nx7685)) ;
    INV_X0P5B_A12TS ix7852 (.Y (nx7851), .A (idat_cur_10)) ;
    MXIT2_X0P5M_A12TS ix7854 (.Y (nx7853), .A (idat_cur_2), .B (idat_cur_10), .S0 (
                      op_pos_0)) ;
    OAI222_X0P5M_A12TS ix1279 (.Y (op1_n_0), .A0 (nx7856), .A1 (nx7572), .B0 (
                       nx7864), .B1 (nx7575), .C0 (nx7867), .C1 (nx7687)) ;
    INV_X0P5B_A12TS ix7857 (.Y (nx7856), .A (cdata_0)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_0 (.Q (cdata_0), .CK (wb_clk_i), .D (nx6114), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6115 (.Y (nx6114), .A0 (nx7860), .A1 (nx7555), .B0 (
                      nx7862)) ;
    AOI32_X0P5M_A12TS ix7861 (.Y (nx7860), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[0]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7863 (.Y (nx7862), .A (cdata_0), .B (nx7555)) ;
    INV_X0P5B_A12TS ix7865 (.Y (nx7864), .A (ddat_ir_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_0 (.Q (ddat_ir_0), .CK (wb_clk_i), .D (
                        wbd_dat_i[0]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_0)) ;
    AOI211_X0P5M_A12TS ix7868 (.Y (nx7867), .A0 (idat_old_8), .A1 (nx5675), .B0 (
                       nx618), .C0 (nx1481)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_8 (.Q (idat_old_8), .CK (wb_clk_i), .D (
                        idat_cur_8), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_8)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_8 (.Q (idat_cur_8), .CK (wb_clk_i), .D (
                       nx6054), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6055 (.Y (nx6054), .A0 (nx7872), .A1 (NOT_nx5673), .B0 (
                      nx7874)) ;
    AOI32_X0P5M_A12TS ix7873 (.Y (nx7872), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[8]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7875 (.Y (nx7874), .A (idat_cur_8), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix1280 (.Y (nx618), .A0 (nx7877), .A1 (nx7654), .B0 (
                      nx7893), .B1 (nx7663)) ;
    MXIT2_X0P5M_A12TS ix7878 (.Y (nx7877), .A (idat_old_16), .B (idat_old_24), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_16 (.Q (idat_old_16), .CK (wb_clk_i), .D (
                        idat_cur_16), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_16)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_16 (.Q (idat_cur_16), .CK (wb_clk_i), .D (
                       nx6524), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6525 (.Y (nx6524), .A0 (nx7882), .A1 (NOT_nx5673), .B0 (
                      nx7884)) ;
    AOI32_X0P5M_A12TS ix7883 (.Y (nx7882), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[16]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7885 (.Y (nx7884), .A (idat_cur_16), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_24 (.Q (idat_old_24), .CK (wb_clk_i), .D (
                        idat_cur_24), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_24)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_24 (.Q (idat_cur_24), .CK (wb_clk_i), .D (
                       nx6094), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6095 (.Y (nx6094), .A0 (nx7889), .A1 (NOT_nx5673), .B0 (
                      nx7891)) ;
    AOI32_X0P5M_A12TS ix7890 (.Y (nx7889), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[24]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7892 (.Y (nx7891), .A (idat_cur_24), .B (NOT_nx5673)) ;
    INV_X0P5B_A12TS ix7894 (.Y (nx7893), .A (idat_old_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_0 (.Q (idat_old_0), .CK (wb_clk_i), .D (
                        idat_cur_0), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_0)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_0 (.Q (idat_cur_0), .CK (wb_clk_i), .D (
                       nx6074), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6075 (.Y (nx6074), .A0 (nx7860), .A1 (NOT_nx5673), .B0 (
                      nx7898)) ;
    NAND2_X0P5A_A12TS ix7899 (.Y (nx7898), .A (idat_cur_0), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix1281 (.Y (nx1481), .A0 (nx7901), .A1 (nx7670), .B0 (
                      nx7903), .B1 (nx7685)) ;
    INV_X0P5B_A12TS ix7902 (.Y (nx7901), .A (idat_cur_8)) ;
    MXIT2_X0P5M_A12TS ix7904 (.Y (nx7903), .A (idat_cur_0), .B (idat_cur_8), .S0 (
                      op_pos_0)) ;
    OAI222_X0P5M_A12TS ix1282 (.Y (op1_n_6), .A0 (nx7908), .A1 (nx7572), .B0 (
                       nx7916), .B1 (nx7575), .C0 (nx7919), .C1 (nx7687)) ;
    INV_X0P5B_A12TS ix7909 (.Y (nx7908), .A (cdata_6)) ;
    DFFRPQ_X0P5M_A12TS reg_cdata_6 (.Q (cdata_6), .CK (wb_clk_i), .D (nx6314), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6315 (.Y (nx6314), .A0 (nx7912), .A1 (nx7555), .B0 (
                      nx7914)) ;
    AOI32_X0P5M_A12TS ix7913 (.Y (nx7912), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[6]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7915 (.Y (nx7914), .A (cdata_6), .B (nx7555)) ;
    INV_X0P5B_A12TS ix7917 (.Y (nx7916), .A (ddat_ir_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_ddat_ir_6 (.Q (ddat_ir_6), .CK (wb_clk_i), .D (
                        wbd_dat_i[6]), .R (wb_rst_i), .SE (NOT_dack_i), .SI (
                        ddat_ir_6)) ;
    AOI211_X0P5M_A12TS ix7920 (.Y (nx7919), .A0 (idat_old_14), .A1 (nx5675), .B0 (
                       nx880), .C0 (nx828)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_14 (.Q (idat_old_14), .CK (wb_clk_i), .D (
                        idat_cur_14), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_14)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_14 (.Q (idat_cur_14), .CK (wb_clk_i), .D (
                       nx6234), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6235 (.Y (nx6234), .A0 (nx7924), .A1 (NOT_nx5673), .B0 (
                      nx7926)) ;
    AOI32_X0P5M_A12TS ix7925 (.Y (nx7924), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[14]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7927 (.Y (nx7926), .A (idat_cur_14), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix1284 (.Y (nx880), .A0 (nx7929), .A1 (nx7654), .B0 (
                      nx7945), .B1 (nx7663)) ;
    MXIT2_X0P5M_A12TS ix7930 (.Y (nx7929), .A (idat_old_22), .B (idat_old_30), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_22 (.Q (idat_old_22), .CK (wb_clk_i), .D (
                        idat_cur_22), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_22)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_22 (.Q (idat_cur_22), .CK (wb_clk_i), .D (
                       nx6274), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6275 (.Y (nx6274), .A0 (nx7934), .A1 (NOT_nx5673), .B0 (
                      nx7936)) ;
    AOI32_X0P5M_A12TS ix7935 (.Y (nx7934), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[22]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7937 (.Y (nx7936), .A (idat_cur_22), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_30 (.Q (idat_old_30), .CK (wb_clk_i), .D (
                        idat_cur_30), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_30)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_30 (.Q (idat_cur_30), .CK (wb_clk_i), .D (
                       nx6294), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6295 (.Y (nx6294), .A0 (nx7941), .A1 (NOT_nx5673), .B0 (
                      nx7943)) ;
    AOI32_X0P5M_A12TS ix7942 (.Y (nx7941), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[30]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7944 (.Y (nx7943), .A (idat_cur_30), .B (NOT_nx5673)) ;
    INV_X0P5B_A12TS ix7946 (.Y (nx7945), .A (idat_old_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_6 (.Q (idat_old_6), .CK (wb_clk_i), .D (
                        idat_cur_6), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_6)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_6 (.Q (idat_cur_6), .CK (wb_clk_i), .D (
                       nx6254), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6255 (.Y (nx6254), .A0 (nx7912), .A1 (NOT_nx5673), .B0 (
                      nx7950)) ;
    NAND2_X0P5A_A12TS ix7951 (.Y (nx7950), .A (idat_cur_6), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix829 (.Y (nx828), .A0 (nx7953), .A1 (nx7670), .B0 (nx7955
                      ), .B1 (nx7685)) ;
    INV_X0P5B_A12TS ix7954 (.Y (nx7953), .A (idat_cur_14)) ;
    MXIT2_X0P5M_A12TS ix7956 (.Y (nx7955), .A (idat_cur_6), .B (idat_cur_14), .S0 (
                      op_pos_0)) ;
    AOI21_X0P5M_A12TS ix7959 (.Y (nx7958), .A0 (op1_n_2), .A1 (op1_n_1), .B0 (
                      op1_n_3)) ;
    AOI211_X0P5M_A12TS ix7966 (.Y (nx7965), .A0 (idat_old_10), .A1 (nx5675), .B0 (
                       nx1488), .C0 (nx1487)) ;
    OAI22_X0P5M_A12TS ix1005 (.Y (nx1488), .A0 (nx7818), .A1 (nx7654), .B0 (
                      nx7834), .B1 (nx7663)) ;
    AOI211_X0P5M_A12TS ix7976 (.Y (nx7975), .A0 (idat_old_13), .A1 (nx5675), .B0 (
                       nx518), .C0 (nx466)) ;
    OAI22_X0P5M_A12TS ix519 (.Y (nx518), .A0 (nx7714), .A1 (nx7654), .B0 (nx7730
                      ), .B1 (nx7663)) ;
    AOI222_X0P5M_A12TS ix7982 (.Y (nx7981), .A0 (cdata_7), .A1 (nx270), .B0 (
                       ddat_ir_7), .B1 (dack_ir), .C0 (nx1493), .C1 (nx260)) ;
    MXIT2_X0P5M_A12TS ix7985 (.Y (nx7984), .A (idat_old_23), .B (idat_old_31), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_23 (.Q (idat_old_23), .CK (wb_clk_i), .D (
                        idat_cur_23), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_23)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_23 (.Q (idat_cur_23), .CK (wb_clk_i), .D (
                       nx6454), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6455 (.Y (nx6454), .A0 (nx7989), .A1 (NOT_nx5673), .B0 (
                      nx7991)) ;
    AOI32_X0P5M_A12TS ix7990 (.Y (nx7989), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[23]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7992 (.Y (nx7991), .A (idat_cur_23), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_31 (.Q (idat_old_31), .CK (wb_clk_i), .D (
                        idat_cur_31), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_31)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_31 (.Q (idat_cur_31), .CK (wb_clk_i), .D (
                       nx6474), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6475 (.Y (nx6474), .A0 (nx7996), .A1 (NOT_nx5673), .B0 (
                      nx7998)) ;
    AOI32_X0P5M_A12TS ix7997 (.Y (nx7996), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[31]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix7999 (.Y (nx7998), .A (idat_cur_31), .B (NOT_nx5673)) ;
    INV_X0P5B_A12TS ix8001 (.Y (nx8000), .A (idat_old_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_7 (.Q (idat_old_7), .CK (wb_clk_i), .D (
                        idat_cur_7), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_7)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_7 (.Q (idat_cur_7), .CK (wb_clk_i), .D (
                       nx6434), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6435 (.Y (nx6434), .A0 (nx7553), .A1 (NOT_nx5673), .B0 (
                      nx8005)) ;
    NAND2_X0P5A_A12TS ix8006 (.Y (nx8005), .A (idat_cur_7), .B (NOT_nx5673)) ;
    OAI22_X0P5M_A12TS ix1115 (.Y (nx1114), .A0 (nx8010), .A1 (nx7670), .B0 (
                      nx8012), .B1 (nx7685)) ;
    INV_X0P5B_A12TS ix8011 (.Y (nx8010), .A (idat_cur_15)) ;
    MXIT2_X0P5M_A12TS ix8013 (.Y (nx8012), .A (idat_cur_7), .B (idat_cur_15), .S0 (
                      op_pos_0)) ;
    AOI211_X0P5M_A12TS ix1245 (.Y (nx1497), .A0 (nx8017), .A1 (op1_n_0), .B0 (
                       op1_n_3), .C0 (nx8019)) ;
    OA21A1OI2_X0P5M_A12TS ix1319 (.Y (nx1318), .A0 (op1_n_7), .A1 (nx8022), .B0 (
                          nx8025), .C0 (op1_n_6)) ;
    NOR2_X0P5A_A12TS ix8023 (.Y (nx8022), .A (nx1276), .B (op1_n_1)) ;
    AOI21_X0P5M_A12TS ix1285 (.Y (nx1276), .A0 (op1_n_2), .A1 (op1_n_5), .B0 (
                      op1_n_0)) ;
    OA21A1OI2_X0P5M_A12TS ix8026 (.Y (nx8025), .A0 (nx1306), .A1 (op1_n_3), .B0 (
                          op1_n_4), .C0 (nx1500)) ;
    NOR3_X0P5A_A12TS ix1307 (.Y (nx1306), .A (nx8028), .B (op1_n_1), .C (op1_n_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix1286 (.Y (nx1500), .A0 (op1_n_4), .A1 (nx8031), .B0 (
                          nx778), .C0 (nx8019)) ;
    AOI32_X0P5M_A12TS ix8036 (.Y (nx8035), .A0 (op1_n_1), .A1 (nx7704), .A2 (
                      op1_n_2), .B0 (op1_n_3), .B1 (nx778)) ;
    AOI31_X0P5M_A12TS ix8038 (.Y (nx8037), .A0 (nx8014), .A1 (op1_n_7), .A2 (
                      op1_n_3), .B0 (nx1496)) ;
    NOR3_X0P5A_A12TS ix1287 (.Y (nx1496), .A (nx8040), .B (op1_n_3), .C (nx8043)
                     ) ;
    AOI22_X0P5M_A12TS ix8041 (.Y (nx8040), .A0 (nx7808), .A1 (op1_n_0), .B0 (
                      op1_n_4), .B1 (nx1491)) ;
    AOI222_X0P5M_A12TS ix8044 (.Y (nx8043), .A0 (cdata_1), .A1 (nx270), .B0 (
                       ddat_ir_1), .B1 (dack_ir), .C0 (nx1478), .C1 (nx260)) ;
    OAI31_X0P5M_A12TS ix1043 (.Y (nx1042), .A0 (nx8046), .A1 (op1_n_3), .A2 (
                      op1_n_2), .B0 (nx8049)) ;
    AOI31_X0P5M_A12TS ix8047 (.Y (nx8046), .A0 (nx778), .A1 (nx7981), .A2 (
                      op1_n_6), .B0 (nx1482)) ;
    NOR3_X0P5A_A12TS ix1288 (.Y (nx1482), .A (nx416), .B (op1_n_5), .C (op1_n_0)
                     ) ;
    OAI211_X0P5M_A12TS ix8050 (.Y (nx8049), .A0 (op1_n_3), .A1 (op1_n_2), .B0 (
                       op1_n_7), .C0 (nx1038)) ;
    NOR2_X0P5A_A12TS ix1039 (.Y (nx1038), .A (op1_n_6), .B (nx778)) ;
    XOR2_X0P5M_A12TS ix1355 (.Y (nx1354), .A (nx1352), .B (op_pos_2)) ;
    CGENI_X1M_A12TS ix1353 (.CON (nx1352), .A (nx7541), .B (nx7595), .CI (nx7613
                    )) ;
    OAI22_X0P5M_A12TS ix1167 (.Y (nx1166), .A0 (nx7984), .A1 (nx7654), .B0 (
                      nx8000), .B1 (nx7663)) ;
    OA21A1OI2_X0P5M_A12TS ix8057 (.Y (nx8056), .A0 (nx1499), .A1 (nx1498), .B0 (
                          op1_n_6), .C0 (nx1318)) ;
    OAI22_X0P5M_A12TS ix1289 (.Y (nx1499), .A0 (op1_n_0), .A1 (nx8059), .B0 (
                      op1_n_4), .B1 (nx7958)) ;
    AOI222_X0P5M_A12TS ix8068 (.Y (nx8067), .A0 (cdata_4), .A1 (nx270), .B0 (
                       ddat_ir_4), .B1 (dack_ir), .C0 (nx1485), .C1 (nx260)) ;
    NOR2_X0P5A_A12TS ix8070 (.Y (nx8069), .A (pc_wr_r2), .B (rd)) ;
    XOR2_X0P5M_A12TS ix8072 (.Y (nx8071), .A (op_pos_1), .B (nx7613)) ;
    NAND2_X0P5A_A12TS ix8074 (.Y (nx8073), .A (op_pos_1), .B (nx8069)) ;
    NAND2_X0P5A_A12TS ix8076 (.Y (nx8075), .A (idat_cur_1), .B (NOT_nx5673)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_9 (.Q (idat_cur_9), .CK (wb_clk_i), .D (
                       nx5854), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5855 (.Y (nx5854), .A0 (nx8079), .A1 (NOT_nx5673), .B0 (
                      nx8081)) ;
    AOI32_X0P5M_A12TS ix8080 (.Y (nx8079), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[9]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix8082 (.Y (nx8081), .A (idat_cur_9), .B (NOT_nx5673)) ;
    AOI31_X0P5M_A12TS ix8084 (.Y (nx8083), .A0 (op_pos_1), .A1 (idat_cur_9), .A2 (
                      op_pos_2), .B0 (nx378)) ;
    OA21A1OI2_X0P5M_A12TS ix379 (.Y (nx378), .A0 (nx7595), .A1 (nx8086), .B0 (
                          nx8102), .C0 (op_pos_2)) ;
    MXIT2_X0P5M_A12TS ix8087 (.Y (nx8086), .A (idat_old_17), .B (idat_old_25), .S0 (
                      op_pos_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_17 (.Q (idat_old_17), .CK (wb_clk_i), .D (
                        idat_cur_17), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_17)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_17 (.Q (idat_cur_17), .CK (wb_clk_i), .D (
                       nx5864), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5865 (.Y (nx5864), .A0 (nx8091), .A1 (NOT_nx5673), .B0 (
                      nx8093)) ;
    AOI32_X0P5M_A12TS ix8092 (.Y (nx8091), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[17]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix8094 (.Y (nx8093), .A (idat_cur_17), .B (NOT_nx5673)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_25 (.Q (idat_old_25), .CK (wb_clk_i), .D (
                        idat_cur_25), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_25)) ;
    DFFRPQ_X0P5M_A12TS reg_idat_cur_25 (.Q (idat_cur_25), .CK (wb_clk_i), .D (
                       nx5884), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5885 (.Y (nx5884), .A0 (nx8098), .A1 (NOT_nx5673), .B0 (
                      nx8100)) ;
    AOI32_X0P5M_A12TS ix8099 (.Y (nx8098), .A0 (ea_int), .A1 (ea_int), .A2 (
                      ea_in), .B0 (wbi_dat_i[25]), .B1 (nx7521)) ;
    NAND2_X0P5A_A12TS ix8101 (.Y (nx8100), .A (idat_cur_25), .B (NOT_nx5673)) ;
    AOI32_X0P5M_A12TS ix8103 (.Y (nx8102), .A0 (op_pos_0), .A1 (idat_old_9), .A2 (
                      nx7595), .B0 (idat_old_1), .B1 (nx7665)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_9 (.Q (idat_old_9), .CK (wb_clk_i), .D (
                        idat_cur_9), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_9)) ;
    SDFFRPQ_X0P5M_A12TS reg_idat_old_1 (.Q (idat_old_1), .CK (wb_clk_i), .D (
                        idat_cur_1), .R (wb_rst_i), .SE (NOT_nx5673), .SI (
                        idat_old_1)) ;
    NAND2_X0P5A_A12TS ix8107 (.Y (nx8106), .A (nx7965), .B (nx7628)) ;
    NAND4B_X0P5M_A12TS ix8109 (.Y (nx8108), .AN (mem_wait), .B (nx7919), .C (
                       nx3944), .D (nx7581)) ;
    OR3_X0P5M_A12TS ix3959 (.Y (mem_wait), .A (wbd_stb_o), .B (imem_wait), .C (
                    pc_wr_r2)) ;
    DFFRPQ_X0P5M_A12TS reg_int_ack (.Q (int_ack), .CK (wb_clk_i), .D (nx3924), .R (
                       wb_rst_i)) ;
    NOR2B_X0P7M_A12TS ix3925 (.Y (nx3924), .AN (int_ack_buff), .B (int_ack_t)) ;
    DFFRPQ_X0P5M_A12TS reg_int_ack_buff (.Q (int_ack_buff), .CK (wb_clk_i), .D (
                       int_ack_t), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_0 (.Q (wbd_dat_o[0]), .CK (wb_clk_i), .D (
                       nx7104), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7105 (.Y (nx7104), .A0N (nx8119), .B0 (wbd_dat_o[0]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8120 (.Y (nx8119), .A (acc_0), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_1 (.Q (wbd_dat_o[1]), .CK (wb_clk_i), .D (
                       nx7114), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7115 (.Y (nx7114), .A0N (nx8123), .B0 (wbd_dat_o[1]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8124 (.Y (nx8123), .A (acc_1), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_2 (.Q (wbd_dat_o[2]), .CK (wb_clk_i), .D (
                       nx7124), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7125 (.Y (nx7124), .A0N (nx8127), .B0 (wbd_dat_o[2]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8128 (.Y (nx8127), .A (acc_2), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_3 (.Q (wbd_dat_o[3]), .CK (wb_clk_i), .D (
                       nx7134), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7135 (.Y (nx7134), .A0N (nx8131), .B0 (wbd_dat_o[3]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8132 (.Y (nx8131), .A (acc_3), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_4 (.Q (wbd_dat_o[4]), .CK (wb_clk_i), .D (
                       nx7144), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7145 (.Y (nx7144), .A0N (nx8135), .B0 (wbd_dat_o[4]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8136 (.Y (nx8135), .A (acc_4), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_5 (.Q (wbd_dat_o[5]), .CK (wb_clk_i), .D (
                       nx7154), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7155 (.Y (nx7154), .A0N (nx8139), .B0 (wbd_dat_o[5]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8140 (.Y (nx8139), .A (acc_5), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_6 (.Q (wbd_dat_o[6]), .CK (wb_clk_i), .D (
                       nx7164), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7165 (.Y (nx7164), .A0N (nx8143), .B0 (wbd_dat_o[6]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8144 (.Y (nx8143), .A (acc_6), .B (mem_act_0), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ddat_o_7 (.Q (wbd_dat_o[7]), .CK (wb_clk_i), .D (
                       nx7174), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7175 (.Y (nx7174), .A0N (nx8147), .B0 (wbd_dat_o[7]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8148 (.Y (nx8147), .A (mem_act_0), .B (acc_7), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dwe_o (.Q (wbd_we_o), .CK (wb_clk_i), .D (nx3976), .R (
                       wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix3977 (.Y (nx3976), .A (nx7568), .B (wbd_ack_i)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_0 (.Q (wbd_adr_o[0]), .CK (wb_clk_i), .D (
                        nx4036), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[0])) ;
    NAND2_X0P5A_A12TS ix8156 (.Y (nx8155), .A (dptr_lo_0), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_1 (.Q (wbd_adr_o[1]), .CK (wb_clk_i), .D (
                        nx4048), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[1])) ;
    NAND2_X0P5A_A12TS ix8162 (.Y (nx8161), .A (dptr_lo_1), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_2 (.Q (wbd_adr_o[2]), .CK (wb_clk_i), .D (
                        nx4060), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[2])) ;
    NAND2_X0P5A_A12TS ix8168 (.Y (nx8167), .A (dptr_lo_2), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_3 (.Q (wbd_adr_o[3]), .CK (wb_clk_i), .D (
                        nx4072), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[3])) ;
    NAND2_X0P5A_A12TS ix8174 (.Y (nx8173), .A (dptr_lo_3), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_4 (.Q (wbd_adr_o[4]), .CK (wb_clk_i), .D (
                        nx4084), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[4])) ;
    NAND2_X0P5A_A12TS ix8180 (.Y (nx8179), .A (dptr_lo_4), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_5 (.Q (wbd_adr_o[5]), .CK (wb_clk_i), .D (
                        nx4096), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[5])) ;
    INV_X0P5B_A12TS ix8184 (.Y (nx8183), .A (ri_5)) ;
    NAND2_X0P5A_A12TS ix8186 (.Y (nx8185), .A (dptr_lo_5), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_6 (.Q (wbd_adr_o[6]), .CK (wb_clk_i), .D (
                        nx4108), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[6])) ;
    INV_X0P5B_A12TS ix8190 (.Y (nx8189), .A (ri_6)) ;
    NAND2_X0P5A_A12TS ix8192 (.Y (nx8191), .A (dptr_lo_6), .B (nx7566)) ;
    SDFFRPQ_X0P5M_A12TS reg_dadr_ot_7 (.Q (wbd_adr_o[7]), .CK (wb_clk_i), .D (
                        nx4120), .R (wb_rst_i), .SE (wbd_ack_i), .SI (
                        wbd_adr_o[7])) ;
    NAND2_X0P5A_A12TS ix8198 (.Y (nx8197), .A (nx7566), .B (dptr_lo_7)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_8 (.Q (wbd_adr_o[8]), .CK (wb_clk_i), .D (
                       nx7264), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7265 (.Y (nx7264), .A0N (nx8201), .B0 (wbd_adr_o[8]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8202 (.Y (nx8201), .A (dptr_hi_0), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_9 (.Q (wbd_adr_o[9]), .CK (wb_clk_i), .D (
                       nx7274), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7275 (.Y (nx7274), .A0N (nx8205), .B0 (wbd_adr_o[9]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8206 (.Y (nx8205), .A (dptr_hi_1), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_10 (.Q (wbd_adr_o[10]), .CK (wb_clk_i), .D (
                       nx7284), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7285 (.Y (nx7284), .A0N (nx8209), .B0 (wbd_adr_o[10]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8210 (.Y (nx8209), .A (dptr_hi_2), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_11 (.Q (wbd_adr_o[11]), .CK (wb_clk_i), .D (
                       nx7294), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7295 (.Y (nx7294), .A0N (nx8213), .B0 (wbd_adr_o[11]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8214 (.Y (nx8213), .A (dptr_hi_3), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_12 (.Q (wbd_adr_o[12]), .CK (wb_clk_i), .D (
                       nx7304), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7305 (.Y (nx7304), .A0N (nx8217), .B0 (wbd_adr_o[12]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8218 (.Y (nx8217), .A (dptr_hi_4), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_13 (.Q (wbd_adr_o[13]), .CK (wb_clk_i), .D (
                       nx7314), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7315 (.Y (nx7314), .A0N (nx8221), .B0 (wbd_adr_o[13]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8222 (.Y (nx8221), .A (dptr_hi_5), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_14 (.Q (wbd_adr_o[14]), .CK (wb_clk_i), .D (
                       nx7324), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7325 (.Y (nx7324), .A0N (nx8225), .B0 (wbd_adr_o[14]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8226 (.Y (nx8225), .A (dptr_hi_6), .B (nx7566), .C (
                      NOT_dack_i)) ;
    DFFRPQ_X0P5M_A12TS reg_dadr_ot_15 (.Q (wbd_adr_o[15]), .CK (wb_clk_i), .D (
                       nx7334), .R (wb_rst_i)) ;
    AO1B2_X0P5M_A12TS ix7335 (.Y (nx7334), .A0N (nx8229), .B0 (wbd_adr_o[15]), .B1 (
                      wbd_ack_i)) ;
    NAND3_X0P5A_A12TS ix8230 (.Y (nx8229), .A (dptr_hi_7), .B (nx7566), .C (
                      NOT_dack_i)) ;
    OAI21_X0P5M_A12TS ix1593 (.Y (op3_n_0), .A0 (rd), .A1 (nx8235), .B0 (nx8253)
                      ) ;
    INV_X0P5B_A12TS ix8236 (.Y (nx8235), .A (op3_buff_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_0 (.Q (op3_buff_0), .CK (wb_clk_i), .D (
                        nx1580), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_0)
                        ) ;
    OAI211_X0P5M_A12TS ix1581 (.Y (nx1580), .A0 (nx7877), .A1 (nx7593), .B0 (
                       nx8239), .C0 (nx8246)) ;
    AOI22_X0P5M_A12TS ix8240 (.Y (nx8239), .A0 (int_vec_buff_0), .A1 (nx1473), .B0 (
                      nx576), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_0 (.Q (int_vec_buff_0), .CK (wb_clk_i)
                        , .D (int_src_1), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_0)) ;
    AOI22_X0P5M_A12TS ix8247 (.Y (nx8246), .A0 (idat_cur_16), .A1 (nx1503), .B0 (
                      idat_cur_24), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8254 (.Y (nx8253), .A (rd), .B (nx1580)) ;
    OAI21_X0P5M_A12TS ix1695 (.Y (op3_n_1), .A0 (rd), .A1 (nx8256), .B0 (nx8270)
                      ) ;
    INV_X0P5B_A12TS ix8257 (.Y (nx8256), .A (op3_buff_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_1 (.Q (op3_buff_1), .CK (wb_clk_i), .D (
                        nx1682), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_1)
                        ) ;
    OAI211_X0P5M_A12TS ix1683 (.Y (nx1682), .A0 (nx8086), .A1 (nx7593), .B0 (
                       nx8260), .C0 (nx8268)) ;
    AOI22_X0P5M_A12TS ix8261 (.Y (nx8260), .A0 (int_vec_buff_1), .A1 (nx1473), .B0 (
                      nx388), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_1 (.Q (int_vec_buff_1), .CK (wb_clk_i)
                        , .D (int_src_1), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_1)) ;
    INV_X0P5B_A12TS ix8265 (.Y (nx8264), .A (idat_cur_9)) ;
    AOI22_X0P5M_A12TS ix8269 (.Y (nx8268), .A0 (idat_cur_17), .A1 (nx1503), .B0 (
                      idat_cur_25), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8271 (.Y (nx8270), .A (rd), .B (nx1682)) ;
    OAI21_X0P5M_A12TS ix1797 (.Y (op3_n_2), .A0 (rd), .A1 (nx8273), .B0 (nx8285)
                      ) ;
    INV_X0P5B_A12TS ix8274 (.Y (nx8273), .A (op3_buff_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_2 (.Q (op3_buff_2), .CK (wb_clk_i), .D (
                        nx1784), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_2)
                        ) ;
    OAI211_X0P5M_A12TS ix1785 (.Y (nx1784), .A0 (nx7818), .A1 (nx7593), .B0 (
                       nx8277), .C0 (nx8283)) ;
    AOI22_X0P5M_A12TS ix8278 (.Y (nx8277), .A0 (int_vec_buff_2), .A1 (nx1473), .B0 (
                      nx1486), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_2 (.Q (int_vec_buff_2), .CK (wb_clk_i)
                        , .D (int_src_7), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_2)) ;
    AOI22_X0P5M_A12TS ix8284 (.Y (nx8283), .A0 (idat_cur_18), .A1 (nx1503), .B0 (
                      idat_cur_26), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8286 (.Y (nx8285), .A (rd), .B (nx1784)) ;
    OAI21_X0P5M_A12TS ix1865 (.Y (op3_n_3), .A0 (rd), .A1 (nx8288), .B0 (nx8300)
                      ) ;
    INV_X0P5B_A12TS ix8289 (.Y (nx8288), .A (op3_buff_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_3 (.Q (op3_buff_3), .CK (wb_clk_i), .D (
                        nx1852), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_3)
                        ) ;
    OAI211_X0P5M_A12TS ix1853 (.Y (nx1852), .A0 (nx7638), .A1 (nx7593), .B0 (
                       nx8292), .C0 (nx8298)) ;
    AOI22_X0P5M_A12TS ix8293 (.Y (nx8292), .A0 (int_vec_buff_3), .A1 (nx1473), .B0 (
                      nx120), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_3 (.Q (int_vec_buff_3), .CK (wb_clk_i)
                        , .D (int_src_3), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_3)) ;
    AOI22_X0P5M_A12TS ix8299 (.Y (nx8298), .A0 (idat_cur_19), .A1 (nx1503), .B0 (
                      idat_cur_27), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8301 (.Y (nx8300), .A (rd), .B (nx1852)) ;
    OAI21_X0P5M_A12TS ix1937 (.Y (op3_n_4), .A0 (rd), .A1 (nx8303), .B0 (nx8317)
                      ) ;
    INV_X0P5B_A12TS ix8304 (.Y (nx8303), .A (op3_buff_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_4 (.Q (op3_buff_4), .CK (wb_clk_i), .D (
                        nx1508), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_4)
                        ) ;
    OAI211_X0P5M_A12TS ix1292 (.Y (nx1508), .A0 (nx7788), .A1 (nx7593), .B0 (
                       nx8307), .C0 (nx8315)) ;
    AOI22_X0P5M_A12TS ix8308 (.Y (nx8307), .A0 (int_vec_buff_4), .A1 (nx1473), .B0 (
                      nx754), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_4 (.Q (int_vec_buff_4), .CK (wb_clk_i)
                        , .D (int_src_4), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_4)) ;
    INV_X0P5B_A12TS ix8312 (.Y (nx8311), .A (idat_cur_12)) ;
    AOI22_X0P5M_A12TS ix8316 (.Y (nx8315), .A0 (idat_cur_20), .A1 (nx1503), .B0 (
                      idat_cur_28), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8318 (.Y (nx8317), .A (rd), .B (nx1508)) ;
    OAI21_X0P5M_A12TS ix1294 (.Y (op3_n_5), .A0 (rd), .A1 (nx8320), .B0 (nx8332)
                      ) ;
    INV_X0P5B_A12TS ix8321 (.Y (nx8320), .A (op3_buff_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_5 (.Q (op3_buff_5), .CK (wb_clk_i), .D (
                        nx2088), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_5)
                        ) ;
    OAI211_X0P5M_A12TS ix2089 (.Y (nx2088), .A0 (nx7714), .A1 (nx7593), .B0 (
                       nx8324), .C0 (nx8330)) ;
    AOI22_X0P5M_A12TS ix8325 (.Y (nx8324), .A0 (int_vec_buff_5), .A1 (nx1473), .B0 (
                      nx1479), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_5 (.Q (int_vec_buff_5), .CK (wb_clk_i)
                        , .D (int_src_5), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_5)) ;
    AOI22_X0P5M_A12TS ix8331 (.Y (nx8330), .A0 (idat_cur_21), .A1 (nx1503), .B0 (
                      idat_cur_29), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8333 (.Y (nx8332), .A (rd), .B (nx2088)) ;
    OAI21_X0P5M_A12TS ix1295 (.Y (op3_n_6), .A0 (rd), .A1 (nx8335), .B0 (nx8347)
                      ) ;
    INV_X0P5B_A12TS ix8336 (.Y (nx8335), .A (op3_buff_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_6 (.Q (op3_buff_6), .CK (wb_clk_i), .D (
                        nx1516), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_6)
                        ) ;
    OAI211_X0P5M_A12TS ix1296 (.Y (nx1516), .A0 (nx7929), .A1 (nx7593), .B0 (
                       nx8339), .C0 (nx8345)) ;
    AOI22_X0P5M_A12TS ix8340 (.Y (nx8339), .A0 (int_vec_buff_6), .A1 (nx1473), .B0 (
                      nx822), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_6 (.Q (int_vec_buff_6), .CK (wb_clk_i)
                        , .D (int_src_7), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_6)) ;
    AOI22_X0P5M_A12TS ix8346 (.Y (nx8345), .A0 (idat_cur_22), .A1 (nx1503), .B0 (
                      idat_cur_30), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8348 (.Y (nx8347), .A (rd), .B (nx1516)) ;
    OAI21_X0P5M_A12TS ix2295 (.Y (op3_n_7), .A0 (rd), .A1 (nx8350), .B0 (nx8362)
                      ) ;
    INV_X0P5B_A12TS ix8351 (.Y (nx8350), .A (op3_buff_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_op3_buff_7 (.Q (op3_buff_7), .CK (wb_clk_i), .D (
                        nx2282), .R (wb_rst_i), .SE (NOT_rd), .SI (op3_buff_7)
                        ) ;
    OAI211_X0P5M_A12TS ix2283 (.Y (nx2282), .A0 (nx7984), .A1 (nx7593), .B0 (
                       nx8354), .C0 (nx8360)) ;
    AOI22_X0P5M_A12TS ix8355 (.Y (nx8354), .A0 (int_vec_buff_7), .A1 (nx1473), .B0 (
                      nx1108), .B1 (nx1476)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_buff_7 (.Q (int_vec_buff_7), .CK (wb_clk_i)
                        , .D (int_src_7), .R (wb_rst_i), .SE (NOT_intr), .SI (
                        int_vec_buff_7)) ;
    AOI22_X0P5M_A12TS ix8361 (.Y (nx8360), .A0 (idat_cur_23), .A1 (nx1503), .B0 (
                      idat_cur_31), .B1 (nx1420)) ;
    NAND2_X0P5A_A12TS ix8363 (.Y (nx8362), .A (rd), .B (nx2282)) ;
    OAI21_X0P5M_A12TS ix1441 (.Y (op2_n_0), .A0 (rd), .A1 (nx8365), .B0 (nx8378)
                      ) ;
    INV_X0P5B_A12TS ix8366 (.Y (nx8365), .A (op2_buff_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_0 (.Q (op2_buff_0), .CK (wb_clk_i), .D (
                        nx1428), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_0)
                        ) ;
    OAI211_X0P5M_A12TS ix1429 (.Y (nx1428), .A0 (nx7901), .A1 (nx8369), .B0 (
                       nx8371), .C0 (nx8374)) ;
    NAND2_X0P5A_A12TS ix8370 (.Y (nx8369), .A (nx7665), .B (nx138)) ;
    AOI22_X0P5M_A12TS ix8372 (.Y (nx8371), .A0 (idat_cur_16), .A1 (nx1420), .B0 (
                      idat_old_8), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8375 (.Y (nx8374), .A0 (idat_old_24), .A1 (nx1404), .B0 (
                       idat_cur_0), .B1 (nx1502), .C0 (idat_old_16), .C1 (nx5675
                       )) ;
    NOR2_X0P5A_A12TS ix1405 (.Y (nx1404), .A (op_pos_0), .B (nx7654)) ;
    NOR2_X0P5A_A12TS ix1297 (.Y (nx1502), .A (nx7591), .B (nx7654)) ;
    NAND2_X0P5A_A12TS ix8379 (.Y (nx8378), .A (rd), .B (nx1428)) ;
    OAI21_X0P5M_A12TS ix1298 (.Y (op2_n_1), .A0 (rd), .A1 (nx8381), .B0 (nx8389)
                      ) ;
    INV_X0P5B_A12TS ix8382 (.Y (nx8381), .A (op2_buff_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_1 (.Q (op2_buff_1), .CK (wb_clk_i), .D (
                        nx1734), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_1)
                        ) ;
    OAI211_X0P5M_A12TS ix1735 (.Y (nx1734), .A0 (nx8264), .A1 (nx8369), .B0 (
                       nx8385), .C0 (nx8387)) ;
    AOI22_X0P5M_A12TS ix8386 (.Y (nx8385), .A0 (idat_cur_17), .A1 (nx1420), .B0 (
                      idat_old_9), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8388 (.Y (nx8387), .A0 (idat_old_25), .A1 (nx1404), .B0 (
                       idat_cur_1), .B1 (nx1502), .C0 (idat_old_17), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8390 (.Y (nx8389), .A (rd), .B (nx1734)) ;
    OAI21_X0P5M_A12TS ix1299 (.Y (op2_n_2), .A0 (rd), .A1 (nx8392), .B0 (nx8400)
                      ) ;
    INV_X0P5B_A12TS ix8393 (.Y (nx8392), .A (op2_buff_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_2 (.Q (op2_buff_2), .CK (wb_clk_i), .D (
                        nx1506), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_2)
                        ) ;
    OAI211_X0P5M_A12TS ix1300 (.Y (nx1506), .A0 (nx7851), .A1 (nx8369), .B0 (
                       nx8396), .C0 (nx8398)) ;
    AOI22_X0P5M_A12TS ix8397 (.Y (nx8396), .A0 (idat_cur_18), .A1 (nx1420), .B0 (
                      idat_old_10), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8399 (.Y (nx8398), .A0 (idat_old_26), .A1 (nx1404), .B0 (
                       idat_cur_2), .B1 (nx1502), .C0 (idat_old_18), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8401 (.Y (nx8400), .A (rd), .B (nx1506)) ;
    OAI21_X0P5M_A12TS ix1551 (.Y (op2_n_3), .A0 (rd), .A1 (nx8403), .B0 (nx8411)
                      ) ;
    INV_X0P5B_A12TS ix8404 (.Y (nx8403), .A (op2_buff_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_3 (.Q (op2_buff_3), .CK (wb_clk_i), .D (
                        nx1538), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_3)
                        ) ;
    OAI211_X0P5M_A12TS ix1539 (.Y (nx1538), .A0 (nx7668), .A1 (nx8369), .B0 (
                       nx8407), .C0 (nx8409)) ;
    AOI22_X0P5M_A12TS ix8408 (.Y (nx8407), .A0 (idat_cur_19), .A1 (nx1420), .B0 (
                      idat_old_11), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8410 (.Y (nx8409), .A0 (idat_old_27), .A1 (nx1404), .B0 (
                       idat_cur_3), .B1 (nx1502), .C0 (idat_old_19), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8412 (.Y (nx8411), .A (rd), .B (nx1538)) ;
    OAI21_X0P5M_A12TS ix1302 (.Y (op2_n_4), .A0 (rd), .A1 (nx8414), .B0 (nx8422)
                      ) ;
    INV_X0P5B_A12TS ix8415 (.Y (nx8414), .A (op2_buff_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_4 (.Q (op2_buff_4), .CK (wb_clk_i), .D (
                        nx1512), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_4)
                        ) ;
    OAI211_X0P5M_A12TS ix1304 (.Y (nx1512), .A0 (nx8311), .A1 (nx8369), .B0 (
                       nx8418), .C0 (nx8420)) ;
    AOI22_X0P5M_A12TS ix8419 (.Y (nx8418), .A0 (idat_cur_20), .A1 (nx1420), .B0 (
                      idat_old_12), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8421 (.Y (nx8420), .A0 (idat_old_28), .A1 (nx1404), .B0 (
                       idat_cur_4), .B1 (nx1502), .C0 (idat_old_20), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8423 (.Y (nx8422), .A (rd), .B (nx1512)) ;
    OAI21_X0P5M_A12TS ix1306 (.Y (op2_n_5), .A0 (rd), .A1 (nx8425), .B0 (nx8433)
                      ) ;
    INV_X0P5B_A12TS ix8426 (.Y (nx8425), .A (op2_buff_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_5 (.Q (op2_buff_5), .CK (wb_clk_i), .D (
                        nx1514), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_5)
                        ) ;
    OAI211_X0P5M_A12TS ix1308 (.Y (nx1514), .A0 (nx7747), .A1 (nx8369), .B0 (
                       nx8429), .C0 (nx8431)) ;
    AOI22_X0P5M_A12TS ix8430 (.Y (nx8429), .A0 (idat_cur_21), .A1 (nx1420), .B0 (
                      idat_old_13), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8432 (.Y (nx8431), .A0 (idat_old_29), .A1 (nx1404), .B0 (
                       idat_cur_5), .B1 (nx1502), .C0 (idat_old_21), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8434 (.Y (nx8433), .A (rd), .B (nx1514)) ;
    OAI21_X0P5M_A12TS ix1309 (.Y (op2_n_6), .A0 (rd), .A1 (nx8436), .B0 (nx8444)
                      ) ;
    INV_X0P5B_A12TS ix8437 (.Y (nx8436), .A (op2_buff_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_6 (.Q (op2_buff_6), .CK (wb_clk_i), .D (
                        nx1515), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_6)
                        ) ;
    OAI211_X0P5M_A12TS ix1310 (.Y (nx1515), .A0 (nx7953), .A1 (nx8369), .B0 (
                       nx8440), .C0 (nx8442)) ;
    AOI22_X0P5M_A12TS ix8441 (.Y (nx8440), .A0 (idat_cur_22), .A1 (nx1420), .B0 (
                      idat_old_14), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8443 (.Y (nx8442), .A0 (idat_old_30), .A1 (nx1404), .B0 (
                       idat_cur_6), .B1 (nx1502), .C0 (idat_old_22), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8445 (.Y (nx8444), .A (rd), .B (nx1515)) ;
    OAI21_X0P5M_A12TS ix2245 (.Y (op2_n_7), .A0 (rd), .A1 (nx8447), .B0 (nx8455)
                      ) ;
    INV_X0P5B_A12TS ix8448 (.Y (nx8447), .A (op2_buff_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_op2_buff_7 (.Q (op2_buff_7), .CK (wb_clk_i), .D (
                        nx2232), .R (wb_rst_i), .SE (NOT_rd), .SI (op2_buff_7)
                        ) ;
    OAI211_X0P5M_A12TS ix2233 (.Y (nx2232), .A0 (nx8010), .A1 (nx8369), .B0 (
                       nx8451), .C0 (nx8453)) ;
    AOI22_X0P5M_A12TS ix8452 (.Y (nx8451), .A0 (idat_cur_23), .A1 (nx1420), .B0 (
                      idat_old_15), .B1 (nx1475)) ;
    AOI222_X0P5M_A12TS ix8454 (.Y (nx8453), .A0 (idat_old_31), .A1 (nx1404), .B0 (
                       idat_cur_7), .B1 (nx1502), .C0 (idat_old_23), .C1 (nx5675
                       )) ;
    NAND2_X0P5A_A12TS ix8456 (.Y (nx8455), .A (rd), .B (nx2232)) ;
    OAI21_X0P5M_A12TS ix4201 (.Y (wbi_adr_o[0]), .A0 (istb_t), .A1 (nx8458), .B0 (
                      nx8494)) ;
    INV_X0P5B_A12TS ix8459 (.Y (nx8458), .A (pc_buf_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_0 (.Q (pc_buf_0), .CK (wb_clk_i), .D (nx2488)
                        , .R (wb_rst_i), .SE (NOT_nx2430), .SI (pc_buf_0)) ;
    NAND3_X0P5A_A12TS ix2489 (.Y (nx2488), .A (nx8462), .B (nx8466), .C (nx8474)
                      ) ;
    AOI22_X0P5M_A12TS ix8463 (.Y (nx8462), .A0 (nx7537), .A1 (pc_buf_0), .B0 (
                      nx2438), .B1 (nx2478)) ;
    NOR3_X0P5A_A12TS ix2479 (.Y (nx2478), .A (nx7533), .B (nx7537), .C (
                     pc_wr_sel_1)) ;
    AO21A1AI2_X0P5M_A12TS ix8467 (.Y (nx8466), .A0 (nx8468), .A1 (nx2464), .B0 (
                          nx2454), .C0 (des_acc_0)) ;
    INV_X0P5B_A12TS ix8469 (.Y (nx8468), .A (pc_wr_sel_0)) ;
    NOR3_X0P5A_A12TS ix2465 (.Y (nx2464), .A (pc_wr_sel_2), .B (nx7537), .C (
                     pc_wr_sel_1)) ;
    NOR2_X0P5A_A12TS ix2455 (.Y (nx2454), .A (nx7533), .B (nx8472)) ;
    NAND2_X0P5A_A12TS ix8473 (.Y (nx8472), .A (pc_wr_sel_1), .B (pc_wr_dup_1371)
                      ) ;
    OAI211_X0P5M_A12TS ix8475 (.Y (nx8474), .A0 (nx2438), .A1 (pc_0), .B0 (
                       nx8489), .C0 (nx2446)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_0 (.Q (pc_0), .CK (wb_clk_i), .D (nx6794), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8479 (.Y (nx8478), .A0 (pc_buf_0), .A1 (pc_wr_r2), .B0 (
                          nx2512), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix1311 (.Y (nx2512), .A0 (nx8481), .A1 (nx7905), .B0 (
                       pc_wr_r2), .C0 (nx2504)) ;
    OAI21_X0P5M_A12TS ix8482 (.Y (nx8481), .A0 (pc_buf_0), .A1 (op_pos_0), .B0 (
                      nx8483)) ;
    NAND2_X0P5A_A12TS ix8484 (.Y (nx8483), .A (op_pos_0), .B (pc_buf_0)) ;
    NOR2_X0P5A_A12TS ix2505 (.Y (nx2504), .A (nx7905), .B (nx8481)) ;
    OAI21_X0P5M_A12TS ix1312 (.Y (nx1518), .A0 (NOT_rd), .A1 (int_ack_t), .B0 (
                      nx7603)) ;
    NAND2_X0P5A_A12TS ix8490 (.Y (nx8489), .A (pc_0), .B (nx2438)) ;
    NOR2_X0P5A_A12TS ix2447 (.Y (nx2446), .A (pc_wr_sel_2), .B (nx8472)) ;
    NAND2_X0P5A_A12TS ix8495 (.Y (nx8494), .A (istb_t), .B (iadr_t_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_0 (.Q (iadr_t_0), .CK (wb_clk_i), .D (
                        des_acc_0), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_0)) ;
    OAI21_X0P5M_A12TS ix1314 (.Y (wbi_adr_o[1]), .A0 (istb_t), .A1 (nx8498), .B0 (
                      nx8533)) ;
    INV_X0P5B_A12TS ix8499 (.Y (nx8498), .A (pc_buf_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_1 (.Q (pc_buf_1), .CK (wb_clk_i), .D (nx2572)
                        , .R (wb_rst_i), .SE (NOT_nx2430), .SI (pc_buf_1)) ;
    OAI221_X0P5M_A12TS ix2573 (.Y (nx2572), .A0 (nx8502), .A1 (nx8504), .B0 (
                       nx8506), .B1 (nx8523), .C0 (nx8525)) ;
    MXIT2_X0P5M_A12TS ix8503 (.Y (nx8502), .A (op2_n_1), .B (op3_n_1), .S0 (
                      pc_wr_sel_0)) ;
    XNOR2_X0P5M_A12TS ix8507 (.Y (nx8506), .A (nx8489), .B (nx8508)) ;
    XOR2_X0P5M_A12TS ix8509 (.Y (nx8508), .A (pc_1), .B (nx8502)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_1 (.Q (pc_1), .CK (wb_clk_i), .D (nx6814), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8513 (.Y (nx8512), .A0 (pc_buf_1), .A1 (pc_wr_r2), .B0 (
                          nx2588), .C0 (nx1518)) ;
    NOR2_X0P5A_A12TS ix2589 (.Y (nx2588), .A (pc_wr_r2), .B (nx8515)) ;
    XOR2_X0P5M_A12TS ix8516 (.Y (nx8515), .A (nx2504), .B (nx8517)) ;
    XNOR2_X0P5M_A12TS ix8518 (.Y (nx8517), .A (nx7613), .B (nx8519)) ;
    XNOR2_X0P5M_A12TS ix8520 (.Y (nx8519), .A (nx8483), .B (nx8521)) ;
    XNOR2_X0P5M_A12TS ix8522 (.Y (nx8521), .A (op_pos_1), .B (pc_buf_1)) ;
    NAND3_X0P5A_A12TS ix8524 (.Y (nx8523), .A (pc_wr_dup_1371), .B (pc_wr_sel_1)
                      , .C (nx7533)) ;
    AOI22_X0P5M_A12TS ix8526 (.Y (nx8525), .A0 (nx7537), .A1 (pc_buf_1), .B0 (
                      des_acc_1), .B1 (nx2562)) ;
    NAND3_X0P5A_A12TS ix8529 (.Y (nx8528), .A (pc_wr_dup_1371), .B (pc_wr_sel_1)
                      , .C (pc_wr_sel_2)) ;
    NOR3_X0P5A_A12TS ix8532 (.Y (NOT_nx2552), .A (nx7537), .B (pc_wr_sel_1), .C (
                     pc_wr_sel_0)) ;
    NAND2_X0P5A_A12TS ix8534 (.Y (nx8533), .A (istb_t), .B (iadr_t_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_1 (.Q (iadr_t_1), .CK (wb_clk_i), .D (
                        des_acc_1), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_1)) ;
    OAI21_X0P5M_A12TS ix4225 (.Y (wbi_adr_o[2]), .A0 (istb_t), .A1 (nx8537), .B0 (
                      nx8585)) ;
    XNOR2_X0P5M_A12TS ix8538 (.Y (nx8537), .A (pc_buf_2), .B (nx5672)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_buf_2 (.Q (pc_buf_2), .CK (wb_clk_i), .D (nx6824)
                       , .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6825 (.Y (nx6824), .A0 (nx8541), .A1 (nx2430), .B0 (
                      nx8546)) ;
    INV_X0P5B_A12TS ix8542 (.Y (nx8541), .A (pc_buf_2)) ;
    NAND2_X0P5A_A12TS ix2431 (.Y (nx2430), .A (nx8544), .B (pc_wr_dup_1371)) ;
    OAI31_X0P5M_A12TS ix8545 (.Y (nx8544), .A0 (nx8468), .A1 (pc_wr_sel_2), .A2 (
                      pc_wr_sel_1), .B0 (pc_wr_dup_1371)) ;
    OAI21_X0P5M_A12TS ix8547 (.Y (nx8546), .A0 (nx2648), .A1 (nx2638), .B0 (
                      nx2430)) ;
    OAI22_X0P5M_A12TS ix2649 (.Y (nx2648), .A0 (nx8549), .A1 (nx8551), .B0 (
                      pc_wr_dup_1371), .B1 (nx8537)) ;
    INV_X0P5B_A12TS ix8550 (.Y (nx8549), .A (des_acc_2)) ;
    OAI22_X0P5M_A12TS ix2639 (.Y (nx2638), .A0 (nx8560), .A1 (nx8504), .B0 (
                      nx8562), .B1 (nx8523)) ;
    MXIT2_X0P5M_A12TS ix8561 (.Y (nx8560), .A (op2_n_2), .B (op3_n_2), .S0 (
                      pc_wr_sel_0)) ;
    XNOR2_X0P5M_A12TS ix8563 (.Y (nx8562), .A (nx8564), .B (nx8570)) ;
    MXIT2_X0P5M_A12TS ix8568 (.Y (nx8567), .A (op2_n_0), .B (op3_n_0), .S0 (
                      pc_wr_sel_0)) ;
    XOR2_X0P5M_A12TS ix8571 (.Y (nx8570), .A (pc_2), .B (nx8560)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_2 (.Q (pc_2), .CK (wb_clk_i), .D (nx2674), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_2)) ;
    OAI211_X0P5M_A12TS ix8575 (.Y (nx8574), .A0 (nx2658), .A1 (nx2604), .B0 (
                       nx7603), .C0 (nx8583)) ;
    CGENI_X1M_A12TS ix2613 (.CON (nx2612), .A (nx8483), .B (nx7595), .CI (nx8498
                    )) ;
    XNOR2_X0P5M_A12TS ix8579 (.Y (nx8578), .A (op_pos_2), .B (pc_buf_2)) ;
    MXIT2_X0P5M_A12TS ix2605 (.Y (nx2604), .A (nx8581), .B (nx8519), .S0 (nx8517
                      )) ;
    NAND2_X0P5A_A12TS ix8584 (.Y (nx8583), .A (nx2604), .B (nx2658)) ;
    NAND2_X0P5A_A12TS ix8586 (.Y (nx8585), .A (istb_t), .B (iadr_t_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_2 (.Q (iadr_t_2), .CK (wb_clk_i), .D (
                        des_acc_2), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_3 (.Q (iadr_t_3), .CK (wb_clk_i), .D (
                        des_acc_3), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_3)) ;
    NAND2_X0P5A_A12TS ix8593 (.Y (nx8592), .A (nx7555), .B (nx2722)) ;
    OAI21_X0P5M_A12TS ix2723 (.Y (nx2722), .A0 (nx8595), .A1 (nx5672), .B0 (
                      nx8626)) ;
    INV_X0P5B_A12TS ix8596 (.Y (nx8595), .A (pc_buf_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_3 (.Q (pc_buf_3), .CK (wb_clk_i), .D (nx2730)
                        , .R (wb_rst_i), .SE (NOT_nx2430), .SI (pc_buf_3)) ;
    OAI221_X0P5M_A12TS ix2731 (.Y (nx2730), .A0 (nx8599), .A1 (nx8504), .B0 (
                       nx8601), .B1 (nx8523), .C0 (nx8624)) ;
    MXIT2_X0P5M_A12TS ix8600 (.Y (nx8599), .A (op2_n_3), .B (op3_n_3), .S0 (
                      pc_wr_sel_0)) ;
    XOR2_X0P5M_A12TS ix8602 (.Y (nx8601), .A (nx2696), .B (nx8606)) ;
    CGENI_X1M_A12TS ix2697 (.CON (nx2696), .A (nx8564), .B (nx8604), .CI (nx8560
                    )) ;
    INV_X0P5B_A12TS ix8605 (.Y (nx8604), .A (pc_2)) ;
    XOR2_X0P5M_A12TS ix8607 (.Y (nx8606), .A (pc_3), .B (nx8599)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_3 (.Q (pc_3), .CK (wb_clk_i), .D (nx2770), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_3)) ;
    OAI211_X0P5M_A12TS ix8611 (.Y (nx8610), .A0 (nx2754), .A1 (nx2662), .B0 (
                       nx7603), .C0 (nx8622)) ;
    AOI21_X0P5M_A12TS ix2755 (.Y (nx2754), .A0 (nx8613), .A1 (pc_buf_3), .B0 (
                      nx2746)) ;
    CGENI_X1M_A12TS ix8614 (.CON (nx8613), .A (nx2612), .B (op_pos_2), .CI (
                    pc_buf_2)) ;
    NOR2_X0P5A_A12TS ix2747 (.Y (nx2746), .A (pc_buf_3), .B (nx8613)) ;
    XOR2_X0P5M_A12TS ix8621 (.Y (nx8620), .A (nx2612), .B (nx8578)) ;
    NAND2_X0P5A_A12TS ix8623 (.Y (nx8622), .A (nx2662), .B (nx2754)) ;
    AOI22_X0P5M_A12TS ix8625 (.Y (nx8624), .A0 (des_acc_3), .A1 (nx2562), .B0 (
                      nx7537), .B1 (nx2722)) ;
    OAI211_X0P5M_A12TS ix8627 (.Y (nx8626), .A0 (pc_buf_2), .A1 (pc_buf_3), .B0 (
                       nx5672), .C0 (nx8628)) ;
    NAND2_X0P5A_A12TS ix8629 (.Y (nx8628), .A (pc_buf_3), .B (pc_buf_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_4 (.Q (iadr_t_4), .CK (wb_clk_i), .D (
                        des_acc_4), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_4)) ;
    NAND2_X0P5A_A12TS ix8635 (.Y (nx8634), .A (nx7555), .B (nx2818)) ;
    OAI21_X0P5M_A12TS ix2819 (.Y (nx2818), .A0 (nx8637), .A1 (nx5672), .B0 (
                      nx8666)) ;
    INV_X0P5B_A12TS ix8638 (.Y (nx8637), .A (pc_buf_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_4 (.Q (pc_buf_4), .CK (wb_clk_i), .D (nx2826)
                        , .R (wb_rst_i), .SE (NOT_nx2430), .SI (pc_buf_4)) ;
    OAI221_X0P5M_A12TS ix2827 (.Y (nx2826), .A0 (nx8641), .A1 (nx8504), .B0 (
                       nx8643), .B1 (nx8523), .C0 (nx8664)) ;
    MXIT2_X0P5M_A12TS ix8642 (.Y (nx8641), .A (op2_n_4), .B (op3_n_4), .S0 (
                      pc_wr_sel_0)) ;
    XNOR2_X0P5M_A12TS ix8644 (.Y (nx8643), .A (nx8645), .B (nx8648)) ;
    CGENI_X1M_A12TS ix8646 (.CON (nx8645), .A (nx2696), .B (pc_3), .CI (nx2686)
                    ) ;
    XOR2_X0P5M_A12TS ix8649 (.Y (nx8648), .A (pc_4), .B (nx8641)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_4 (.Q (pc_4), .CK (wb_clk_i), .D (nx6874), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8653 (.Y (nx8652), .A0 (pc_buf_4), .A1 (pc_wr_r2), .B0 (
                          nx2858), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix2859 (.Y (nx2858), .A0 (nx8655), .A1 (nx8622), .B0 (
                       pc_wr_r2), .C0 (nx2850)) ;
    OAI21_X0P5M_A12TS ix8656 (.Y (nx8655), .A0 (nx2838), .A1 (nx2746), .B0 (
                      nx8659)) ;
    AO21A1AI2_X0P5M_A12TS ix8660 (.Y (nx8659), .A0 (pc_buf_4), .A1 (pc_buf_3), .B0 (
                          nx8661), .C0 (nx2746)) ;
    NOR2_X0P5A_A12TS ix8662 (.Y (nx8661), .A (pc_buf_3), .B (pc_buf_4)) ;
    NOR2_X0P5A_A12TS ix2851 (.Y (nx2850), .A (nx8622), .B (nx8655)) ;
    AOI22_X0P5M_A12TS ix8665 (.Y (nx8664), .A0 (des_acc_4), .A1 (nx2562), .B0 (
                      nx7537), .B1 (nx2818)) ;
    OAI211_X0P5M_A12TS ix8667 (.Y (nx8666), .A0 (nx2710), .A1 (pc_buf_4), .B0 (
                       nx5672), .C0 (nx8669)) ;
    NAND3_X0P5A_A12TS ix8670 (.Y (nx8669), .A (pc_buf_4), .B (pc_buf_3), .C (
                      pc_buf_2)) ;
    OAI21_X0P5M_A12TS ix4261 (.Y (wbi_adr_o[5]), .A0 (istb_t), .A1 (nx8672), .B0 (
                      nx8710)) ;
    AOI21_X0P5M_A12TS ix8673 (.Y (nx8672), .A0 (pc_buf_5), .A1 (nx8705), .B0 (
                      nx2904)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_buf_5 (.Q (pc_buf_5), .CK (wb_clk_i), .D (nx6884)
                       , .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6885 (.Y (nx6884), .A0 (nx8676), .A1 (nx2430), .B0 (
                      nx8678)) ;
    INV_X0P5B_A12TS ix8677 (.Y (nx8676), .A (pc_buf_5)) ;
    OAI21_X0P5M_A12TS ix8679 (.Y (nx8678), .A0 (nx2916), .A1 (nx2892), .B0 (
                      nx2430)) ;
    OAI22_X0P5M_A12TS ix2917 (.Y (nx2916), .A0 (nx8681), .A1 (nx8551), .B0 (
                      pc_wr_dup_1371), .B1 (nx8672)) ;
    INV_X0P5B_A12TS ix8682 (.Y (nx8681), .A (des_acc_5)) ;
    OAI22_X0P5M_A12TS ix2893 (.Y (nx2892), .A0 (nx8684), .A1 (nx8504), .B0 (
                      nx8686), .B1 (nx8523)) ;
    MXIT2_X0P5M_A12TS ix8685 (.Y (nx8684), .A (op2_n_5), .B (op3_n_5), .S0 (
                      pc_wr_sel_0)) ;
    XOR2_X0P5M_A12TS ix8687 (.Y (nx8686), .A (nx2884), .B (nx8691)) ;
    CGENI_X1M_A12TS ix2885 (.CON (nx2884), .A (nx8645), .B (nx8689), .CI (nx8641
                    )) ;
    INV_X0P5B_A12TS ix8690 (.Y (nx8689), .A (pc_4)) ;
    XOR2_X0P5M_A12TS ix8692 (.Y (nx8691), .A (pc_5), .B (nx8684)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_5 (.Q (pc_5), .CK (wb_clk_i), .D (nx2954), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_5)) ;
    OAI211_X0P5M_A12TS ix8696 (.Y (nx8695), .A0 (nx2938), .A1 (nx2850), .B0 (
                       nx7603), .C0 (nx8703)) ;
    AOI21_X0P5M_A12TS ix2939 (.Y (nx2938), .A0 (nx8698), .A1 (nx8659), .B0 (
                      nx2932)) ;
    OA21A1OI2_X0P5M_A12TS ix8699 (.Y (nx8698), .A0 (pc_buf_3), .A1 (pc_buf_4), .B0 (
                          pc_buf_5), .C0 (nx8700)) ;
    NOR3_X0P5A_A12TS ix8701 (.Y (nx8700), .A (pc_buf_3), .B (pc_buf_4), .C (
                     pc_buf_5)) ;
    NOR2_X0P5A_A12TS ix2933 (.Y (nx2932), .A (nx8659), .B (nx8698)) ;
    NAND2_X0P5A_A12TS ix8704 (.Y (nx8703), .A (nx2850), .B (nx2938)) ;
    AOI211_X0P5M_A12TS ix2905 (.Y (nx2904), .A0 (nx8669), .A1 (nx8676), .B0 (
                       nx8705), .C0 (nx2898)) ;
    NOR2_X0P5A_A12TS ix2899 (.Y (nx2898), .A (nx8676), .B (nx8669)) ;
    NAND2_X0P5A_A12TS ix8711 (.Y (nx8710), .A (istb_t), .B (iadr_t_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_5 (.Q (iadr_t_5), .CK (wb_clk_i), .D (
                        des_acc_5), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_6 (.Q (iadr_t_6), .CK (wb_clk_i), .D (
                        des_acc_6), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_6)) ;
    NAND2_X0P5A_A12TS ix8718 (.Y (nx8717), .A (nx7555), .B (nx3002)) ;
    OAI21_X0P5M_A12TS ix3003 (.Y (nx3002), .A0 (nx8720), .A1 (nx5672), .B0 (
                      nx8747)) ;
    INV_X0P5B_A12TS ix8721 (.Y (nx8720), .A (pc_buf_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_6 (.Q (pc_buf_6), .CK (wb_clk_i), .D (nx3010)
                        , .R (wb_rst_i), .SE (NOT_nx2430), .SI (pc_buf_6)) ;
    OAI221_X0P5M_A12TS ix3011 (.Y (nx3010), .A0 (nx8724), .A1 (nx8504), .B0 (
                       nx8726), .B1 (nx8523), .C0 (nx8745)) ;
    MXIT2_X0P5M_A12TS ix8725 (.Y (nx8724), .A (op2_n_6), .B (op3_n_6), .S0 (
                      pc_wr_sel_0)) ;
    XNOR2_X0P5M_A12TS ix8727 (.Y (nx8726), .A (nx8728), .B (nx8731)) ;
    CGENI_X1M_A12TS ix8729 (.CON (nx8728), .A (nx2884), .B (pc_5), .CI (nx2874)
                    ) ;
    XOR2_X0P5M_A12TS ix8732 (.Y (nx8731), .A (pc_6), .B (nx8724)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_6 (.Q (pc_6), .CK (wb_clk_i), .D (nx6914), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8736 (.Y (nx8735), .A0 (pc_buf_6), .A1 (pc_wr_r2), .B0 (
                          nx3042), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix3043 (.Y (nx3042), .A0 (nx8738), .A1 (nx8703), .B0 (
                       pc_wr_r2), .C0 (nx3034)) ;
    OAI21_X0P5M_A12TS ix8739 (.Y (nx8738), .A0 (nx3022), .A1 (nx2932), .B0 (
                      nx8742)) ;
    OAI21_X0P5M_A12TS ix3023 (.Y (nx3022), .A0 (nx8720), .A1 (nx8700), .B0 (
                      nx3016)) ;
    NAND2_X0P5A_A12TS ix3017 (.Y (nx3016), .A (nx8700), .B (nx8720)) ;
    NAND2_X0P5A_A12TS ix8743 (.Y (nx8742), .A (nx2932), .B (nx3022)) ;
    NOR2_X0P5A_A12TS ix3035 (.Y (nx3034), .A (nx8703), .B (nx8738)) ;
    AOI22_X0P5M_A12TS ix8746 (.Y (nx8745), .A0 (des_acc_6), .A1 (nx2562), .B0 (
                      nx7537), .B1 (nx3002)) ;
    OAI211_X0P5M_A12TS ix8748 (.Y (nx8747), .A0 (nx2898), .A1 (pc_buf_6), .B0 (
                       nx5672), .C0 (nx8749)) ;
    NAND2_X0P5A_A12TS ix8750 (.Y (nx8749), .A (pc_buf_6), .B (nx2898)) ;
    OAI21_X0P5M_A12TS ix4285 (.Y (wbi_adr_o[7]), .A0 (istb_t), .A1 (nx8752), .B0 (
                      nx8787)) ;
    AOI21_X0P5M_A12TS ix8753 (.Y (nx8752), .A0 (pc_buf_7), .A1 (nx8705), .B0 (
                      nx3088)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_buf_7 (.Q (pc_buf_7), .CK (wb_clk_i), .D (nx6924)
                       , .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix6925 (.Y (nx6924), .A0 (nx8756), .A1 (nx2430), .B0 (
                      nx8758)) ;
    INV_X0P5B_A12TS ix8757 (.Y (nx8756), .A (pc_buf_7)) ;
    OAI21_X0P5M_A12TS ix8759 (.Y (nx8758), .A0 (nx3100), .A1 (nx3076), .B0 (
                      nx2430)) ;
    OAI22_X0P5M_A12TS ix3101 (.Y (nx3100), .A0 (nx8761), .A1 (nx8551), .B0 (
                      pc_wr_dup_1371), .B1 (nx8752)) ;
    INV_X0P5B_A12TS ix8762 (.Y (nx8761), .A (des_acc_7)) ;
    OAI22_X0P5M_A12TS ix3077 (.Y (nx3076), .A0 (nx8764), .A1 (nx8504), .B0 (
                      nx8766), .B1 (nx8523)) ;
    MXIT2_X0P5M_A12TS ix8765 (.Y (nx8764), .A (op2_n_7), .B (op3_n_7), .S0 (
                      pc_wr_sel_0)) ;
    XOR2_X0P5M_A12TS ix8767 (.Y (nx8766), .A (nx3068), .B (nx8771)) ;
    CGENI_X1M_A12TS ix3069 (.CON (nx3068), .A (nx8728), .B (nx8769), .CI (nx8724
                    )) ;
    INV_X0P5B_A12TS ix8770 (.Y (nx8769), .A (pc_6)) ;
    XOR2_X0P5M_A12TS ix8772 (.Y (nx8771), .A (pc_7), .B (nx8764)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_7 (.Q (pc_7), .CK (wb_clk_i), .D (nx3138), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_7)) ;
    OAI211_X0P5M_A12TS ix8776 (.Y (nx8775), .A0 (nx3122), .A1 (nx3034), .B0 (
                       nx7603), .C0 (nx8783)) ;
    AOI21_X0P5M_A12TS ix3123 (.Y (nx3122), .A0 (nx8778), .A1 (nx8742), .B0 (
                      nx3116)) ;
    AOI21_X0P5M_A12TS ix8779 (.Y (nx8778), .A0 (pc_buf_7), .A1 (nx3016), .B0 (
                      nx8780)) ;
    NOR2_X0P5A_A12TS ix8781 (.Y (nx8780), .A (nx3016), .B (pc_buf_7)) ;
    NOR2_X0P5A_A12TS ix3117 (.Y (nx3116), .A (nx8742), .B (nx8778)) ;
    NAND2_X0P5A_A12TS ix8784 (.Y (nx8783), .A (nx3034), .B (nx3122)) ;
    AOI211_X0P5M_A12TS ix3089 (.Y (nx3088), .A0 (nx8749), .A1 (nx8756), .B0 (
                       nx8705), .C0 (nx3082)) ;
    NOR2_X0P5A_A12TS ix3083 (.Y (nx3082), .A (nx8756), .B (nx8749)) ;
    NAND2_X0P5A_A12TS ix8788 (.Y (nx8787), .A (istb_t), .B (iadr_t_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_7 (.Q (iadr_t_7), .CK (wb_clk_i), .D (
                        des_acc_7), .R (wb_rst_i), .SE (NOT_nx226), .SI (
                        iadr_t_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_8 (.Q (iadr_t_8), .CK (wb_clk_i), .D (des2_0)
                        , .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_8)) ;
    NAND2_X0P5A_A12TS ix8795 (.Y (nx8794), .A (nx7555), .B (nx3206)) ;
    OAI21_X0P5M_A12TS ix3207 (.Y (nx3206), .A0 (nx8797), .A1 (nx5672), .B0 (
                      nx8830)) ;
    INV_X0P5B_A12TS ix8798 (.Y (nx8797), .A (pc_buf_8)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_8 (.Q (pc_buf_8), .CK (wb_clk_i), .D (nx3222)
                        , .R (wb_rst_i), .SE (NOT_nx2554), .SI (pc_buf_8)) ;
    NAND3_X0P5A_A12TS ix3223 (.Y (nx3222), .A (nx8801), .B (nx8803), .C (nx8806)
                      ) ;
    AOI222_X0P5M_A12TS ix8802 (.Y (nx8801), .A0 (des_acc_0), .A1 (NOT_nx2430), .B0 (
                       des2_0), .B1 (nx2558), .C0 (nx7537), .C1 (nx3206)) ;
    AOI32_X0P5M_A12TS ix8804 (.Y (nx8803), .A0 (op1_n_5), .A1 (pc_wr_sel_2), .A2 (
                      NOT_nx2552), .B0 (op2_n_0), .B1 (nx3184)) ;
    NOR3_X0P5A_A12TS ix3185 (.Y (nx3184), .A (nx8544), .B (pc_wr_sel_1), .C (
                     NOT_nx2552)) ;
    MXIT2_X0P5M_A12TS ix8807 (.Y (nx8806), .A (nx3168), .B (nx3146), .S0 (nx8811
                      )) ;
    NOR2_X0P5A_A12TS ix3169 (.Y (nx3168), .A (nx8764), .B (nx8523)) ;
    NOR2_X0P5A_A12TS ix3147 (.Y (nx3146), .A (nx3058), .B (nx8523)) ;
    NOR2_X0P5A_A12TS ix8812 (.Y (nx8811), .A (nx8813), .B (nx3156)) ;
    NOR2B_X0P7M_A12TS ix8814 (.Y (nx8813), .AN (nx8815), .B (pc_8)) ;
    CGENI_X1M_A12TS ix8816 (.CON (nx8815), .A (nx3068), .B (pc_7), .CI (nx3058)
                    ) ;
    DFFRPQ_X0P5M_A12TS reg_pc_8 (.Q (pc_8), .CK (wb_clk_i), .D (nx6954), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8820 (.Y (nx8819), .A0 (pc_buf_8), .A1 (pc_wr_r2), .B0 (
                          nx3254), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix3255 (.Y (nx3254), .A0 (nx8822), .A1 (nx8783), .B0 (
                       pc_wr_r2), .C0 (nx3246)) ;
    OAI21_X0P5M_A12TS ix8823 (.Y (nx8822), .A0 (nx3234), .A1 (nx3116), .B0 (
                      nx8826)) ;
    OAI21_X0P5M_A12TS ix3235 (.Y (nx3234), .A0 (nx8797), .A1 (nx8780), .B0 (
                      nx3228)) ;
    NAND2_X0P5A_A12TS ix3229 (.Y (nx3228), .A (nx8780), .B (nx8797)) ;
    NAND2_X0P5A_A12TS ix8827 (.Y (nx8826), .A (nx3116), .B (nx3234)) ;
    NOR2_X0P5A_A12TS ix3247 (.Y (nx3246), .A (nx8783), .B (nx8822)) ;
    OAI211_X0P5M_A12TS ix8831 (.Y (nx8830), .A0 (nx3082), .A1 (pc_buf_8), .B0 (
                       nx5672), .C0 (nx8832)) ;
    NAND2_X0P5A_A12TS ix8833 (.Y (nx8832), .A (pc_buf_8), .B (nx3082)) ;
    OAI21_X0P5M_A12TS ix1315 (.Y (wbi_adr_o[9]), .A0 (istb_t), .A1 (nx8835), .B0 (
                      nx8879)) ;
    AOI21_X0P5M_A12TS ix8836 (.Y (nx8835), .A0 (pc_buf_9), .A1 (nx8705), .B0 (
                      nx3302)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_9 (.Q (pc_buf_9), .CK (wb_clk_i), .D (nx3324)
                        , .R (wb_rst_i), .SE (NOT_nx2554), .SI (pc_buf_9)) ;
    NAND4_X0P5A_A12TS ix3325 (.Y (nx3324), .A (nx8839), .B (nx8854), .C (nx8856)
                      , .D (nx8873)) ;
    AOI222_X0P5M_A12TS ix8840 (.Y (nx8839), .A0 (des_acc_1), .A1 (NOT_nx2430), .B0 (
                       des2_1), .B1 (nx2558), .C0 (nx7537), .C1 (nx3308)) ;
    INV_X0P5B_A12TS ix8843 (.Y (nx8842), .A (pc_buf_9)) ;
    AOI32_X0P5M_A12TS ix8855 (.Y (nx8854), .A0 (op1_n_6), .A1 (pc_wr_sel_2), .A2 (
                      NOT_nx2552), .B0 (op2_n_1), .B1 (nx3184)) ;
    AO21A1AI2_X0P5M_A12TS ix8857 (.Y (nx8856), .A0 (pc_9), .A1 (nx3158), .B0 (
                          nx8871), .C0 (nx3168)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_9 (.Q (pc_9), .CK (wb_clk_i), .D (nx3360), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_9)) ;
    OAI211_X0P5M_A12TS ix8861 (.Y (nx8860), .A0 (nx3344), .A1 (nx3246), .B0 (
                       nx7603), .C0 (nx8868)) ;
    AOI21_X0P5M_A12TS ix3345 (.Y (nx3344), .A0 (nx8863), .A1 (nx8826), .B0 (
                      nx3338)) ;
    AOI21_X0P5M_A12TS ix8864 (.Y (nx8863), .A0 (pc_buf_9), .A1 (nx3228), .B0 (
                      nx8865)) ;
    NOR2_X0P5A_A12TS ix8866 (.Y (nx8865), .A (nx3228), .B (pc_buf_9)) ;
    NOR2_X0P5A_A12TS ix3339 (.Y (nx3338), .A (nx8826), .B (nx8863)) ;
    NAND2_X0P5A_A12TS ix8869 (.Y (nx8868), .A (nx3246), .B (nx3344)) ;
    NOR2_X0P5A_A12TS ix8872 (.Y (nx8871), .A (nx3158), .B (pc_9)) ;
    OAI211_X0P5M_A12TS ix8874 (.Y (nx8873), .A0 (nx3156), .A1 (pc_9), .B0 (
                       nx8875), .C0 (nx3146)) ;
    NAND2_X0P5A_A12TS ix8876 (.Y (nx8875), .A (pc_9), .B (nx3156)) ;
    AOI211_X0P5M_A12TS ix3303 (.Y (nx3302), .A0 (nx8832), .A1 (nx8842), .B0 (
                       nx8705), .C0 (nx3296)) ;
    NOR2_X0P5A_A12TS ix3297 (.Y (nx3296), .A (nx8842), .B (nx8832)) ;
    NAND2_X0P5A_A12TS ix8880 (.Y (nx8879), .A (istb_t), .B (iadr_t_9)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_9 (.Q (iadr_t_9), .CK (wb_clk_i), .D (des2_1)
                        , .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_9)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_10 (.Q (iadr_t_10), .CK (wb_clk_i), .D (
                        des2_2), .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_10)
                        ) ;
    NAND2_X0P5A_A12TS ix8887 (.Y (nx8886), .A (nx7555), .B (nx3410)) ;
    OAI21_X0P5M_A12TS ix3411 (.Y (nx3410), .A0 (nx8889), .A1 (nx5672), .B0 (
                      nx8921)) ;
    INV_X0P5B_A12TS ix8890 (.Y (nx8889), .A (pc_buf_10)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_10 (.Q (pc_buf_10), .CK (wb_clk_i), .D (
                        nx3426), .R (wb_rst_i), .SE (NOT_nx2554), .SI (pc_buf_10
                        )) ;
    NAND4_X0P5A_A12TS ix3427 (.Y (nx3426), .A (nx8893), .B (nx8895), .C (nx8897)
                      , .D (nx8914)) ;
    AOI222_X0P5M_A12TS ix8894 (.Y (nx8893), .A0 (des_acc_2), .A1 (NOT_nx2430), .B0 (
                       des2_2), .B1 (nx2558), .C0 (nx7537), .C1 (nx3410)) ;
    AOI32_X0P5M_A12TS ix8896 (.Y (nx8895), .A0 (op1_n_7), .A1 (pc_wr_sel_2), .A2 (
                      NOT_nx2552), .B0 (op2_n_2), .B1 (nx3184)) ;
    AO21A1AI2_X0P5M_A12TS ix8898 (.Y (nx8897), .A0 (pc_10), .A1 (nx3274), .B0 (
                          nx8912), .C0 (nx3168)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_10 (.Q (pc_10), .CK (wb_clk_i), .D (nx6994), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8902 (.Y (nx8901), .A0 (pc_buf_10), .A1 (pc_wr_r2), 
                          .B0 (nx3458), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix3459 (.Y (nx3458), .A0 (nx8904), .A1 (nx8868), .B0 (
                       pc_wr_r2), .C0 (nx3450)) ;
    OAI21_X0P5M_A12TS ix8905 (.Y (nx8904), .A0 (nx3438), .A1 (nx3338), .B0 (
                      nx8908)) ;
    OAI21_X0P5M_A12TS ix3439 (.Y (nx3438), .A0 (nx8889), .A1 (nx8865), .B0 (
                      nx3432)) ;
    NAND2_X0P5A_A12TS ix3433 (.Y (nx3432), .A (nx8865), .B (nx8889)) ;
    NAND2_X0P5A_A12TS ix8909 (.Y (nx8908), .A (nx3338), .B (nx3438)) ;
    NOR2_X0P5A_A12TS ix3451 (.Y (nx3450), .A (nx8868), .B (nx8904)) ;
    NOR2_X0P5A_A12TS ix8913 (.Y (nx8912), .A (nx3274), .B (pc_10)) ;
    OAI211_X0P5M_A12TS ix8915 (.Y (nx8914), .A0 (nx3266), .A1 (pc_10), .B0 (
                       nx8919), .C0 (nx3146)) ;
    NAND2B_X0P7M_A12TS ix8918 (.Y (nx8917), .AN (nx8815), .B (pc_8)) ;
    NAND2_X0P5A_A12TS ix8920 (.Y (nx8919), .A (pc_10), .B (nx3266)) ;
    OAI211_X0P5M_A12TS ix8922 (.Y (nx8921), .A0 (nx3296), .A1 (pc_buf_10), .B0 (
                       nx5672), .C0 (nx8923)) ;
    NAND2_X0P5A_A12TS ix8924 (.Y (nx8923), .A (pc_buf_10), .B (nx3296)) ;
    OAI21_X0P5M_A12TS ix1316 (.Y (wbi_adr_o[11]), .A0 (istb_t), .A1 (nx8926), .B0 (
                      nx8966)) ;
    AOI21_X0P5M_A12TS ix8927 (.Y (nx8926), .A0 (pc_buf_11), .A1 (nx8705), .B0 (
                      nx3508)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_11 (.Q (pc_buf_11), .CK (wb_clk_i), .D (
                        nx3528), .R (wb_rst_i), .SE (NOT_nx2552), .SI (pc_buf_11
                        )) ;
    OAI211_X0P5M_A12TS ix3529 (.Y (nx3528), .A0 (pc_wr_dup_1371), .A1 (nx8926), 
                       .B0 (nx8930), .C0 (nx8932)) ;
    AOI22_X0P5M_A12TS ix8931 (.Y (nx8930), .A0 (des2_3), .A1 (nx2454), .B0 (
                      op2_n_3), .B1 (nx2478)) ;
    AOI21_X0P5M_A12TS ix8933 (.Y (nx8932), .A0 (des_acc_3), .A1 (nx2464), .B0 (
                      nx3496)) ;
    OAI21_X0P5M_A12TS ix3497 (.Y (nx3496), .A0 (nx8935), .A1 (nx8937), .B0 (
                      nx8956)) ;
    NAND2_X0P5A_A12TS ix8936 (.Y (nx8935), .A (nx3058), .B (nx2446)) ;
    AOI21_X0P5M_A12TS ix8938 (.Y (nx8937), .A0 (pc_11), .A1 (nx3376), .B0 (
                      nx8954)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_11 (.Q (pc_11), .CK (wb_clk_i), .D (nx3564), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_11)) ;
    INV_X0P5B_A12TS ix8942 (.Y (nx8941), .A (pc_buf_11)) ;
    OAI211_X0P5M_A12TS ix8944 (.Y (nx8943), .A0 (nx3548), .A1 (nx3450), .B0 (
                       nx7603), .C0 (nx8951)) ;
    AOI21_X0P5M_A12TS ix3549 (.Y (nx3548), .A0 (nx8946), .A1 (nx8908), .B0 (
                      nx3542)) ;
    AOI21_X0P5M_A12TS ix8947 (.Y (nx8946), .A0 (pc_buf_11), .A1 (nx3432), .B0 (
                      nx8948)) ;
    NOR2_X0P5A_A12TS ix8949 (.Y (nx8948), .A (nx3432), .B (pc_buf_11)) ;
    NOR2_X0P5A_A12TS ix3543 (.Y (nx3542), .A (nx8908), .B (nx8946)) ;
    NAND2_X0P5A_A12TS ix8952 (.Y (nx8951), .A (nx3450), .B (nx3548)) ;
    NOR2_X0P5A_A12TS ix8955 (.Y (nx8954), .A (nx3376), .B (pc_11)) ;
    OAI211_X0P5M_A12TS ix8957 (.Y (nx8956), .A0 (nx3368), .A1 (pc_11), .B0 (
                       nx8959), .C0 (nx3476)) ;
    NAND2_X0P5A_A12TS ix8960 (.Y (nx8959), .A (pc_11), .B (nx3368)) ;
    AOI211_X0P5M_A12TS ix3509 (.Y (nx3508), .A0 (nx8923), .A1 (nx8941), .B0 (
                       nx8705), .C0 (nx3502)) ;
    NOR2_X0P5A_A12TS ix3503 (.Y (nx3502), .A (nx8941), .B (nx8923)) ;
    NAND2_X0P5A_A12TS ix8967 (.Y (nx8966), .A (istb_t), .B (iadr_t_11)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_11 (.Q (iadr_t_11), .CK (wb_clk_i), .D (
                        des2_3), .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_11)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_12 (.Q (iadr_t_12), .CK (wb_clk_i), .D (
                        des2_4), .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_12)
                        ) ;
    NAND2_X0P5A_A12TS ix8974 (.Y (nx8973), .A (nx7555), .B (nx3610)) ;
    OAI21_X0P5M_A12TS ix3611 (.Y (nx3610), .A0 (nx8976), .A1 (nx5672), .B0 (
                      nx9007)) ;
    INV_X0P5B_A12TS ix8977 (.Y (nx8976), .A (pc_buf_12)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_12 (.Q (pc_buf_12), .CK (wb_clk_i), .D (
                        nx3624), .R (wb_rst_i), .SE (NOT_nx2552), .SI (pc_buf_12
                        )) ;
    NAND4_X0P5A_A12TS ix3625 (.Y (nx3624), .A (nx8980), .B (nx8982), .C (nx9000)
                      , .D (nx9005)) ;
    AOI222_X0P5M_A12TS ix8981 (.Y (nx8980), .A0 (des2_4), .A1 (nx2454), .B0 (
                       nx7537), .B1 (nx3610), .C0 (op2_n_4), .C1 (nx2478)) ;
    AO21A1AI2_X0P5M_A12TS ix8983 (.Y (nx8982), .A0 (pc_12), .A1 (nx3486), .B0 (
                          nx8997), .C0 (nx3484)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_12 (.Q (pc_12), .CK (wb_clk_i), .D (nx7034), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix8987 (.Y (nx8986), .A0 (pc_buf_12), .A1 (pc_wr_r2), 
                          .B0 (nx3656), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix3657 (.Y (nx3656), .A0 (nx8989), .A1 (nx8951), .B0 (
                       pc_wr_r2), .C0 (nx3648)) ;
    OAI21_X0P5M_A12TS ix8990 (.Y (nx8989), .A0 (nx3636), .A1 (nx3542), .B0 (
                      nx8993)) ;
    OAI21_X0P5M_A12TS ix3637 (.Y (nx3636), .A0 (nx8976), .A1 (nx8948), .B0 (
                      nx3630)) ;
    NAND2_X0P5A_A12TS ix3631 (.Y (nx3630), .A (nx8948), .B (nx8976)) ;
    NAND2_X0P5A_A12TS ix8994 (.Y (nx8993), .A (nx3542), .B (nx3636)) ;
    NOR2_X0P5A_A12TS ix3649 (.Y (nx3648), .A (nx8951), .B (nx8989)) ;
    NOR2_X0P5A_A12TS ix8998 (.Y (nx8997), .A (nx3486), .B (pc_12)) ;
    OAI211_X0P5M_A12TS ix9001 (.Y (nx9000), .A0 (nx3472), .A1 (pc_12), .B0 (
                       nx9003), .C0 (nx3476)) ;
    NAND2_X0P5A_A12TS ix9004 (.Y (nx9003), .A (pc_12), .B (nx3472)) ;
    NAND2_X0P5A_A12TS ix9006 (.Y (nx9005), .A (des_acc_4), .B (nx2464)) ;
    OAI211_X0P5M_A12TS ix9008 (.Y (nx9007), .A0 (nx3502), .A1 (pc_buf_12), .B0 (
                       nx5672), .C0 (nx9009)) ;
    NAND2_X0P5A_A12TS ix9010 (.Y (nx9009), .A (pc_buf_12), .B (nx3502)) ;
    OAI21_X0P5M_A12TS ix1318 (.Y (wbi_adr_o[13]), .A0 (istb_t), .A1 (nx9012), .B0 (
                      nx9047)) ;
    AOI21_X0P5M_A12TS ix9013 (.Y (nx9012), .A0 (pc_buf_13), .A1 (nx8705), .B0 (
                      nx3700)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_13 (.Q (pc_buf_13), .CK (wb_clk_i), .D (
                        nx3720), .R (wb_rst_i), .SE (NOT_nx2552), .SI (pc_buf_13
                        )) ;
    OAI211_X0P5M_A12TS ix3721 (.Y (nx3720), .A0 (pc_wr_dup_1371), .A1 (nx9012), 
                       .B0 (nx9016), .C0 (nx9018)) ;
    AOI22_X0P5M_A12TS ix9017 (.Y (nx9016), .A0 (des2_5), .A1 (nx2454), .B0 (
                      op2_n_5), .B1 (nx2478)) ;
    AOI21_X0P5M_A12TS ix9019 (.Y (nx9018), .A0 (des_acc_5), .A1 (nx2464), .B0 (
                      nx3688)) ;
    OAI21_X0P5M_A12TS ix3689 (.Y (nx3688), .A0 (nx8935), .A1 (nx9021), .B0 (
                      nx9040)) ;
    AOI21_X0P5M_A12TS ix9022 (.Y (nx9021), .A0 (pc_13), .A1 (nx3582), .B0 (
                      nx9038)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_13 (.Q (pc_13), .CK (wb_clk_i), .D (nx3756), .R (
                        wb_rst_i), .SE (NOT_nx2426), .SI (pc_13)) ;
    INV_X0P5B_A12TS ix9026 (.Y (nx9025), .A (pc_buf_13)) ;
    OAI211_X0P5M_A12TS ix9028 (.Y (nx9027), .A0 (nx3740), .A1 (nx3648), .B0 (
                       nx7603), .C0 (nx9035)) ;
    AOI21_X0P5M_A12TS ix3741 (.Y (nx3740), .A0 (nx9030), .A1 (nx8993), .B0 (
                      nx3734)) ;
    AOI21_X0P5M_A12TS ix9031 (.Y (nx9030), .A0 (pc_buf_13), .A1 (nx3630), .B0 (
                      nx9032)) ;
    NOR2_X0P5A_A12TS ix9033 (.Y (nx9032), .A (nx3630), .B (pc_buf_13)) ;
    NOR2_X0P5A_A12TS ix3735 (.Y (nx3734), .A (nx8993), .B (nx9030)) ;
    NAND2_X0P5A_A12TS ix9036 (.Y (nx9035), .A (nx3648), .B (nx3740)) ;
    NOR2_X0P5A_A12TS ix9039 (.Y (nx9038), .A (nx3582), .B (pc_13)) ;
    OAI211_X0P5M_A12TS ix9041 (.Y (nx9040), .A0 (nx3574), .A1 (pc_13), .B0 (
                       nx9043), .C0 (nx3476)) ;
    NAND2_X0P5A_A12TS ix9044 (.Y (nx9043), .A (pc_13), .B (nx3574)) ;
    AOI211_X0P5M_A12TS ix3701 (.Y (nx3700), .A0 (nx9009), .A1 (nx9025), .B0 (
                       nx8705), .C0 (nx3694)) ;
    NOR2_X0P5A_A12TS ix3695 (.Y (nx3694), .A (nx9025), .B (nx9009)) ;
    NAND2_X0P5A_A12TS ix9048 (.Y (nx9047), .A (istb_t), .B (iadr_t_13)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_13 (.Q (iadr_t_13), .CK (wb_clk_i), .D (
                        des2_5), .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_13)
                        ) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_14 (.Q (iadr_t_14), .CK (wb_clk_i), .D (
                        des2_6), .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_14)
                        ) ;
    NAND2_X0P5A_A12TS ix9055 (.Y (nx9054), .A (nx7555), .B (nx3802)) ;
    OAI21_X0P5M_A12TS ix3803 (.Y (nx3802), .A0 (nx9057), .A1 (nx5672), .B0 (
                      nx9085)) ;
    INV_X0P5B_A12TS ix9058 (.Y (nx9057), .A (pc_buf_14)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_14 (.Q (pc_buf_14), .CK (wb_clk_i), .D (
                        nx3816), .R (wb_rst_i), .SE (NOT_nx2552), .SI (pc_buf_14
                        )) ;
    NAND4_X0P5A_A12TS ix3817 (.Y (nx3816), .A (nx9061), .B (nx9063), .C (nx9078)
                      , .D (nx9083)) ;
    AOI222_X0P5M_A12TS ix9062 (.Y (nx9061), .A0 (des2_6), .A1 (nx2454), .B0 (
                       nx7537), .B1 (nx3802), .C0 (op2_n_6), .C1 (nx2478)) ;
    AO21A1AI2_X0P5M_A12TS ix9064 (.Y (nx9063), .A0 (pc_14), .A1 (nx3678), .B0 (
                          nx9076), .C0 (nx3484)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_14 (.Q (pc_14), .CK (wb_clk_i), .D (nx7074), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix9068 (.Y (nx9067), .A0 (pc_buf_14), .A1 (pc_wr_r2), 
                          .B0 (nx3848), .C0 (nx1518)) ;
    AOI211_X0P5M_A12TS ix3849 (.Y (nx3848), .A0 (nx9070), .A1 (nx9035), .B0 (
                       pc_wr_r2), .C0 (nx3840)) ;
    XNOR2_X0P5M_A12TS ix9071 (.Y (nx9070), .A (nx3734), .B (nx3828)) ;
    OAI21_X0P5M_A12TS ix3829 (.Y (nx3828), .A0 (nx9057), .A1 (nx9032), .B0 (
                      nx3822)) ;
    NAND2_X0P5A_A12TS ix3823 (.Y (nx3822), .A (nx9032), .B (nx9057)) ;
    NOR2_X0P5A_A12TS ix3841 (.Y (nx3840), .A (nx9035), .B (nx9070)) ;
    NOR2_X0P5A_A12TS ix9077 (.Y (nx9076), .A (nx3678), .B (pc_14)) ;
    OAI211_X0P5M_A12TS ix9079 (.Y (nx9078), .A0 (nx3670), .A1 (pc_14), .B0 (
                       nx9081), .C0 (nx3476)) ;
    NAND2_X0P5A_A12TS ix9082 (.Y (nx9081), .A (pc_14), .B (nx3670)) ;
    NAND2_X0P5A_A12TS ix9084 (.Y (nx9083), .A (des_acc_6), .B (nx2464)) ;
    OAI211_X0P5M_A12TS ix9086 (.Y (nx9085), .A0 (nx3694), .A1 (pc_buf_14), .B0 (
                       nx5672), .C0 (nx9087)) ;
    NAND2_X0P5A_A12TS ix9088 (.Y (nx9087), .A (pc_buf_14), .B (nx3694)) ;
    OAI21_X0P5M_A12TS ix4381 (.Y (wbi_adr_o[15]), .A0 (istb_t), .A1 (nx9090), .B0 (
                      nx9112)) ;
    MXIT2_X0P5M_A12TS ix9091 (.Y (nx9090), .A (pc_buf_15), .B (nx3872), .S0 (
                      nx5672)) ;
    SDFFRPQ_X0P5M_A12TS reg_pc_buf_15 (.Q (pc_buf_15), .CK (wb_clk_i), .D (
                        nx3894), .R (wb_rst_i), .SE (NOT_nx2552), .SI (pc_buf_15
                        )) ;
    OAI211_X0P5M_A12TS ix3895 (.Y (nx3894), .A0 (pc_wr_dup_1371), .A1 (nx9090), 
                       .B0 (nx9094), .C0 (nx9109)) ;
    AOI22_X0P5M_A12TS ix9095 (.Y (nx9094), .A0 (nx3886), .A1 (nx3476), .B0 (
                      nx3882), .B1 (nx3484)) ;
    XNOR2_X0P5M_A12TS ix3887 (.Y (nx3886), .A (nx9081), .B (pc_15)) ;
    DFFRPQ_X0P5M_A12TS reg_pc_15 (.Q (pc_15), .CK (wb_clk_i), .D (nx7094), .R (
                       wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix9100 (.Y (nx9099), .A0 (pc_buf_15), .A1 (pc_wr_r2), 
                          .B0 (nx3908), .C0 (nx1518)) ;
    NOR2_X0P5A_A12TS ix3909 (.Y (nx3908), .A (pc_wr_r2), .B (nx9102)) ;
    XOR2_X0P5M_A12TS ix9103 (.Y (nx9102), .A (nx3840), .B (nx9104)) ;
    XNOR3_X0P5M_A12TS ix9105 (.Y (nx9104), .A (nx9106), .B (pc_buf_15), .C (
                      nx3822)) ;
    NAND2_X0P5A_A12TS ix9107 (.Y (nx9106), .A (nx3734), .B (nx3828)) ;
    XOR2_X0P5M_A12TS ix3883 (.Y (nx3882), .A (pc_15), .B (nx9076)) ;
    AOI222_X0P5M_A12TS ix9110 (.Y (nx9109), .A0 (des2_7), .A1 (nx2454), .B0 (
                       des_acc_7), .B1 (nx2464), .C0 (op2_n_7), .C1 (nx2478)) ;
    XNOR2_X0P5M_A12TS ix3873 (.Y (nx3872), .A (pc_buf_15), .B (nx9087)) ;
    NAND2_X0P5A_A12TS ix9113 (.Y (nx9112), .A (istb_t), .B (iadr_t_15)) ;
    SDFFRPQ_X0P5M_A12TS reg_iadr_t_15 (.Q (iadr_t_15), .CK (wb_clk_i), .D (
                        des2_7), .R (wb_rst_i), .SE (NOT_nx226), .SI (iadr_t_15)
                        ) ;
    MXT2_X0P5M_A12TS ix1320 (.Y (ram_out_0), .A (sfr_out_0), .B (ram_data_0), .S0 (
                     nx9116)) ;
    NAND2B_X0P7M_A12TS ix9117 (.Y (nx9116), .AN (rd_ind), .B (rd_addr_r)) ;
    DFFRPQ_X0P5M_A12TS reg_rd_ind (.Q (rd_ind), .CK (wb_clk_i), .D (nx2324), .R (
                       wb_rst_i)) ;
    INV_X0P5B_A12TS ix9121 (.Y (nx9120), .A (ram_rd_sel_0)) ;
    DFFRPQ_X0P5M_A12TS reg_rd_addr_r (.Q (rd_addr_r), .CK (wb_clk_i), .D (
                       rd_addr_7), .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix2421 (.Y (rd_addr_7), .A (nx9124), .B (nx9129)) ;
    AOI21_X0P5M_A12TS ix9125 (.Y (nx9124), .A0 (op2_n_7), .A1 (nx1504), .B0 (
                      ram_rd_sel_2)) ;
    NOR3_X0P5A_A12TS ix1321 (.Y (nx1504), .A (ram_rd_sel_0), .B (ram_rd_sel_2), 
                     .C (nx9127)) ;
    INV_X0P5B_A12TS ix9128 (.Y (nx9127), .A (ram_rd_sel_1)) ;
    AOI32_X0P5M_A12TS ix9130 (.Y (nx9129), .A0 (sp_7), .A1 (ram_rd_sel_1), .A2 (
                      ram_rd_sel_0), .B0 (ri_7), .B1 (nx1465)) ;
    NOR2_X0P5A_A12TS ix1322 (.Y (nx1465), .A (ram_rd_sel_1), .B (nx9120)) ;
    MXT2_X0P5M_A12TS ix4409 (.Y (ram_out_1), .A (sfr_out_1), .B (ram_data_1), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix4417 (.Y (ram_out_2), .A (sfr_out_2), .B (ram_data_2), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix1324 (.Y (ram_out_3), .A (sfr_out_3), .B (ram_data_3), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix1326 (.Y (ram_out_4), .A (sfr_out_4), .B (ram_data_4), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix4441 (.Y (ram_out_5), .A (sfr_out_5), .B (ram_data_5), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix1327 (.Y (ram_out_6), .A (sfr_out_6), .B (ram_data_6), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix1328 (.Y (ram_out_7), .A (sfr_out_7), .B (ram_data_7), .S0 (
                     nx9116)) ;
    MXT2_X0P5M_A12TS ix4465 (.Y (bit_out), .A (sfr_bit), .B (bit_data), .S0 (
                     nx9116)) ;
    NAND2_X2M_A12TS ix1329 (.Y (wr_addr_0), .A (nx9141), .B (nx9149)) ;
    AOI22_X0P5M_A12TS ix9142 (.Y (nx9141), .A0 (rn_r_0), .A1 (nx1654), .B0 (
                      imm_r_0), .B1 (nx1638)) ;
    DFFRPQ_X0P5M_A12TS reg_rn_r_0 (.Q (rn_r_0), .CK (wb_clk_i), .D (op1_cur_0), 
                       .R (wb_rst_i)) ;
    NOR3_X0P5A_A12TS ix1655 (.Y (nx1654), .A (ram_wr_sel_0), .B (ram_wr_sel_2), 
                     .C (ram_wr_sel_1)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_0 (.Q (imm_r_0), .CK (wb_clk_i), .D (op2_n_0), 
                       .R (wb_rst_i)) ;
    NOR3_X0P5A_A12TS ix1639 (.Y (nx1638), .A (ram_wr_sel_1), .B (ram_wr_sel_2), 
                     .C (nx9147)) ;
    INV_X0P5B_A12TS ix9148 (.Y (nx9147), .A (ram_wr_sel_0)) ;
    AOI222_X0P5M_A12TS ix9150 (.Y (nx9149), .A0 (sp_w_0), .A1 (nx1624), .B0 (
                       imm2_r_0), .B1 (nx1602), .C0 (ri_r_0), .C1 (nx1616)) ;
    NOR3_X0P5A_A12TS ix1625 (.Y (nx1624), .A (nx7505), .B (ram_wr_sel_2), .C (
                     nx9147)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_0 (.Q (imm2_r_0), .CK (wb_clk_i), .D (op3_n_0)
                       , .R (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix1603 (.Y (nx1602), .A (ram_wr_sel_1), .B (nx9154)) ;
    NAND2_X0P5A_A12TS ix9155 (.Y (nx9154), .A (ram_wr_sel_2), .B (ram_wr_sel_0)
                      ) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_0 (.Q (ri_r_0), .CK (wb_clk_i), .D (ri_0), .R (
                       wb_rst_i)) ;
    NAND2_X1M_A12TS ix1330 (.Y (wr_addr_1), .A (nx9159), .B (nx9163)) ;
    AOI22_X0P5M_A12TS ix9160 (.Y (nx9159), .A0 (rn_r_1), .A1 (nx1654), .B0 (
                      imm_r_1), .B1 (nx1638)) ;
    DFFRPQ_X0P5M_A12TS reg_rn_r_1 (.Q (rn_r_1), .CK (wb_clk_i), .D (op1_cur_1), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_1 (.Q (imm_r_1), .CK (wb_clk_i), .D (op2_n_1), 
                       .R (wb_rst_i)) ;
    AOI222_X0P5M_A12TS ix9164 (.Y (nx9163), .A0 (sp_w_1), .A1 (nx1624), .B0 (
                       imm2_r_1), .B1 (nx1602), .C0 (ri_r_1), .C1 (nx1616)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_1 (.Q (imm2_r_1), .CK (wb_clk_i), .D (op3_n_1)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_1 (.Q (ri_r_1), .CK (wb_clk_i), .D (ri_1), .R (
                       wb_rst_i)) ;
    NAND2_X1M_A12TS ix1831 (.Y (wr_addr_2), .A (nx9168), .B (nx9172)) ;
    AOI22_X0P5M_A12TS ix9169 (.Y (nx9168), .A0 (rn_r_2), .A1 (nx1654), .B0 (
                      imm_r_2), .B1 (nx1638)) ;
    DFFRPQ_X0P5M_A12TS reg_rn_r_2 (.Q (rn_r_2), .CK (wb_clk_i), .D (op1_cur_2), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_2 (.Q (imm_r_2), .CK (wb_clk_i), .D (op2_n_2), 
                       .R (wb_rst_i)) ;
    AOI222_X0P5M_A12TS ix9173 (.Y (nx9172), .A0 (sp_w_2), .A1 (nx1624), .B0 (
                       imm2_r_2), .B1 (nx1602), .C0 (ri_r_2), .C1 (nx1616)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_2 (.Q (imm2_r_2), .CK (wb_clk_i), .D (op3_n_2)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_2 (.Q (ri_r_2), .CK (wb_clk_i), .D (ri_2), .R (
                       wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix1331 (.Y (wr_addr_3), .A (nx9177), .B (nx9181)) ;
    AOI22_X0P5M_A12TS ix9178 (.Y (nx9177), .A0 (rn_r_3), .A1 (nx1654), .B0 (
                      imm_r_3), .B1 (nx1638)) ;
    DFFRPQ_X0P5M_A12TS reg_rn_r_3 (.Q (rn_r_3), .CK (wb_clk_i), .D (bank_sel_0)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_3 (.Q (imm_r_3), .CK (wb_clk_i), .D (op2_n_3), 
                       .R (wb_rst_i)) ;
    AOI222_X0P5M_A12TS ix9182 (.Y (nx9181), .A0 (sp_w_3), .A1 (nx1624), .B0 (
                       imm2_r_3), .B1 (nx1602), .C0 (ri_r_3), .C1 (nx1616)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_3 (.Q (imm2_r_3), .CK (wb_clk_i), .D (op3_n_3)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_3 (.Q (ri_r_3), .CK (wb_clk_i), .D (ri_3), .R (
                       wb_rst_i)) ;
    NAND4_X1M_A12TS ix1332 (.Y (wr_addr_4), .A (nx9186), .B (nx9190), .C (nx9193
                    ), .D (nx9199)) ;
    AOI22_X0P5M_A12TS ix9187 (.Y (nx9186), .A0 (rn_r_4), .A1 (nx1654), .B0 (
                      imm_r_4), .B1 (nx1638)) ;
    DFFRPQ_X0P5M_A12TS reg_rn_r_4 (.Q (rn_r_4), .CK (wb_clk_i), .D (bank_sel_1)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_4 (.Q (imm_r_4), .CK (wb_clk_i), .D (op2_n_4), 
                       .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix9191 (.Y (nx9190), .A (ri_r_4), .B (nx1616)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_4 (.Q (ri_r_4), .CK (wb_clk_i), .D (ri_4), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix9194 (.Y (nx9193), .A0 (imm2_r_4), .A1 (ram_wr_sel_1), .B0 (
                      nx1507)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_4 (.Q (imm2_r_4), .CK (wb_clk_i), .D (op3_n_4)
                       , .R (wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix9200 (.Y (nx9199), .A (sp_w_4), .B (ram_wr_sel_1), .C (
                      ram_wr_sel_0)) ;
    OAI211_X1M_A12TS ix2111 (.Y (wr_addr_5), .A0 (nx9202), .A1 (nx9205), .B0 (
                     nx9207), .C0 (nx9210)) ;
    INV_X0P5B_A12TS ix9203 (.Y (nx9202), .A (ri_r_5)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_5 (.Q (ri_r_5), .CK (wb_clk_i), .D (ri_5), .R (
                       wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix9206 (.Y (nx9205), .A (nx9147), .B (wr_ind)) ;
    OAI211_X0P5M_A12TS ix9208 (.Y (nx9207), .A0 (imm2_r_5), .A1 (ram_wr_sel_1), 
                       .B0 (ram_wr_sel_2), .C0 (ram_wr_sel_0)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_5 (.Q (imm2_r_5), .CK (wb_clk_i), .D (op3_n_5)
                       , .R (wb_rst_i)) ;
    AOI32_X0P5M_A12TS ix9211 (.Y (nx9210), .A0 (wr_ind), .A1 (sp_w_5), .A2 (
                      ram_wr_sel_0), .B0 (imm_r_5), .B1 (nx2056)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_5 (.Q (imm_r_5), .CK (wb_clk_i), .D (op2_n_5), 
                       .R (wb_rst_i)) ;
    NOR3_X0P5A_A12TS ix2057 (.Y (nx2056), .A (ram_wr_sel_2), .B (ram_wr_sel_1), 
                     .C (nx9147)) ;
    OAI211_X0P5M_A12TS ix2209 (.Y (wr_addr_6), .A0 (nx9215), .A1 (nx9205), .B0 (
                       nx9218), .C0 (nx9221)) ;
    INV_X0P5B_A12TS ix9216 (.Y (nx9215), .A (ri_r_6)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_6 (.Q (ri_r_6), .CK (wb_clk_i), .D (ri_6), .R (
                       wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix9219 (.Y (nx9218), .A0 (imm2_r_6), .A1 (ram_wr_sel_1), 
                       .B0 (ram_wr_sel_2), .C0 (ram_wr_sel_0)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_6 (.Q (imm2_r_6), .CK (wb_clk_i), .D (op3_n_6)
                       , .R (wb_rst_i)) ;
    AOI32_X0P5M_A12TS ix9222 (.Y (nx9221), .A0 (wr_ind), .A1 (sp_w_6), .A2 (
                      ram_wr_sel_0), .B0 (imm_r_6), .B1 (nx2056)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_6 (.Q (imm_r_6), .CK (wb_clk_i), .D (op2_n_6), 
                       .R (wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix1333 (.Y (wr_addr_7), .A (nx9225), .B (nx9228)) ;
    OAI211_X0P5M_A12TS ix9226 (.Y (nx9225), .A0 (imm2_r_7), .A1 (ram_wr_sel_1), 
                       .B0 (ram_wr_sel_2), .C0 (ram_wr_sel_0)) ;
    DFFRPQ_X0P5M_A12TS reg_imm2_r_7 (.Q (imm2_r_7), .CK (wb_clk_i), .D (op3_n_7)
                       , .R (wb_rst_i)) ;
    AOI222_X0P5M_A12TS ix9229 (.Y (nx9228), .A0 (imm_r_7), .A1 (nx2056), .B0 (
                       sp_w_7), .B1 (nx1900), .C0 (ri_r_7), .C1 (nx1616)) ;
    DFFRPQ_X0P5M_A12TS reg_imm_r_7 (.Q (imm_r_7), .CK (wb_clk_i), .D (op2_n_7), 
                       .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ri_r_7 (.Q (ri_r_7), .CK (wb_clk_i), .D (ri_7), .R (
                       wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix1463 (.Y (rd_addr_0), .A (nx9234), .B (nx9239)) ;
    AOI22_X0P5M_A12TS ix9235 (.Y (nx9234), .A0 (sp_0), .A1 (nx1456), .B0 (
                      op2_n_0), .B1 (nx1504)) ;
    NOR2_X0P5A_A12TS ix1334 (.Y (nx1456), .A (ram_rd_sel_2), .B (nx9237)) ;
    NAND2_X0P5A_A12TS ix9238 (.Y (nx9237), .A (ram_rd_sel_1), .B (ram_rd_sel_0)
                      ) ;
    AOI22_X0P5M_A12TS ix9240 (.Y (nx9239), .A0 (op1_cur_0), .A1 (nx1468), .B0 (
                      ri_0), .B1 (nx1467)) ;
    NOR3_X0P5A_A12TS ix1335 (.Y (nx1468), .A (ram_rd_sel_0), .B (ram_rd_sel_2), 
                     .C (ram_rd_sel_1)) ;
    NOR3_X0P5A_A12TS ix1336 (.Y (nx1467), .A (ram_rd_sel_2), .B (ram_rd_sel_1), 
                     .C (nx9120)) ;
    OAI211_X0P5M_A12TS ix2321 (.Y (rd_addr_1), .A0 (nx9244), .A1 (nx9246), .B0 (
                       nx9250), .C0 (nx9252)) ;
    INV_X0P5B_A12TS ix9245 (.Y (nx9244), .A (op1_cur_1)) ;
    INV_X0P5B_A12TS ix9249 (.Y (nx9248), .A (ram_rd_sel_2)) ;
    AOI22_X0P5M_A12TS ix9251 (.Y (nx9250), .A0 (sp_1), .A1 (nx1456), .B0 (
                      op2_n_1), .B1 (nx1504)) ;
    OAI21_X0P5M_A12TS ix9253 (.Y (nx9252), .A0 (ri_1), .A1 (ram_rd_sel_2), .B0 (
                      nx1465)) ;
    NAND2_X0P5A_A12TS ix1337 (.Y (rd_addr_2), .A (nx9255), .B (nx9257)) ;
    AOI22_X0P5M_A12TS ix9256 (.Y (nx9255), .A0 (sp_2), .A1 (nx1456), .B0 (
                      op2_n_2), .B1 (nx1504)) ;
    AOI22_X0P5M_A12TS ix9258 (.Y (nx9257), .A0 (op1_cur_2), .A1 (nx1468), .B0 (
                      ri_2), .B1 (nx1467)) ;
    NAND2_X0P5A_A12TS ix1559 (.Y (rd_addr_3), .A (nx9260), .B (nx9262)) ;
    AOI22_X0P5M_A12TS ix9261 (.Y (nx9260), .A0 (sp_3), .A1 (nx1456), .B0 (
                      op2_n_3), .B1 (nx1504)) ;
    AOI22_X0P5M_A12TS ix9263 (.Y (nx9262), .A0 (bank_sel_0), .A1 (nx1468), .B0 (
                      ri_3), .B1 (nx1467)) ;
    AO1B2_X0P5M_A12TS ix1338 (.Y (rd_addr_4), .A0N (nx9265), .B0 (ri_4), .B1 (
                      nx1517)) ;
    AOI31_X0P5M_A12TS ix9266 (.Y (nx9265), .A0 (nx2332), .A1 (sp_4), .A2 (nx2324
                      ), .B0 (nx2356)) ;
    OAI21_X0P5M_A12TS ix2333 (.Y (nx2332), .A0 (ram_rd_sel_1), .A1 (ram_rd_sel_0
                      ), .B0 (nx9237)) ;
    AOI21_X0P5M_A12TS ix2357 (.Y (nx2356), .A0 (nx9269), .A1 (nx9248), .B0 (
                      ram_rd_sel_0)) ;
    MXIT2_X0P5M_A12TS ix9270 (.Y (nx9269), .A (op2_n_4), .B (bank_sel_1), .S0 (
                      nx2332)) ;
    NOR2_X0P5A_A12TS ix1339 (.Y (nx1517), .A (nx9272), .B (nx2332)) ;
    NAND2_X0P5A_A12TS ix9273 (.Y (nx9272), .A (nx9248), .B (ram_rd_sel_0)) ;
    OAI211_X0P5M_A12TS ix2385 (.Y (rd_addr_5), .A0 (nx8183), .A1 (nx9275), .B0 (
                       nx9277), .C0 (nx9279)) ;
    AO21A1AI2_X0P5M_A12TS ix9278 (.Y (nx9277), .A0 (sp_5), .A1 (ram_rd_sel_0), .B0 (
                          ram_rd_sel_2), .C0 (nx2332)) ;
    NAND4_X0P5A_A12TS ix9280 (.Y (nx9279), .A (nx9248), .B (nx9120), .C (op2_n_5
                      ), .D (ram_rd_sel_1)) ;
    OAI211_X0P5M_A12TS ix2409 (.Y (rd_addr_6), .A0 (nx8189), .A1 (nx9275), .B0 (
                       nx9282), .C0 (nx9284)) ;
    AO21A1AI2_X0P5M_A12TS ix9283 (.Y (nx9282), .A0 (op2_n_6), .A1 (ram_rd_sel_1)
                          , .B0 (ram_rd_sel_2), .C0 (nx9120)) ;
    OAI211_X0P5M_A12TS ix9285 (.Y (nx9284), .A0 (ram_rd_sel_2), .A1 (sp_6), .B0 (
                       ram_rd_sel_0), .C0 (ram_rd_sel_1)) ;
    INV_X0P5B_A12TS ix3679 (.Y (nx3678), .A (nx9038)) ;
    INV_X0P5B_A12TS ix3671 (.Y (nx3670), .A (nx9043)) ;
    INV_X0P5B_A12TS ix3583 (.Y (nx3582), .A (nx8997)) ;
    INV_X0P5B_A12TS ix3575 (.Y (nx3574), .A (nx9003)) ;
    INV_X0P5B_A12TS ix3487 (.Y (nx3486), .A (nx8954)) ;
    INV_X0P5B_A12TS ix3485 (.Y (nx3484), .A (nx8935)) ;
    INV_X0P5B_A12TS ix3473 (.Y (nx3472), .A (nx8959)) ;
    INV_X0P5B_A12TS ix3377 (.Y (nx3376), .A (nx8912)) ;
    INV_X0P5B_A12TS ix3369 (.Y (nx3368), .A (nx8919)) ;
    INV_X0P5B_A12TS ix3309 (.Y (nx3308), .A (nx8835)) ;
    INV_X0P5B_A12TS ix3275 (.Y (nx3274), .A (nx8871)) ;
    INV_X0P5B_A12TS ix3267 (.Y (nx3266), .A (nx8875)) ;
    INV_X0P5B_A12TS ix3159 (.Y (nx3158), .A (nx8813)) ;
    INV_X0P5B_A12TS ix3157 (.Y (nx3156), .A (nx8917)) ;
    INV_X0P5B_A12TS ix3059 (.Y (nx3058), .A (nx8764)) ;
    INV_X0P5B_A12TS ix2875 (.Y (nx2874), .A (nx8684)) ;
    INV_X0P5B_A12TS ix2711 (.Y (nx2710), .A (nx8628)) ;
    INV_X0P5B_A12TS ix2687 (.Y (nx2686), .A (nx8599)) ;
    INV_X0P5B_A12TS ix2663 (.Y (nx2662), .A (nx8583)) ;
    INV_X0P5B_A12TS ix2659 (.Y (nx2658), .A (nx8620)) ;
    INV_X0P5B_A12TS ix8552 (.Y (nx8551), .A (nx2562)) ;
    INV_X0P5B_A12TS ix2559 (.Y (nx2558), .A (nx8528)) ;
    INV_X0P5B_A12TS ix8582 (.Y (nx8581), .A (nx2504)) ;
    INV_X0P5B_A12TS ix1340 (.Y (nx2438), .A (nx8567)) ;
    INV_X0P5B_A12TS ix8493 (.Y (NOT_nx2430), .A (nx2430)) ;
    INV_X0P5B_A12TS ix8488 (.Y (NOT_nx2426), .A (nx1518)) ;
    INV_X0P5B_A12TS ix9276 (.Y (nx9275), .A (nx1517)) ;
    INV_X0P5B_A12TS ix2325 (.Y (nx2324), .A (nx9272)) ;
    INV_X0P5B_A12TS ix1617 (.Y (nx1616), .A (nx9205)) ;
    INV_X0P5B_A12TS ix1342 (.Y (nx1507), .A (nx9154)) ;
    INV_X0P5B_A12TS ix1343 (.Y (nx1503), .A (nx8369)) ;
    INV_X0P5B_A12TS ix1344 (.Y (nx1493), .A (nx7581)) ;
    INV_X0P5B_A12TS ix1109 (.Y (nx1108), .A (nx8012)) ;
    INV_X0P5B_A12TS ix1345 (.Y (nx1070), .A (nx8071)) ;
    INV_X0P5B_A12TS ix7906 (.Y (nx7905), .A (nx5677)) ;
    INV_X0P5B_A12TS ix1346 (.Y (nx1491), .A (nx8019)) ;
    INV_X0P5B_A12TS ix1348 (.Y (nx1489), .A (nx7965)) ;
    INV_X0P5B_A12TS ix1349 (.Y (nx1486), .A (nx7853)) ;
    INV_X0P5B_A12TS ix823 (.Y (nx822), .A (nx7955)) ;
    INV_X0P5B_A12TS ix8015 (.Y (nx8014), .A (nx778)) ;
    INV_X0P5B_A12TS ix755 (.Y (nx754), .A (nx7766)) ;
    INV_X0P5B_A12TS ix577 (.Y (nx576), .A (nx7903)) ;
    INV_X0P5B_A12TS ix1350 (.Y (nx1480), .A (nx7975)) ;
    INV_X0P5B_A12TS ix1352 (.Y (nx1479), .A (nx7749)) ;
    INV_X0P5B_A12TS ix8032 (.Y (nx8031), .A (nx416)) ;
    INV_X0P5B_A12TS ix393 (.Y (nx392), .A (nx7778)) ;
    INV_X0P5B_A12TS ix389 (.Y (nx388), .A (nx7515)) ;
    INV_X0P5B_A12TS ix1354 (.Y (nx270), .A (nx7572)) ;
    INV_X0P5B_A12TS ix7688 (.Y (nx7687), .A (nx260)) ;
    INV_X0P5B_A12TS ix1356 (.Y (nx1476), .A (nx7654)) ;
    INV_X0P5B_A12TS ix1358 (.Y (nx1475), .A (nx7663)) ;
    INV_X0P5B_A12TS ix7781 (.Y (nx7780), .A (nx1473)) ;
    INV_X0P5B_A12TS ix121 (.Y (nx120), .A (nx7683)) ;
    INV_X0P5B_A12TS ix1360 (.Y (nx1470), .A (nx8069)) ;
    INV_X0P5B_A12TS ix8706 (.Y (nx8705), .A (nx5672)) ;
    INV_X0P5B_A12TS ix37 (.Y (nx36), .A (nx8544)) ;
    INV_X0P5B_A12TS ix27 (.Y (nx26), .A (nx7679)) ;
    INV_X0P5B_A12TS ix1361 (.Y (nx1469), .A (nx7521)) ;
    INV_X0P5B_A12TS ix9247 (.Y (nx9246), .A (nx1468)) ;
    INV_X0P5B_A12TS ix1362 (.Y (op1_n_1), .A (nx8043)) ;
    INV_X0P5B_A12TS ix1364 (.Y (op1_n_2), .A (nx7808)) ;
    INV_X0P5B_A12TS ix773 (.Y (op1_n_4), .A (nx8067)) ;
    INV_X0P5B_A12TS ix1365 (.Y (op1_n_5), .A (nx7704)) ;
    INV_X0P5B_A12TS ix1366 (.Y (op1_n_7), .A (nx7981)) ;
    AO1B2_X0P5M_A12TS ix5825 (.Y (nx5824), .A0N (NOT_nx226), .B0 (istb_t), .B1 (
                      imem_wait)) ;
    OAI31_X0P5M_A12TS ix7979 (.Y (nx1498), .A0 (nx8062), .A1 (nx778), .A2 (
                      nx8031), .B0 (nx9295)) ;
    INV_X0P5B_A12TS ix9294 (.Y (nx9295), .A (nx1497)) ;
    NAND2_X0P5A_A12TS ix8018 (.Y (nx8017), .A (nx7704), .B (op1_n_4)) ;
    OR2_X0P5M_A12TS ix8020 (.Y (nx8019), .A (nx7981), .B (nx7808)) ;
    NAND2_X0P5A_A12TS ix8029 (.Y (nx8028), .A (nx7704), .B (nx7808)) ;
    OR2_X0P5M_A12TS ix779 (.Y (nx778), .A (nx8067), .B (nx7704)) ;
    OR2_X0P5M_A12TS ix8060 (.Y (nx8059), .A (nx7981), .B (nx7704)) ;
    NAND3_X0P5A_A12TS ix8063 (.Y (nx8062), .A (nx7981), .B (op1_n_0), .C (
                      op1_n_2)) ;
    NOR2B_X0P7M_A12TS ix3945 (.Y (nx3944), .AN (nx1485), .B (nx7975)) ;
    AO1B2_X0P5M_A12TS ix4037 (.Y (nx4036), .A0N (nx8155), .B0 (ri_0), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4049 (.Y (nx4048), .A0N (nx8161), .B0 (ri_1), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4061 (.Y (nx4060), .A0N (nx8167), .B0 (ri_2), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4073 (.Y (nx4072), .A0N (nx8173), .B0 (ri_3), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4085 (.Y (nx4084), .A0N (nx8179), .B0 (ri_4), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4097 (.Y (nx4096), .A0N (nx8185), .B0 (ri_5), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4109 (.Y (nx4108), .A0N (nx8191), .B0 (ri_6), .B1 (
                      mem_act_1)) ;
    AO1B2_X0P5M_A12TS ix4121 (.Y (nx4120), .A0N (nx8197), .B0 (mem_act_1), .B1 (
                      ri_7)) ;
    NOR2B_X0P7M_A12TS ix1421 (.Y (nx1420), .AN (nx138), .B (nx7665)) ;
    OAI2XB1_X0P5M_A12TS ix6795 (.Y (nx6794), .A0 (nx1518), .A1N (pc_0), .B0 (
                        nx8478)) ;
    NAND3B_X0P5M_A12TS ix8505 (.Y (nx8504), .AN (pc_wr_sel_1), .B (
                       pc_wr_dup_1371), .C (pc_wr_sel_2)) ;
    OAI2XB1_X0P5M_A12TS ix6815 (.Y (nx6814), .A0 (nx1518), .A1N (pc_1), .B0 (
                        nx8512)) ;
    NAND2B_X0P7M_A12TS ix2563 (.Y (nx2562), .AN (NOT_nx2554), .B (nx8528)) ;
    NOR2B_X0P7M_A12TS ix8555 (.Y (NOT_nx2554), .AN (NOT_nx2552), .B (pc_wr_sel_2
                      )) ;
    CGEN_X1M_A12TS ix8565 (.CO (nx8564), .A (nx8489), .B (nx9297), .CI (nx8502)
                   ) ;
    INV_X0P5B_A12TS ix9296 (.Y (nx9297), .A (pc_1)) ;
    AO1B2_X0P5M_A12TS ix2675 (.Y (nx2674), .A0N (nx8574), .B0 (pc_buf_2), .B1 (
                      pc_wr_r2)) ;
    AO1B2_X0P5M_A12TS ix4237 (.Y (wbi_adr_o[3]), .A0N (nx8592), .B0 (istb_t), .B1 (
                      iadr_t_3)) ;
    AO1B2_X0P5M_A12TS ix2771 (.Y (nx2770), .A0N (nx8610), .B0 (pc_buf_3), .B1 (
                      pc_wr_r2)) ;
    AO1B2_X0P5M_A12TS ix4249 (.Y (wbi_adr_o[4]), .A0N (nx8634), .B0 (istb_t), .B1 (
                      iadr_t_4)) ;
    OAI2XB1_X0P5M_A12TS ix6875 (.Y (nx6874), .A0 (nx1518), .A1N (pc_4), .B0 (
                        nx8652)) ;
    AO21_X0P5M_A12TS ix2839 (.Y (nx2838), .A0 (pc_buf_4), .A1 (pc_buf_3), .B0 (
                     nx8661)) ;
    AO1B2_X0P5M_A12TS ix2955 (.Y (nx2954), .A0N (nx8695), .B0 (pc_buf_5), .B1 (
                      pc_wr_r2)) ;
    AO1B2_X0P5M_A12TS ix4273 (.Y (wbi_adr_o[6]), .A0N (nx8717), .B0 (istb_t), .B1 (
                      iadr_t_6)) ;
    OAI2XB1_X0P5M_A12TS ix6915 (.Y (nx6914), .A0 (nx1518), .A1N (pc_6), .B0 (
                        nx8735)) ;
    AO1B2_X0P5M_A12TS ix3139 (.Y (nx3138), .A0N (nx8775), .B0 (pc_buf_7), .B1 (
                      pc_wr_r2)) ;
    AO1B2_X0P5M_A12TS ix4297 (.Y (wbi_adr_o[8]), .A0N (nx8794), .B0 (istb_t), .B1 (
                      iadr_t_8)) ;
    OAI2XB1_X0P5M_A12TS ix6955 (.Y (nx6954), .A0 (nx1518), .A1N (pc_8), .B0 (
                        nx8819)) ;
    AO1B2_X0P5M_A12TS ix3361 (.Y (nx3360), .A0N (nx8860), .B0 (pc_buf_9), .B1 (
                      pc_wr_r2)) ;
    AO1B2_X0P5M_A12TS ix4321 (.Y (wbi_adr_o[10]), .A0N (nx8886), .B0 (istb_t), .B1 (
                      iadr_t_10)) ;
    OAI2XB1_X0P5M_A12TS ix6995 (.Y (nx6994), .A0 (nx1518), .A1N (pc_10), .B0 (
                        nx8901)) ;
    AO1B2_X0P5M_A12TS ix3565 (.Y (nx3564), .A0N (nx8943), .B0 (pc_buf_11), .B1 (
                      pc_wr_r2)) ;
    AND2_X0P5M_A12TS ix3477 (.Y (nx3476), .A (nx8764), .B (nx2446)) ;
    AO1B2_X0P5M_A12TS ix1367 (.Y (wbi_adr_o[12]), .A0N (nx8973), .B0 (istb_t), .B1 (
                      iadr_t_12)) ;
    OAI2XB1_X0P5M_A12TS ix7035 (.Y (nx7034), .A0 (nx1518), .A1N (pc_12), .B0 (
                        nx8986)) ;
    AO1B2_X0P5M_A12TS ix3757 (.Y (nx3756), .A0N (nx9027), .B0 (pc_buf_13), .B1 (
                      pc_wr_r2)) ;
    AO1B2_X0P5M_A12TS ix4369 (.Y (wbi_adr_o[14]), .A0N (nx9054), .B0 (istb_t), .B1 (
                      iadr_t_14)) ;
    OAI2XB1_X0P5M_A12TS ix7075 (.Y (nx7074), .A0 (nx1518), .A1N (pc_14), .B0 (
                        nx9067)) ;
    OAI2XB1_X0P5M_A12TS ix7095 (.Y (nx7094), .A0 (nx1518), .A1N (pc_15), .B0 (
                        nx9099)) ;
    AND2_X0P5M_A12TS ix1901 (.Y (nx1900), .A (ram_wr_sel_1), .B (ram_wr_sel_0)
                     ) ;
    DFFRPQ_X0P5M_A12TS reg_wr_bit_r_dup_66146 (.Q (wr_bit_r_dup_1790), .CK (
                       wb_clk_i), .D (bit_addr), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_pres_ow (.Q (pres_ow), .CK (wb_clk_i), .D (nx2080), .R (
                       wb_rst_i)) ;
    NOR3_X0P5A_A12TS ix1519 (.Y (nx2080), .A (nx1884), .B (nx2183), .C (
                     prescaler_2)) ;
    NAND2_X0P5A_A12TS ix1523 (.Y (nx1884), .A (prescaler_1), .B (prescaler_0)) ;
    DFFRPQ_X0P5M_A12TS reg_prescaler_1 (.Q (prescaler_1), .CK (wb_clk_i), .D (
                       nx1792), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix2178 (.Y (nx1791), .A (prescaler_0)) ;
    DFFRPQ_X0P5M_A12TS reg_prescaler_0 (.Q (prescaler_0), .CK (wb_clk_i), .D (
                       nx1791), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix2184 (.Y (nx2183), .A (prescaler_3)) ;
    DFFRPQ_X0P5M_A12TS reg_prescaler_3 (.Q (prescaler_3), .CK (wb_clk_i), .D (
                       nx1794), .R (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix1525 (.Y (nx1794), .A (nx2080), .B (nx2187)) ;
    XOR2_X0P5M_A12TS ix2188 (.Y (nx2187), .A (prescaler_3), .B (nx2189)) ;
    NAND3_X0P5A_A12TS ix2190 (.Y (nx2189), .A (prescaler_2), .B (prescaler_1), .C (
                      prescaler_0)) ;
    DFFRPQ_X0P5M_A12TS reg_prescaler_2 (.Q (prescaler_2), .CK (wb_clk_i), .D (
                       nx34), .R (wb_rst_i)) ;
    OA21A1OI2_X0P5M_A12TS ix35 (.Y (nx34), .A0 (nx1884), .A1 (prescaler_3), .B0 (
                          nx2193), .C0 (nx2082)) ;
    INV_X0P5B_A12TS ix2194 (.Y (nx2193), .A (prescaler_2)) ;
    DFFRPQ_X0P5M_A12TS reg_wait_data (.Q (wait_data), .CK (wb_clk_i), .D (
                       NOT_NOT__68049), .R (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix1526 (.Y (NOT_NOT__68049), .A (wait_data), .B (nx1885)) ;
    AOI22_X0P5M_A12TS ix1528 (.Y (nx1885), .A0 (rd_addr_7), .A1 (nx848), .B0 (
                      nx2220), .B1 (nx1838)) ;
    OAI21_X0P5M_A12TS ix1529 (.Y (nx848), .A0 (nx2201), .A1 (nx2203), .B0 (
                      nx1886)) ;
    XNOR2_X0P5M_A12TS ix2202 (.Y (nx2201), .A (wr_sfr_1), .B (wr_sfr_0)) ;
    NAND4_X0P5A_A12TS ix2204 (.Y (nx2203), .A (rd_addr_5), .B (rd_addr_6), .C (
                      nx1801), .D (nx1812)) ;
    NOR2_X0P5A_A12TS ix1530 (.Y (nx1801), .A (rd_addr_3), .B (rd_addr_4)) ;
    NOR3_X0P5A_A12TS ix1531 (.Y (nx1812), .A (rd_addr_2), .B (rd_addr_0), .C (
                     rd_addr_1)) ;
    OAI21_X0P5M_A12TS ix1532 (.Y (nx1886), .A0 (psw_set_1), .A1 (psw_set_0), .B0 (
                      nx1840)) ;
    NOR2_X0P5A_A12TS ix1533 (.Y (nx1840), .A (nx2210), .B (nx2214)) ;
    NAND2_X0P5A_A12TS ix2211 (.Y (nx2210), .A (nx2212), .B (rd_addr_6)) ;
    INV_X0P5B_A12TS ix2213 (.Y (nx2212), .A (rd_addr_5)) ;
    NAND2_X0P5A_A12TS ix2215 (.Y (nx2214), .A (nx1807), .B (nx830)) ;
    NOR2_X0P5A_A12TS ix1536 (.Y (nx1807), .A (rd_addr_3), .B (nx2217)) ;
    INV_X0P5B_A12TS ix2218 (.Y (nx2217), .A (rd_addr_4)) ;
    NOR3_X0P5A_A12TS ix1537 (.Y (nx830), .A (rd_addr_2), .B (rd_addr_0), .C (
                     rd_addr_1)) ;
    NAND4_X0P5A_A12TS ix2221 (.Y (nx2220), .A (nx2222), .B (wr_sfr_1), .C (
                      wr_sfr_0), .D (nx1832)) ;
    INV_X0P5B_A12TS ix2223 (.Y (nx2222), .A (rd_addr_3)) ;
    NOR2_X0P5A_A12TS ix1545 (.Y (nx1832), .A (nx1830), .B (nx2227)) ;
    NAND3_X0P5A_A12TS ix1546 (.Y (nx1830), .A (nx2217), .B (rd_addr_7), .C (
                      nx158)) ;
    NOR2_X0P5A_A12TS ix159 (.Y (nx158), .A (rd_addr_5), .B (rd_addr_6)) ;
    INV_X0P5B_A12TS ix2232 (.Y (nx2231), .A (rd_addr_0)) ;
    OAI211_X0P5M_A12TS ix1549 (.Y (nx1838), .A0 (nx2234), .A1 (nx2236), .B0 (
                       nx2251), .C0 (nx2256)) ;
    NAND3_X0P5A_A12TS ix2235 (.Y (nx2234), .A (wr_bit_r_dup_1790), .B (wr_addr_7
                      ), .C (we)) ;
    NAND2_X0P5A_A12TS ix2237 (.Y (nx2236), .A (nx2238), .B (nx2249)) ;
    NOR3_X0P5A_A12TS ix2239 (.Y (nx2238), .A (nx1799), .B (nx1797), .C (nx1796)
                     ) ;
    XOR2_X0P5M_A12TS ix1550 (.Y (nx1799), .A (wr_addr_4), .B (rd_addr_4)) ;
    XOR2_X0P5M_A12TS ix1552 (.Y (nx1797), .A (wr_addr_5), .B (rd_addr_5)) ;
    NAND3_X0P5A_A12TS ix1553 (.Y (nx1796), .A (nx2243), .B (nx2245), .C (nx2247)
                      ) ;
    XNOR2_X0P5M_A12TS ix2244 (.Y (nx2243), .A (wr_addr_7), .B (rd_addr_7)) ;
    XNOR2_X0P5M_A12TS ix2246 (.Y (nx2245), .A (wr_addr_3), .B (rd_addr_3)) ;
    XNOR2_X0P5M_A12TS ix2248 (.Y (nx2247), .A (wr_addr_6), .B (rd_addr_6)) ;
    NAND3_X0P5A_A12TS ix2250 (.Y (nx2249), .A (rd_addr_2), .B (rd_addr_0), .C (
                      rd_addr_1)) ;
    NAND4_X0P5A_A12TS ix2252 (.Y (nx2251), .A (nx2222), .B (wr_sfr_1), .C (
                      wr_sfr_0), .D (nx1836)) ;
    NOR2_X0P5A_A12TS ix1554 (.Y (nx1836), .A (nx1830), .B (nx2254)) ;
    NAND3_X0P5A_A12TS ix2257 (.Y (nx2256), .A (wr_addr_7), .B (we), .C (nx1834)
                      ) ;
    NOR2_X0P5A_A12TS ix1555 (.Y (nx1834), .A (wr_bit_r_dup_1790), .B (nx2259)) ;
    NAND4_X0P5A_A12TS ix2260 (.Y (nx2259), .A (nx2238), .B (nx2261), .C (nx2263)
                      , .D (nx2265)) ;
    XNOR2_X0P5M_A12TS ix2262 (.Y (nx2261), .A (wr_addr_0), .B (rd_addr_0)) ;
    XNOR2_X0P5M_A12TS ix2264 (.Y (nx2263), .A (wr_addr_2), .B (rd_addr_2)) ;
    XNOR2_X0P5M_A12TS ix2266 (.Y (nx2265), .A (wr_addr_1), .B (rd_addr_1)) ;
    INV_X0P5B_A12TS ix1905 (.Y (comp_wait), .A (nx2268)) ;
    AO21A1AI2_X0P5M_A12TS ix2269 (.Y (nx2268), .A0 (comp_sel_0), .A1 (nx2270), .B0 (
                          nx1883), .C0 (nx2256)) ;
    NAND4B_X0P5M_A12TS ix2271 (.Y (nx2270), .AN (wr_bit_r_dup_1790), .B (we), .C (
                       nx2238), .D (nx96)) ;
    NAND3_X0P5A_A12TS ix1556 (.Y (nx96), .A (wr_addr_1), .B (wr_addr_2), .C (
                      wr_addr_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1561 (.Y (nx1883), .A0 (nx2274), .A1 (nx2284), .B0 (
                          comp_sel_1), .C0 (nx2286)) ;
    OAI31_X0P5M_A12TS ix2275 (.Y (nx2274), .A0 (wr_addr_4), .A1 (nx2276), .A2 (
                      nx1879), .B0 (nx2201)) ;
    INV_X0P5B_A12TS ix2277 (.Y (nx2276), .A (wr_addr_5)) ;
    NAND4_X0P5A_A12TS ix1563 (.Y (nx1879), .A (nx2279), .B (we), .C (wr_addr_7)
                      , .D (wr_addr_6)) ;
    NOR2_X0P5A_A12TS ix2280 (.Y (nx2279), .A (nx1878), .B (wr_addr_3)) ;
    NOR2_X0P5A_A12TS ix1861 (.Y (nx1878), .A (wr_bit_r_dup_1790), .B (nx1888)) ;
    NOR3_X0P5A_A12TS ix1567 (.Y (nx1888), .A (wr_addr_1), .B (wr_addr_2), .C (
                     wr_addr_0)) ;
    INV_X0P5B_A12TS ix2285 (.Y (nx2284), .A (comp_sel_0)) ;
    NAND4B_X0P5M_A12TS ix1568 (.Y (nx2286), .AN (psw_set_0), .B (comp_sel_1), .C (
                       nx2284), .D (nx1881)) ;
    AOI31_X0P5M_A12TS ix1879 (.Y (nx1881), .A0 (wr_addr_4), .A1 (nx2276), .A2 (
                      nx2289), .B0 (psw_set_1)) ;
    DFFRPQ_X0P5M_A12TS reg_bit_out (.Q (sfr_bit), .CK (wb_clk_i), .D (nx758), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix759 (.Y (nx758), .A (nx2293), .B (nx1897), .S0 (nx1805)
                      ) ;
    MXIT2_X0P5M_A12TS ix2294 (.Y (nx2293), .A (desCy), .B (nx704), .S0 (nx2450)
                      ) ;
    NAND4_X0P5A_A12TS ix705 (.Y (nx704), .A (nx2296), .B (nx2354), .C (nx2409), 
                      .D (nx2431)) ;
    AOI221_X0P5M_A12TS ix2297 (.Y (nx2296), .A0 (acc_0), .A1 (nx696), .B0 (nx158
                       ), .B1 (nx688), .C0 (nx624)) ;
    AND4_X0P5M_A12TS ix697 (.Y (nx696), .A (rd_addr_5), .B (rd_addr_6), .C (
                     nx1801), .D (nx1812)) ;
    AO21A1AI2_X0P5M_A12TS ix689 (.Y (nx688), .A0 (nx2300), .A1 (nx2306), .B0 (
                          nx2310), .C0 (nx2312)) ;
    AOI22_X0P5M_A12TS ix2301 (.Y (nx2300), .A0 (tcon_7), .A1 (nx1814), .B0 (
                      tcon_1), .B1 (nx284)) ;
    INV_X0P5B_A12TS ix2304 (.Y (nx2303), .A (rd_addr_1)) ;
    NOR3_X0P5A_A12TS ix285 (.Y (nx284), .A (rd_addr_2), .B (nx2231), .C (
                     rd_addr_1)) ;
    AOI222_X0P5M_A12TS ix2307 (.Y (nx2306), .A0 (tcon_0), .A1 (nx1812), .B0 (
                       tcon_3), .B1 (nx1813), .C0 (tcon_2), .C1 (nx1810)) ;
    NOR3_X0P5A_A12TS ix1571 (.Y (nx1810), .A (rd_addr_2), .B (rd_addr_0), .C (
                     nx2303)) ;
    NAND2_X0P5A_A12TS ix2311 (.Y (nx2310), .A (rd_addr_3), .B (nx2217)) ;
    AOI22_X0P5M_A12TS ix2313 (.Y (nx2312), .A0 (nx1801), .A1 (nx682), .B0 (
                      nx1807), .B1 (nx1827)) ;
    NAND2_X0P5A_A12TS ix683 (.Y (nx682), .A (nx2315), .B (nx2317)) ;
    AOI22_X0P5M_A12TS ix2316 (.Y (nx2315), .A0 (p0_data_7), .A1 (nx1814), .B0 (
                      p0_data_1), .B1 (nx284)) ;
    AOI222_X0P5M_A12TS ix2318 (.Y (nx2317), .A0 (p0_data_0), .A1 (nx1812), .B0 (
                       p0_data_3), .B1 (nx1813), .C0 (p0_data_2), .C1 (nx1810)
                       ) ;
    NAND2_X0P5A_A12TS ix1572 (.Y (nx1827), .A (nx2320), .B (nx1889)) ;
    AOI22_X0P5M_A12TS ix1573 (.Y (nx2320), .A0 (p1_data_7), .A1 (nx1814), .B0 (
                      p1_data_1), .B1 (nx284)) ;
    AOI222_X0P5M_A12TS ix1574 (.Y (nx1889), .A0 (p1_data_0), .A1 (nx1812), .B0 (
                       p1_data_3), .B1 (nx1813), .C0 (p1_data_2), .C1 (nx1810)
                       ) ;
    OAI211_X0P5M_A12TS ix625 (.Y (nx624), .A0 (nx2249), .A1 (nx2325), .B0 (
                       nx2340), .C0 (nx2347)) ;
    AOI21_X0P5M_A12TS ix2326 (.Y (nx2325), .A0 (scon_7), .A1 (nx1809), .B0 (
                      nx560)) ;
    INV_X0P5B_A12TS ix2331 (.Y (nx2330), .A (rd_addr_6)) ;
    OAI22_X0P5M_A12TS ix561 (.Y (nx560), .A0 (nx2210), .A1 (nx2333), .B0 (nx1891
                      ), .B1 (nx2338)) ;
    AOI22_X0P5M_A12TS ix2334 (.Y (nx2333), .A0 (t2con_7), .A1 (nx1806), .B0 (cy)
                      , .B1 (nx1807)) ;
    AOI222_X0P5M_A12TS ix2339 (.Y (nx2338), .A0 (p2_data_7), .A1 (nx1801), .B0 (
                       p3_data_7), .B1 (nx1807), .C0 (ie_7), .C1 (nx1806)) ;
    AO21A1AI2_X0P5M_A12TS ix2341 (.Y (nx2340), .A0 (scon_1), .A1 (nx1809), .B0 (
                          nx1825), .C0 (nx284)) ;
    OAI22_X0P5M_A12TS ix1575 (.Y (nx1825), .A0 (nx2210), .A1 (nx2343), .B0 (
                      nx1891), .B1 (nx2345)) ;
    AOI22_X0P5M_A12TS ix2344 (.Y (nx2343), .A0 (t2con_1), .A1 (nx1806), .B0 (
                      psw_1), .B1 (nx1807)) ;
    AOI222_X0P5M_A12TS ix2346 (.Y (nx2345), .A0 (p2_data_1), .A1 (nx1801), .B0 (
                       p3_data_1), .B1 (nx1807), .C0 (ie_1), .C1 (nx1806)) ;
    AO21A1AI2_X0P5M_A12TS ix2348 (.Y (nx2347), .A0 (scon_2), .A1 (nx1809), .B0 (
                          nx1823), .C0 (nx1810)) ;
    OAI22_X0P5M_A12TS ix1576 (.Y (nx1823), .A0 (nx2210), .A1 (nx2350), .B0 (
                      nx1891), .B1 (nx2352)) ;
    AOI22_X0P5M_A12TS ix2351 (.Y (nx2350), .A0 (t2con_2), .A1 (nx1806), .B0 (
                      psw_2), .B1 (nx1807)) ;
    AOI222_X0P5M_A12TS ix2353 (.Y (nx2352), .A0 (p2_data_2), .A1 (nx1801), .B0 (
                       p3_data_2), .B1 (nx1807), .C0 (ie_2), .C1 (nx1806)) ;
    AOI221_X0P5M_A12TS ix2355 (.Y (nx2354), .A0 (nx1812), .A1 (nx528), .B0 (
                       nx1813), .B1 (nx372), .C0 (nx1822)) ;
    OAI222_X0P5M_A12TS ix529 (.Y (nx528), .A0 (nx2210), .A1 (nx2357), .B0 (
                       nx2359), .B1 (nx2361), .C0 (nx1891), .C1 (nx2363)) ;
    AOI22_X0P5M_A12TS ix2358 (.Y (nx2357), .A0 (t2con_0), .A1 (nx1806), .B0 (p)
                      , .B1 (nx1807)) ;
    INV_X0P5B_A12TS ix2360 (.Y (nx2359), .A (scon_0)) ;
    NAND3_X0P5A_A12TS ix2362 (.Y (nx2361), .A (nx158), .B (rd_addr_3), .C (
                      rd_addr_4)) ;
    AOI222_X0P5M_A12TS ix2364 (.Y (nx2363), .A0 (p2_data_0), .A1 (nx1801), .B0 (
                       p3_data_0), .B1 (nx1807), .C0 (ie_0), .C1 (nx1806)) ;
    OAI222_X0P5M_A12TS ix373 (.Y (nx372), .A0 (nx2210), .A1 (nx2366), .B0 (
                       nx2368), .B1 (nx2361), .C0 (nx1891), .C1 (nx2370)) ;
    AOI22_X0P5M_A12TS ix1577 (.Y (nx2366), .A0 (t2con_3), .A1 (nx1806), .B0 (
                      psw_3), .B1 (nx1807)) ;
    INV_X0P5B_A12TS ix2369 (.Y (nx2368), .A (scon_3)) ;
    AOI222_X0P5M_A12TS ix2371 (.Y (nx2370), .A0 (p2_data_3), .A1 (nx1801), .B0 (
                       p3_data_3), .B1 (nx1807), .C0 (ie_3), .C1 (nx1806)) ;
    OA21A1OI2_X0P5M_A12TS ix1578 (.Y (nx1822), .A0 (nx2373), .A1 (nx2375), .B0 (
                          nx2391), .C0 (rd_addr_0)) ;
    NAND2_X0P5A_A12TS ix2374 (.Y (nx2373), .A (nx2303), .B (rd_addr_2)) ;
    AOI211_X0P5M_A12TS ix2376 (.Y (nx2375), .A0 (scon_4), .A1 (nx1809), .B0 (
                       nx1821), .C0 (nx470)) ;
    AOI21_X0P5M_A12TS ix1579 (.Y (nx1821), .A0 (nx2378), .A1 (nx2380), .B0 (
                      nx1891)) ;
    AOI22_X0P5M_A12TS ix2379 (.Y (nx2378), .A0 (p2_data_4), .A1 (nx1801), .B0 (
                      ie_4), .B1 (nx1806)) ;
    AOI32_X0P5M_A12TS ix2381 (.Y (nx2380), .A0 (rd_addr_4), .A1 (ip_4), .A2 (
                      rd_addr_3), .B0 (p3_data_4), .B1 (nx1807)) ;
    OAI222_X0P5M_A12TS ix471 (.Y (nx470), .A0 (nx2210), .A1 (nx2383), .B0 (
                       nx2385), .B1 (nx2387), .C0 (nx2328), .C1 (nx2389)) ;
    AOI22_X0P5M_A12TS ix2384 (.Y (nx2383), .A0 (tclk), .A1 (nx1806), .B0 (psw_4)
                      , .B1 (nx1807)) ;
    AOI22_X0P5M_A12TS ix2386 (.Y (nx2385), .A0 (b_reg_4), .A1 (rd_addr_4), .B0 (
                      acc_4), .B1 (nx1801)) ;
    NAND2_X0P5A_A12TS ix2388 (.Y (nx2387), .A (rd_addr_5), .B (rd_addr_6)) ;
    AOI222_X0P5M_A12TS ix2390 (.Y (nx2389), .A0 (p0_data_4), .A1 (nx1801), .B0 (
                       p1_data_4), .B1 (nx1807), .C0 (tr0), .C1 (nx1806)) ;
    OAI211_X0P5M_A12TS ix2392 (.Y (nx2391), .A0 (nx1818), .A1 (nx408), .B0 (
                       rd_addr_1), .C0 (rd_addr_2)) ;
    AO21A1AI2_X0P5M_A12TS ix1583 (.Y (nx1818), .A0 (nx1892), .A1 (nx2396), .B0 (
                          nx1891), .C0 (nx2398)) ;
    AOI22_X0P5M_A12TS ix1585 (.Y (nx1892), .A0 (p2_data_6), .A1 (nx1801), .B0 (
                      ie_6), .B1 (nx1806)) ;
    AOI32_X0P5M_A12TS ix2397 (.Y (nx2396), .A0 (rd_addr_4), .A1 (ip_6), .A2 (
                      rd_addr_3), .B0 (p3_data_6), .B1 (nx1807)) ;
    NAND2_X0P5A_A12TS ix2399 (.Y (nx2398), .A (scon_6), .B (nx1809)) ;
    OAI222_X0P5M_A12TS ix409 (.Y (nx408), .A0 (nx2210), .A1 (nx2401), .B0 (
                       nx2403), .B1 (nx2405), .C0 (nx2328), .C1 (nx2407)) ;
    AOI22_X0P5M_A12TS ix2402 (.Y (nx2401), .A0 (t2con_6), .A1 (nx1806), .B0 (
                      srcAc), .B1 (nx1807)) ;
    AOI22_X0P5M_A12TS ix2404 (.Y (nx2403), .A0 (b_reg_6), .A1 (rd_addr_4), .B0 (
                      acc_6), .B1 (nx1801)) ;
    NAND2_X0P5A_A12TS ix2406 (.Y (nx2405), .A (rd_addr_5), .B (rd_addr_6)) ;
    AOI222_X0P5M_A12TS ix2408 (.Y (nx2407), .A0 (p0_data_6), .A1 (nx1801), .B0 (
                       p1_data_6), .B1 (nx1807), .C0 (tr1), .C1 (nx1806)) ;
    AOI31_X0P5M_A12TS ix2410 (.Y (nx2409), .A0 (nx1817), .A1 (rd_addr_5), .A2 (
                      rd_addr_6), .B0 (nx300)) ;
    AO21A1AI2_X0P5M_A12TS ix1587 (.Y (nx1817), .A0 (nx2412), .A1 (nx1893), .B0 (
                          nx2416), .C0 (nx2418)) ;
    AOI22_X0P5M_A12TS ix2413 (.Y (nx2412), .A0 (acc_7), .A1 (nx1814), .B0 (acc_1
                      ), .B1 (nx284)) ;
    AOI22_X0P5M_A12TS ix1588 (.Y (nx1893), .A0 (acc_2), .A1 (nx1810), .B0 (acc_3
                      ), .B1 (nx1813)) ;
    AO1B2_X0P5M_A12TS ix2419 (.Y (nx2418), .A0N (rd_addr_4), .B0 (nx2420), .B1 (
                      nx2422)) ;
    AOI22_X0P5M_A12TS ix1589 (.Y (nx2420), .A0 (b_reg_7), .A1 (nx1814), .B0 (
                      b_reg_1), .B1 (nx284)) ;
    AOI222_X0P5M_A12TS ix2423 (.Y (nx2422), .A0 (b_reg_0), .A1 (nx1812), .B0 (
                       b_reg_3), .B1 (nx1813), .C0 (b_reg_2), .C1 (nx1810)) ;
    AOI211_X0P5M_A12TS ix301 (.Y (nx300), .A0 (nx2425), .A1 (nx2427), .B0 (
                       nx2429), .C0 (nx1891)) ;
    AOI22_X0P5M_A12TS ix2426 (.Y (nx2425), .A0 (ip_7), .A1 (nx1814), .B0 (ip_1)
                      , .B1 (nx284)) ;
    AOI222_X0P5M_A12TS ix2428 (.Y (nx2427), .A0 (ip_0), .A1 (nx1812), .B0 (ip_3)
                       , .B1 (nx1813), .C0 (ip_2), .C1 (nx1810)) ;
    NAND2_X0P5A_A12TS ix2430 (.Y (nx2429), .A (rd_addr_3), .B (rd_addr_4)) ;
    OAI211_X0P5M_A12TS ix2432 (.Y (nx2431), .A0 (nx230), .A1 (nx204), .B0 (
                       rd_addr_0), .C0 (nx236)) ;
    AO21A1AI2_X0P5M_A12TS ix231 (.Y (nx230), .A0 (nx2434), .A1 (nx2436), .B0 (
                          nx1891), .C0 (nx1895)) ;
    AOI22_X0P5M_A12TS ix2435 (.Y (nx2434), .A0 (p2_data_5), .A1 (nx1801), .B0 (
                      ie_5), .B1 (nx1806)) ;
    AOI32_X0P5M_A12TS ix2437 (.Y (nx2436), .A0 (rd_addr_4), .A1 (ip_5), .A2 (
                      rd_addr_3), .B0 (p3_data_5), .B1 (nx1807)) ;
    NAND2_X0P5A_A12TS ix1590 (.Y (nx1895), .A (scon_5), .B (nx1809)) ;
    OAI222_X0P5M_A12TS ix205 (.Y (nx204), .A0 (nx2210), .A1 (nx2441), .B0 (
                       nx2443), .B1 (nx2445), .C0 (nx2328), .C1 (nx2447)) ;
    AOI22_X0P5M_A12TS ix2442 (.Y (nx2441), .A0 (rclk), .A1 (nx1806), .B0 (psw_5)
                      , .B1 (nx1807)) ;
    AOI22_X0P5M_A12TS ix2444 (.Y (nx2443), .A0 (b_reg_5), .A1 (rd_addr_4), .B0 (
                      acc_5), .B1 (nx1801)) ;
    NAND2_X0P5A_A12TS ix2446 (.Y (nx2445), .A (rd_addr_5), .B (rd_addr_6)) ;
    AOI222_X0P5M_A12TS ix2448 (.Y (nx2447), .A0 (p0_data_5), .A1 (nx1801), .B0 (
                       p1_data_5), .B1 (nx1807), .C0 (tcon_5), .C1 (nx1806)) ;
    NAND3B_X0P5M_A12TS ix2451 (.Y (nx2450), .AN (nx2259), .B (we), .C (
                       wr_bit_r_dup_1790)) ;
    AOI211_X0P5M_A12TS ix1591 (.Y (nx1897), .A0 (des1_7), .A1 (nx1814), .B0 (
                       nx1829), .C0 (nx742)) ;
    INV_X0P5B_A12TS ix1595 (.Y (nx1829), .A (nx2455)) ;
    AOI22_X0P5M_A12TS ix2456 (.Y (nx2455), .A0 (des1_1), .A1 (nx284), .B0 (
                      des1_2), .B1 (nx1810)) ;
    OAI211_X0P5M_A12TS ix1598 (.Y (nx742), .A0 (rd_addr_0), .A1 (nx2458), .B0 (
                       nx2460), .C0 (nx1899)) ;
    AOI32_X0P5M_A12TS ix2459 (.Y (nx2458), .A0 (rd_addr_2), .A1 (des1_6), .A2 (
                      rd_addr_1), .B0 (des1_4), .B1 (nx236)) ;
    AOI22_X0P5M_A12TS ix2461 (.Y (nx2460), .A0 (des1_0), .A1 (nx1812), .B0 (
                      des1_3), .B1 (nx1813)) ;
    NAND3_X0P5A_A12TS ix1600 (.Y (nx1899), .A (nx236), .B (des1_5), .C (
                      rd_addr_0)) ;
    OAI21_X0P5M_A12TS ix1601 (.Y (nx1805), .A0 (nx2465), .A1 (nx2467), .B0 (
                      nx2270)) ;
    NAND3B_X0P5M_A12TS ix2466 (.Y (nx2465), .AN (wr_sfr_1), .B (wr_sfr_0), .C (
                       rd_addr_7)) ;
    NAND3_X0P5A_A12TS ix2468 (.Y (nx2467), .A (nx1801), .B (rd_addr_5), .C (
                      rd_addr_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_0 (.Q (sfr_out_0), .CK (wb_clk_i), .D (nx1865)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_0)
                        ) ;
    NAND4_X0P5A_A12TS ix1602 (.Y (nx1865), .A (nx2471), .B (nx1902), .C (nx1905)
                      , .D (nx2505)) ;
    AOI222_X0P5M_A12TS ix2472 (.Y (nx2471), .A0 (b_reg_0), .A1 (nx1864), .B0 (
                       des_acc_0), .B1 (nx1833), .C0 (acc_0), .C1 (nx1841)) ;
    NOR3_X0P5A_A12TS ix1605 (.Y (nx1864), .A (nx2214), .B (nx2212), .C (nx2330)
                     ) ;
    AOI222_X0P5M_A12TS ix1607 (.Y (nx1902), .A0 (th1_0), .A1 (nx1030), .B0 (p), 
                       .B1 (nx1840), .C0 (sp_0), .C1 (nx1034)) ;
    NOR3_X0P5A_A12TS ix1609 (.Y (nx1030), .A (nx2481), .B (nx2231), .C (nx2373)
                     ) ;
    NAND3_X0P5A_A12TS ix2482 (.Y (nx2481), .A (rd_addr_3), .B (nx2217), .C (
                      nx158)) ;
    NOR2_X0P5A_A12TS ix1610 (.Y (nx1034), .A (nx1904), .B (nx2486)) ;
    NAND3_X0P5A_A12TS ix2487 (.Y (nx2486), .A (nx1801), .B (nx2220), .C (nx158)
                      ) ;
    AND3_X0P5M_A12TS ix1611 (.Y (nx1905), .A (nx2490), .B (nx2495), .C (nx2499)
                     ) ;
    AOI222_X0P5M_A12TS ix2491 (.Y (nx2490), .A0 (th0_0), .A1 (nx1016), .B0 (
                       tl1_0), .B1 (nx1863), .C0 (dptr_hi_0), .C1 (nx1861)) ;
    NOR3_X0P5A_A12TS ix1614 (.Y (nx1016), .A (nx2481), .B (rd_addr_0), .C (
                     nx2373)) ;
    NOR2_X0P5A_A12TS ix1009 (.Y (nx1863), .A (nx2254), .B (nx2481)) ;
    NOR2_X0P5A_A12TS ix1618 (.Y (nx1861), .A (nx2254), .B (nx2486)) ;
    AOI22_X0P5M_A12TS ix2496 (.Y (nx2495), .A0 (tl0_0), .A1 (nx1860), .B0 (
                      tmod_0), .B1 (nx1858)) ;
    NOR2_X0P5A_A12TS ix997 (.Y (nx1860), .A (nx2227), .B (nx2481)) ;
    NOR2_X0P5A_A12TS ix993 (.Y (nx1858), .A (nx1904), .B (nx2481)) ;
    AOI22_X0P5M_A12TS ix2500 (.Y (nx2499), .A0 (tcon_0), .A1 (nx1857), .B0 (
                      pcon_0), .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix981 (.Y (nx1857), .A (nx2328), .B (nx2502)) ;
    NAND2_X0P5A_A12TS ix2503 (.Y (nx2502), .A (nx1806), .B (nx830)) ;
    NOR2_X0P5A_A12TS ix977 (.Y (nx1856), .A (nx2249), .B (nx2486)) ;
    NOR2_X0P5A_A12TS ix2506 (.Y (nx2505), .A (nx1855), .B (nx918)) ;
    NAND3_X0P5A_A12TS ix973 (.Y (nx1855), .A (nx2508), .B (nx2515), .C (nx2521)
                      ) ;
    AOI222_X0P5M_A12TS ix2509 (.Y (nx2508), .A0 (p1_data_0), .A1 (nx964), .B0 (
                       tl2_0), .B1 (nx960), .C0 (th2_0), .C1 (nx1853)) ;
    NOR2_X0P5A_A12TS ix965 (.Y (nx964), .A (nx2328), .B (nx2214)) ;
    NOR3_X0P5A_A12TS ix961 (.Y (nx960), .A (nx1907), .B (rd_addr_0), .C (nx2373)
                     ) ;
    NAND3_X0P5A_A12TS ix1620 (.Y (nx1907), .A (nx2212), .B (rd_addr_6), .C (
                      nx1806)) ;
    NOR3_X0P5A_A12TS ix1622 (.Y (nx1853), .A (nx1907), .B (nx2231), .C (nx2373)
                     ) ;
    AOI22_X0P5M_A12TS ix2516 (.Y (nx2515), .A0 (p0_data_0), .A1 (nx932), .B0 (
                      dptr_lo_0), .B1 (nx942)) ;
    NOR2_X0P5A_A12TS ix943 (.Y (nx942), .A (nx2227), .B (nx2486)) ;
    AOI22_X0P5M_A12TS ix2522 (.Y (nx2521), .A0 (ie_0), .A1 (nx924), .B0 (
                      rcap2h_0), .B1 (nx920)) ;
    NOR2_X0P5A_A12TS ix925 (.Y (nx924), .A (nx1891), .B (nx2502)) ;
    NOR2_X0P5A_A12TS ix921 (.Y (nx920), .A (nx2254), .B (nx1907)) ;
    NAND3_X0P5A_A12TS ix919 (.Y (nx918), .A (nx2526), .B (nx1908), .C (nx2536)
                      ) ;
    AOI222_X0P5M_A12TS ix2527 (.Y (nx2526), .A0 (t2con_0), .A1 (nx1851), .B0 (
                       rcap2l_0), .B1 (nx894), .C0 (ip_0), .C1 (nx1848)) ;
    NOR2_X0P5A_A12TS ix1623 (.Y (nx1851), .A (nx2210), .B (nx2502)) ;
    NOR2_X0P5A_A12TS ix1627 (.Y (nx894), .A (nx2227), .B (nx1907)) ;
    AND4_X0P5M_A12TS ix1629 (.Y (nx1848), .A (nx1814), .B (nx2220), .C (nx1804)
                     , .D (nx1807)) ;
    NOR2_X0P5A_A12TS ix1632 (.Y (nx1804), .A (nx2212), .B (rd_addr_6)) ;
    AOI22_X0P5M_A12TS ix1633 (.Y (nx1908), .A0 (p3_data_0), .A1 (nx1846), .B0 (
                      p2_data_0), .B1 (nx1845)) ;
    NOR2_X0P5A_A12TS ix1636 (.Y (nx1846), .A (nx1891), .B (nx2214)) ;
    AOI22_X0P5M_A12TS ix2537 (.Y (nx2536), .A0 (sbuf_0), .A1 (nx1844), .B0 (
                      scon_0), .B1 (nx1843)) ;
    NOR3_X0P5A_A12TS ix1637 (.Y (nx1844), .A (nx2361), .B (nx1833), .C (nx1904)
                     ) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_1 (.Q (sfr_out_1), .CK (wb_clk_i), .D (nx1170)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_1)
                        ) ;
    NAND4_X0P5A_A12TS ix1171 (.Y (nx1170), .A (nx2542), .B (nx2544), .C (nx2546)
                      , .D (nx2554)) ;
    AOI222_X0P5M_A12TS ix2543 (.Y (nx2542), .A0 (b_reg_1), .A1 (nx1864), .B0 (
                       des_acc_1), .B1 (nx1833), .C0 (acc_1), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix1641 (.Y (nx2544), .A0 (th1_1), .A1 (nx1030), .B0 (
                       psw_1), .B1 (nx1840), .C0 (sp_1), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix2547 (.Y (nx2546), .A (nx2548), .B (nx2550), .C (nx2552)
                     ) ;
    AOI222_X0P5M_A12TS ix2549 (.Y (nx2548), .A0 (th0_1), .A1 (nx1016), .B0 (
                       tl1_1), .B1 (nx1863), .C0 (dptr_hi_1), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix2551 (.Y (nx2550), .A0 (tl0_1), .A1 (nx1860), .B0 (
                      tmod_1), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix2553 (.Y (nx2552), .A0 (tcon_1), .A1 (nx1857), .B0 (
                      pcon_1), .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix2555 (.Y (nx2554), .A (nx1116), .B (nx1090)) ;
    NAND3_X0P5A_A12TS ix1117 (.Y (nx1116), .A (nx2557), .B (nx2559), .C (nx2561)
                      ) ;
    AOI222_X0P5M_A12TS ix2558 (.Y (nx2557), .A0 (p1_data_1), .A1 (nx964), .B0 (
                       tl2_1), .B1 (nx960), .C0 (th2_1), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2560 (.Y (nx2559), .A0 (p0_data_1), .A1 (nx932), .B0 (
                      dptr_lo_1), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2562 (.Y (nx2561), .A0 (ie_1), .A1 (nx924), .B0 (
                      rcap2h_1), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1643 (.Y (nx1090), .A (nx2564), .B (nx2566), .C (nx2568)
                      ) ;
    AOI222_X0P5M_A12TS ix2565 (.Y (nx2564), .A0 (t2con_1), .A1 (nx1851), .B0 (
                       rcap2l_1), .B1 (nx894), .C0 (ip_1), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix2567 (.Y (nx2566), .A0 (p3_data_1), .A1 (nx1846), .B0 (
                      p2_data_1), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix2569 (.Y (nx2568), .A0 (sbuf_1), .A1 (nx1844), .B0 (
                      scon_1), .B1 (nx1843)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_2 (.Q (sfr_out_2), .CK (wb_clk_i), .D (nx1280)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_2)
                        ) ;
    NAND4_X0P5A_A12TS ix1645 (.Y (nx1280), .A (nx1909), .B (nx2574), .C (nx2576)
                      , .D (nx2584)) ;
    AOI222_X0P5M_A12TS ix1648 (.Y (nx1909), .A0 (b_reg_2), .A1 (nx1864), .B0 (
                       des_acc_2), .B1 (nx1833), .C0 (acc_2), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix2575 (.Y (nx2574), .A0 (th1_2), .A1 (nx1030), .B0 (
                       psw_2), .B1 (nx1840), .C0 (sp_2), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix2577 (.Y (nx2576), .A (nx2578), .B (nx1910), .C (nx2582)
                     ) ;
    AOI222_X0P5M_A12TS ix2579 (.Y (nx2578), .A0 (th0_2), .A1 (nx1016), .B0 (
                       tl1_2), .B1 (nx1863), .C0 (dptr_hi_2), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix1649 (.Y (nx1910), .A0 (tl0_2), .A1 (nx1860), .B0 (
                      tmod_2), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix2583 (.Y (nx2582), .A0 (tcon_2), .A1 (nx1857), .B0 (
                      pcon_2), .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix2585 (.Y (nx2584), .A (nx1226), .B (nx1200)) ;
    NAND3_X0P5A_A12TS ix1227 (.Y (nx1226), .A (nx2587), .B (nx2589), .C (nx2591)
                      ) ;
    AOI222_X0P5M_A12TS ix2588 (.Y (nx2587), .A0 (p1_data_2), .A1 (nx964), .B0 (
                       tl2_2), .B1 (nx960), .C0 (th2_2), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2590 (.Y (nx2589), .A0 (p0_data_2), .A1 (nx932), .B0 (
                      dptr_lo_2), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2592 (.Y (nx2591), .A0 (ie_2), .A1 (nx924), .B0 (
                      rcap2h_2), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1650 (.Y (nx1200), .A (nx2594), .B (nx2596), .C (nx2598)
                      ) ;
    AOI222_X0P5M_A12TS ix2595 (.Y (nx2594), .A0 (t2con_2), .A1 (nx1851), .B0 (
                       rcap2l_2), .B1 (nx894), .C0 (ip_2), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix2597 (.Y (nx2596), .A0 (p3_data_2), .A1 (nx1846), .B0 (
                      p2_data_2), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix2599 (.Y (nx2598), .A0 (sbuf_2), .A1 (nx1844), .B0 (
                      scon_2), .B1 (nx1843)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_3 (.Q (sfr_out_3), .CK (wb_clk_i), .D (nx1390)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_3)
                        ) ;
    NAND4_X0P5A_A12TS ix1391 (.Y (nx1390), .A (nx2602), .B (nx1912), .C (nx2606)
                      , .D (nx2614)) ;
    AOI222_X0P5M_A12TS ix2603 (.Y (nx2602), .A0 (b_reg_3), .A1 (nx1864), .B0 (
                       des_acc_3), .B1 (nx1833), .C0 (acc_3), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix1651 (.Y (nx1912), .A0 (th1_3), .A1 (nx1030), .B0 (
                       psw_3), .B1 (nx1840), .C0 (sp_3), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix2607 (.Y (nx2606), .A (nx2608), .B (nx2610), .C (nx1913)
                     ) ;
    AOI222_X0P5M_A12TS ix2609 (.Y (nx2608), .A0 (th0_3), .A1 (nx1016), .B0 (
                       tl1_3), .B1 (nx1863), .C0 (dptr_hi_3), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix2611 (.Y (nx2610), .A0 (tl0_3), .A1 (nx1860), .B0 (
                      tmod_3), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix1653 (.Y (nx1913), .A0 (tcon_3), .A1 (nx1857), .B0 (
                      pcon_3), .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix2615 (.Y (nx2614), .A (nx1336), .B (nx1310)) ;
    NAND3_X0P5A_A12TS ix1656 (.Y (nx1336), .A (nx2617), .B (nx2619), .C (nx2621)
                      ) ;
    AOI222_X0P5M_A12TS ix2618 (.Y (nx2617), .A0 (p1_data_3), .A1 (nx964), .B0 (
                       tl2_3), .B1 (nx960), .C0 (th2_3), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2620 (.Y (nx2619), .A0 (p0_data_3), .A1 (nx932), .B0 (
                      dptr_lo_3), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2622 (.Y (nx2621), .A0 (ie_3), .A1 (nx924), .B0 (
                      rcap2h_3), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1657 (.Y (nx1310), .A (nx2624), .B (nx2626), .C (nx2628)
                      ) ;
    AOI222_X0P5M_A12TS ix2625 (.Y (nx2624), .A0 (t2con_3), .A1 (nx1851), .B0 (
                       rcap2l_3), .B1 (nx894), .C0 (ip_3), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix2627 (.Y (nx2626), .A0 (p3_data_3), .A1 (nx1846), .B0 (
                      p2_data_3), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix2629 (.Y (nx2628), .A0 (sbuf_3), .A1 (nx1844), .B0 (
                      scon_3), .B1 (nx1843)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_4 (.Q (sfr_out_4), .CK (wb_clk_i), .D (nx1869)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_4)
                        ) ;
    NAND4_X0P5A_A12TS ix1501 (.Y (nx1869), .A (nx2632), .B (nx2634), .C (nx2636)
                      , .D (nx2644)) ;
    AOI222_X0P5M_A12TS ix2633 (.Y (nx2632), .A0 (b_reg_4), .A1 (nx1864), .B0 (
                       des_acc_4), .B1 (nx1833), .C0 (acc_4), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix2635 (.Y (nx2634), .A0 (th1_4), .A1 (nx1030), .B0 (
                       psw_4), .B1 (nx1840), .C0 (sp_4), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix2637 (.Y (nx2636), .A (nx1915), .B (nx2640), .C (nx2642)
                     ) ;
    AOI222_X0P5M_A12TS ix1660 (.Y (nx1915), .A0 (th0_4), .A1 (nx1016), .B0 (
                       tl1_4), .B1 (nx1863), .C0 (dptr_hi_4), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix2641 (.Y (nx2640), .A0 (tl0_4), .A1 (nx1860), .B0 (
                      tmod_4), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix2643 (.Y (nx2642), .A0 (tr0), .A1 (nx1857), .B0 (pcon_4)
                      , .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix2645 (.Y (nx2644), .A (nx1446), .B (nx1867)) ;
    NAND3_X0P5A_A12TS ix1447 (.Y (nx1446), .A (nx2647), .B (nx2649), .C (nx2651)
                      ) ;
    AOI222_X0P5M_A12TS ix2648 (.Y (nx2647), .A0 (p1_data_4), .A1 (nx964), .B0 (
                       tl2_4), .B1 (nx960), .C0 (th2_4), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2650 (.Y (nx2649), .A0 (p0_data_4), .A1 (nx932), .B0 (
                      dptr_lo_4), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2652 (.Y (nx2651), .A0 (ie_4), .A1 (nx924), .B0 (
                      rcap2h_4), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1663 (.Y (nx1867), .A (nx2654), .B (nx2656), .C (nx1916)
                      ) ;
    AOI222_X0P5M_A12TS ix2655 (.Y (nx2654), .A0 (tclk), .A1 (nx1851), .B0 (
                       rcap2l_4), .B1 (nx894), .C0 (ip_4), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix2657 (.Y (nx2656), .A0 (p3_data_4), .A1 (nx1846), .B0 (
                      p2_data_4), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix1666 (.Y (nx1916), .A0 (sbuf_4), .A1 (nx1844), .B0 (
                      scon_4), .B1 (nx1843)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_5 (.Q (sfr_out_5), .CK (wb_clk_i), .D (nx1610)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_5)
                        ) ;
    NAND4_X0P5A_A12TS ix1667 (.Y (nx1610), .A (nx1918), .B (nx2664), .C (nx2666)
                      , .D (nx1919)) ;
    AOI222_X0P5M_A12TS ix1668 (.Y (nx1918), .A0 (b_reg_5), .A1 (nx1864), .B0 (
                       des_acc_5), .B1 (nx1833), .C0 (acc_5), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix2665 (.Y (nx2664), .A0 (th1_5), .A1 (nx1030), .B0 (
                       psw_5), .B1 (nx1840), .C0 (sp_5), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix2667 (.Y (nx2666), .A (nx2668), .B (nx2670), .C (nx2672)
                     ) ;
    AOI222_X0P5M_A12TS ix2669 (.Y (nx2668), .A0 (th0_5), .A1 (nx1016), .B0 (
                       tl1_5), .B1 (nx1863), .C0 (dptr_hi_5), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix2671 (.Y (nx2670), .A0 (tl0_5), .A1 (nx1860), .B0 (
                      tmod_5), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix2673 (.Y (nx2672), .A0 (tcon_5), .A1 (nx1857), .B0 (
                      pcon_5), .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix1670 (.Y (nx1919), .A (nx1871), .B (nx1530)) ;
    NAND3_X0P5A_A12TS ix1671 (.Y (nx1871), .A (nx2677), .B (nx2679), .C (nx2681)
                      ) ;
    AOI222_X0P5M_A12TS ix2678 (.Y (nx2677), .A0 (p1_data_5), .A1 (nx964), .B0 (
                       tl2_5), .B1 (nx960), .C0 (th2_5), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2680 (.Y (nx2679), .A0 (p0_data_5), .A1 (nx932), .B0 (
                      dptr_lo_5), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2682 (.Y (nx2681), .A0 (ie_5), .A1 (nx924), .B0 (
                      rcap2h_5), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1674 (.Y (nx1530), .A (nx2684), .B (nx1921), .C (nx2688)
                      ) ;
    AOI222_X0P5M_A12TS ix2685 (.Y (nx2684), .A0 (rclk), .A1 (nx1851), .B0 (
                       rcap2l_5), .B1 (nx894), .C0 (ip_5), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix1676 (.Y (nx1921), .A0 (p3_data_5), .A1 (nx1846), .B0 (
                      p2_data_5), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix2689 (.Y (nx2688), .A0 (sbuf_5), .A1 (nx1844), .B0 (
                      scon_5), .B1 (nx1843)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_6 (.Q (sfr_out_6), .CK (wb_clk_i), .D (nx1720)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_6)
                        ) ;
    NAND4_X0P5A_A12TS ix1721 (.Y (nx1720), .A (nx2692), .B (nx2694), .C (nx1923)
                      , .D (nx2704)) ;
    AOI222_X0P5M_A12TS ix2693 (.Y (nx2692), .A0 (b_reg_6), .A1 (nx1864), .B0 (
                       des_acc_6), .B1 (nx1833), .C0 (acc_6), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix2695 (.Y (nx2694), .A0 (th1_6), .A1 (nx1030), .B0 (
                       srcAc), .B1 (nx1840), .C0 (sp_6), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix1678 (.Y (nx1923), .A (nx2698), .B (nx2700), .C (nx2702)
                     ) ;
    AOI222_X0P5M_A12TS ix2699 (.Y (nx2698), .A0 (th0_6), .A1 (nx1016), .B0 (
                       tl1_6), .B1 (nx1863), .C0 (dptr_hi_6), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix2701 (.Y (nx2700), .A0 (tl0_6), .A1 (nx1860), .B0 (
                      tmod_6), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix2703 (.Y (nx2702), .A0 (tr1), .A1 (nx1857), .B0 (pcon_6)
                      , .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix2705 (.Y (nx2704), .A (nx1666), .B (nx1640)) ;
    NAND3_X0P5A_A12TS ix1679 (.Y (nx1666), .A (nx2707), .B (nx2709), .C (nx2711)
                      ) ;
    AOI222_X0P5M_A12TS ix2708 (.Y (nx2707), .A0 (p1_data_6), .A1 (nx964), .B0 (
                       tl2_6), .B1 (nx960), .C0 (th2_6), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2710 (.Y (nx2709), .A0 (p0_data_6), .A1 (nx932), .B0 (
                      dptr_lo_6), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2712 (.Y (nx2711), .A0 (ie_6), .A1 (nx924), .B0 (
                      rcap2h_6), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1681 (.Y (nx1640), .A (nx2714), .B (nx2716), .C (nx2718)
                      ) ;
    AOI222_X0P5M_A12TS ix2715 (.Y (nx2714), .A0 (t2con_6), .A1 (nx1851), .B0 (
                       rcap2l_6), .B1 (nx894), .C0 (ip_6), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix2717 (.Y (nx2716), .A0 (p3_data_6), .A1 (nx1846), .B0 (
                      p2_data_6), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix2719 (.Y (nx2718), .A0 (sbuf_6), .A1 (nx1844), .B0 (
                      scon_6), .B1 (nx1843)) ;
    SDFFRPQ_X0P5M_A12TS reg_dat0_7 (.Q (sfr_out_7), .CK (wb_clk_i), .D (nx1876)
                        , .R (wb_rst_i), .SE (NOT_NOT__68049), .SI (sfr_out_7)
                        ) ;
    NAND4_X0P5A_A12TS ix1684 (.Y (nx1876), .A (nx1925), .B (nx2724), .C (nx2726)
                      , .D (nx2734)) ;
    AOI222_X0P5M_A12TS ix1687 (.Y (nx1925), .A0 (b_reg_7), .A1 (nx1864), .B0 (
                       des_acc_7), .B1 (nx1833), .C0 (acc_7), .C1 (nx1841)) ;
    AOI222_X0P5M_A12TS ix2725 (.Y (nx2724), .A0 (th1_7), .A1 (nx1030), .B0 (cy)
                       , .B1 (nx1840), .C0 (sp_7), .C1 (nx1034)) ;
    AND3_X0P5M_A12TS ix2727 (.Y (nx2726), .A (nx2728), .B (nx1927), .C (nx2732)
                     ) ;
    AOI222_X0P5M_A12TS ix2729 (.Y (nx2728), .A0 (th0_7), .A1 (nx1016), .B0 (
                       tl1_7), .B1 (nx1863), .C0 (dptr_hi_7), .C1 (nx1861)) ;
    AOI22_X0P5M_A12TS ix1689 (.Y (nx1927), .A0 (tl0_7), .A1 (nx1860), .B0 (
                      tmod_7), .B1 (nx1858)) ;
    AOI22_X0P5M_A12TS ix2733 (.Y (nx2732), .A0 (tcon_7), .A1 (nx1857), .B0 (
                      pcon_7), .B1 (nx1856)) ;
    NOR2_X0P5A_A12TS ix2735 (.Y (nx2734), .A (nx1875), .B (nx1874)) ;
    NAND3_X0P5A_A12TS ix1691 (.Y (nx1875), .A (nx2737), .B (nx2739), .C (nx2741)
                      ) ;
    AOI222_X0P5M_A12TS ix2738 (.Y (nx2737), .A0 (p1_data_7), .A1 (nx964), .B0 (
                       tl2_7), .B1 (nx960), .C0 (th2_7), .C1 (nx1853)) ;
    AOI22_X0P5M_A12TS ix2740 (.Y (nx2739), .A0 (p0_data_7), .A1 (nx932), .B0 (
                      dptr_lo_7), .B1 (nx942)) ;
    AOI22_X0P5M_A12TS ix2742 (.Y (nx2741), .A0 (ie_7), .A1 (nx924), .B0 (
                      rcap2h_7), .B1 (nx920)) ;
    NAND3_X0P5A_A12TS ix1692 (.Y (nx1874), .A (nx2744), .B (nx1928), .C (nx2748)
                      ) ;
    AOI222_X0P5M_A12TS ix2745 (.Y (nx2744), .A0 (t2con_7), .A1 (nx1851), .B0 (
                       rcap2l_7), .B1 (nx894), .C0 (ip_7), .C1 (nx1848)) ;
    AOI22_X0P5M_A12TS ix1693 (.Y (nx1928), .A0 (p3_data_7), .A1 (nx1846), .B0 (
                      p2_data_7), .B1 (nx1845)) ;
    AOI22_X0P5M_A12TS ix2749 (.Y (nx2748), .A0 (sbuf_7), .A1 (nx1844), .B0 (
                      scon_7), .B1 (nx1843)) ;
    INV_X0P5B_A12TS ix2290 (.Y (nx2289), .A (nx1879)) ;
    INV_X0P5B_A12TS ix1696 (.Y (nx1841), .A (nx2203)) ;
    INV_X0P5B_A12TS ix1698 (.Y (nx1833), .A (nx2220)) ;
    INV_X0P5B_A12TS ix1700 (.Y (nx1814), .A (nx2249)) ;
    INV_X0P5B_A12TS ix1702 (.Y (nx1904), .A (nx284)) ;
    INV_X0P5B_A12TS ix1703 (.Y (nx1813), .A (nx2254)) ;
    INV_X0P5B_A12TS ix2228 (.Y (nx2227), .A (nx1810)) ;
    INV_X0P5B_A12TS ix237 (.Y (nx236), .A (nx2373)) ;
    INV_X0P5B_A12TS ix1704 (.Y (nx1809), .A (nx2361)) ;
    INV_X0P5B_A12TS ix1705 (.Y (nx1806), .A (nx2310)) ;
    INV_X0P5B_A12TS ix2329 (.Y (nx2328), .A (nx158)) ;
    INV_X0P5B_A12TS ix1706 (.Y (nx1891), .A (nx1804)) ;
    INV_X0P5B_A12TS ix2417 (.Y (nx2416), .A (nx1801)) ;
    INV_X0P5B_A12TS ix1708 (.Y (nx2082), .A (nx2189)) ;
    OA21_X0P5M_A12TS ix1709 (.Y (nx1792), .A0 (prescaler_0), .A1 (prescaler_1), 
                     .B0 (nx1884)) ;
    NAND3B_X0P5M_A12TS ix2255 (.Y (nx2254), .AN (rd_addr_2), .B (rd_addr_0), .C (
                       rd_addr_1)) ;
    AND3_X0P5M_A12TS ix933 (.Y (nx932), .A (nx830), .B (nx158), .C (nx1801)) ;
    AND3_X0P5M_A12TS ix1710 (.Y (nx1845), .A (nx830), .B (nx1804), .C (nx1801)
                     ) ;
    NOR2B_X0P7M_A12TS ix1711 (.Y (nx1843), .AN (nx830), .B (nx2361)) ;
    OA21A1OI2_X0P5M_A12TS ix1929 (.Y (mulsrc2_2), .A0 (nx415), .A1 (nx433), .B0 (
                          nx435), .C0 (nx2091)) ;
    INV_X0P5B_A12TS ix416 (.Y (nx415), .A (tmp_mul_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_0 (.Q (tmp_mul_0), .CK (wb_clk_i), .D (
                       mulsrc2_0), .R (wb_rst_i)) ;
    AND2_X0P5M_A12TS ix1930 (.Y (mulsrc2_0), .A (src1_0), .B (nx42)) ;
    MXT4_X0P5M_A12TS ix43 (.Y (nx42), .A (src2_6), .B (src2_4), .C (src2_2), .D (
                     src2_0), .S0 (cycle_0), .S1 (cycle_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_cycle_0 (.Q (cycle_0), .CK (wb_clk_i), .D (
                        NOT_cycle_0), .R (wb_rst_i), .SE (NOT_enable), .SI (
                        cycle_0)) ;
    INV_X0P5B_A12TS ix426 (.Y (NOT_cycle_0), .A (cycle_0)) ;
    INV_X0P5B_A12TS ix1931 (.Y (NOT_enable), .A (enable_mul)) ;
    SDFFRPQ_X0P5M_A12TS reg_cycle_1 (.Q (cycle_1), .CK (wb_clk_i), .D (nx2085), 
                        .R (wb_rst_i), .SE (NOT_enable), .SI (cycle_1)) ;
    AOI21_X0P5M_A12TS ix1935 (.Y (nx2085), .A0 (cycle_0), .A1 (cycle_1), .B0 (
                      nx433)) ;
    NOR2_X0P5A_A12TS ix434 (.Y (nx433), .A (cycle_0), .B (cycle_1)) ;
    XNOR2_X0P5M_A12TS ix436 (.Y (nx435), .A (nx437), .B (nx2116)) ;
    NAND3_X0P5A_A12TS ix438 (.Y (nx437), .A (src1_1), .B (nx72), .C (mulsrc2_0)
                      ) ;
    MXT4_X0P5M_A12TS ix73 (.Y (nx72), .A (src2_7), .B (src2_5), .C (src2_3), .D (
                     src2_1), .S0 (cycle_0), .S1 (cycle_1)) ;
    XNOR2_X0P5M_A12TS ix1938 (.Y (nx2116), .A (nx2118), .B (nx444)) ;
    NAND2_X0P5A_A12TS ix1940 (.Y (nx2118), .A (src1_1), .B (nx72)) ;
    NAND2_X0P5A_A12TS ix1942 (.Y (nx444), .A (src1_2), .B (nx42)) ;
    NOR3_X0P5A_A12TS ix1943 (.Y (nx2091), .A (nx433), .B (nx415), .C (nx435)) ;
    AOI22_X0P5M_A12TS ix450 (.Y (nx449), .A0 (src1_0), .A1 (nx72), .B0 (src1_1)
                      , .B1 (nx42)) ;
    NAND4_X0P5A_A12TS ix433 (.Y (mulOv), .A (nx452), .B (nx609), .C (nx611), .D (
                      nx613)) ;
    NOR2_X0P5A_A12TS ix1945 (.Y (nx452), .A (mulsrc1_6), .B (mulsrc1_7)) ;
    OA21A1OI2_X0P5M_A12TS ix427 (.Y (mulsrc1_6), .A0 (nx2122), .A1 (nx433), .B0 (
                          nx2161), .C0 (nx2115)) ;
    INV_X0P5B_A12TS ix1947 (.Y (nx2122), .A (tmp_mul_12)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_12 (.Q (tmp_mul_12), .CK (wb_clk_i), .D (
                       mulsrc1_4), .R (wb_rst_i)) ;
    OA21A1OI2_X0P5M_A12TS ix1949 (.Y (mulsrc1_4), .A0 (nx459), .A1 (nx433), .B0 (
                          nx583), .C0 (nx374)) ;
    INV_X0P5B_A12TS ix460 (.Y (nx459), .A (tmp_mul_10)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_10 (.Q (tmp_mul_10), .CK (wb_clk_i), .D (
                       mulsrc1_2), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix367 (.Y (mulsrc1_2), .A (nx463)) ;
    AO21A1AI2_X0P5M_A12TS ix464 (.Y (nx463), .A0 (tmp_mul_8), .A1 (nx386), .B0 (
                          nx2110), .C0 (nx581)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_8 (.Q (tmp_mul_8), .CK (wb_clk_i), .D (
                       mulsrc1_0), .R (wb_rst_i)) ;
    XNOR2_X0P5M_A12TS ix1950 (.Y (mulsrc1_0), .A (nx2109), .B (nx556)) ;
    MXIT2_X0P5M_A12TS ix1952 (.Y (nx2109), .A (nx468), .B (nx2150), .S0 (nx2152)
                      ) ;
    MXIT2_X0P5M_A12TS ix1954 (.Y (nx468), .A (nx202), .B (nx2102), .S0 (nx524)
                      ) ;
    MXIT2_X0P5M_A12TS ix1955 (.Y (nx202), .A (nx2126), .B (nx2136), .S0 (nx510)
                      ) ;
    MXIT2_X0P5M_A12TS ix1956 (.Y (nx2126), .A (nx2096), .B (nx178), .S0 (nx495)
                      ) ;
    MXIT2_X0P5M_A12TS ix1957 (.Y (nx2096), .A (nx474), .B (nx480), .S0 (nx2093)
                      ) ;
    NAND2_X0P5A_A12TS ix475 (.Y (nx474), .A (tmp_mul_1), .B (nx386)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_1 (.Q (tmp_mul_1), .CK (wb_clk_i), .D (
                       mulsrc2_1), .R (wb_rst_i)) ;
    XNOR3_X0P5M_A12TS ix1958 (.Y (nx2093), .A (nx2127), .B (nx2129), .C (nx474)
                      ) ;
    OAI211_X0P5M_A12TS ix1960 (.Y (nx2127), .A0 (mulsrc2_0), .A1 (nx2087), .B0 (
                       src1_1), .C0 (nx72)) ;
    XNOR2_X0P5M_A12TS ix1961 (.Y (nx2129), .A (nx489), .B (nx2131)) ;
    NAND2_X0P5A_A12TS ix490 (.Y (nx489), .A (src1_2), .B (nx72)) ;
    NAND2_X0P5A_A12TS ix1962 (.Y (nx2131), .A (src1_3), .B (nx42)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_2 (.Q (tmp_mul_2), .CK (wb_clk_i), .D (
                       mulsrc2_2), .R (wb_rst_i)) ;
    XNOR3_X0P5M_A12TS ix496 (.Y (nx495), .A (nx146), .B (nx2132), .C (nx504)) ;
    CGENI_X1M_A12TS ix1963 (.CON (nx146), .A (nx2127), .B (nx489), .CI (nx2131)
                    ) ;
    XNOR2_X0P5M_A12TS ix1965 (.Y (nx2132), .A (nx500), .B (nx2135)) ;
    NAND2_X0P5A_A12TS ix1966 (.Y (nx500), .A (src1_3), .B (nx72)) ;
    NAND2_X0P5A_A12TS ix1967 (.Y (nx2135), .A (src1_4), .B (nx42)) ;
    NAND2_X0P5A_A12TS ix505 (.Y (nx504), .A (tmp_mul_2), .B (nx386)) ;
    NAND2_X0P5A_A12TS ix1968 (.Y (nx2136), .A (tmp_mul_3), .B (nx386)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_3 (.Q (tmp_mul_3), .CK (wb_clk_i), .D (
                       mulsrc2_3), .R (wb_rst_i)) ;
    XOR2_X0P5M_A12TS ix1970 (.Y (mulsrc2_3), .A (nx2091), .B (nx2093)) ;
    XNOR3_X0P5M_A12TS ix511 (.Y (nx510), .A (nx2095), .B (nx515), .C (nx2136)) ;
    CGENI_X1M_A12TS ix1972 (.CON (nx2095), .A (nx2138), .B (nx500), .CI (nx2135)
                    ) ;
    XNOR2_X0P5M_A12TS ix516 (.Y (nx515), .A (nx517), .B (nx519)) ;
    NAND2_X0P5A_A12TS ix518 (.Y (nx517), .A (src1_4), .B (nx72)) ;
    NAND2_X0P5A_A12TS ix520 (.Y (nx519), .A (src1_5), .B (nx42)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_4 (.Q (tmp_mul_4), .CK (wb_clk_i), .D (
                       mulsrc2_4), .R (wb_rst_i)) ;
    XNOR2_X0P5M_A12TS ix221 (.Y (mulsrc2_4), .A (nx2096), .B (nx495)) ;
    XNOR3_X0P5M_A12TS ix525 (.Y (nx524), .A (nx210), .B (nx2139), .C (nx2149)) ;
    CGENI_X1M_A12TS ix1974 (.CON (nx210), .A (nx527), .B (nx517), .CI (nx519)) ;
    XNOR2_X0P5M_A12TS ix1976 (.Y (nx2139), .A (nx2143), .B (nx2147)) ;
    NAND2_X0P5A_A12TS ix1978 (.Y (nx2143), .A (src1_5), .B (nx72)) ;
    NAND2_X0P5A_A12TS ix1980 (.Y (nx2147), .A (src1_6), .B (nx42)) ;
    NAND2_X0P5A_A12TS ix1981 (.Y (nx2149), .A (tmp_mul_4), .B (nx386)) ;
    NAND2_X0P5A_A12TS ix1983 (.Y (nx2150), .A (tmp_mul_5), .B (nx386)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_5 (.Q (tmp_mul_5), .CK (wb_clk_i), .D (
                       mulsrc2_5), .R (wb_rst_i)) ;
    XOR2_X0P5M_A12TS ix1985 (.Y (mulsrc2_5), .A (nx2126), .B (nx510)) ;
    XNOR3_X0P5M_A12TS ix1986 (.Y (nx2152), .A (nx2105), .B (nx2153), .C (nx2150)
                      ) ;
    CGENI_X1M_A12TS ix1988 (.CON (nx2105), .A (nx546), .B (nx2143), .CI (nx2147)
                    ) ;
    XNOR2_X0P5M_A12TS ix1990 (.Y (nx2153), .A (nx552), .B (nx2155)) ;
    NAND2_X0P5A_A12TS ix1991 (.Y (nx552), .A (src1_6), .B (nx72)) ;
    NAND2_X0P5A_A12TS ix1994 (.Y (nx2155), .A (src1_7), .B (nx42)) ;
    XNOR2_X0P5M_A12TS ix557 (.Y (nx556), .A (nx558), .B (nx2156)) ;
    AO21A1AI2_X0P5M_A12TS ix559 (.Y (nx558), .A0 (src1_7), .A1 (nx72), .B0 (
                          nx2106), .C0 (nx565)) ;
    CGENI_X1M_A12TS ix1997 (.CON (nx2106), .A (nx561), .B (nx552), .CI (nx2155)
                    ) ;
    NAND3_X0P5A_A12TS ix566 (.Y (nx565), .A (nx2106), .B (src1_7), .C (nx72)) ;
    NAND2_X0P5A_A12TS ix1999 (.Y (nx2156), .A (tmp_mul_6), .B (nx386)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_6 (.Q (tmp_mul_6), .CK (wb_clk_i), .D (
                       mulsrc2_6), .R (wb_rst_i)) ;
    XNOR2_X0P5M_A12TS ix2000 (.Y (mulsrc2_6), .A (nx202), .B (nx524)) ;
    MXIT2_X0P5M_A12TS ix2008 (.Y (nx2110), .A (nx2159), .B (nx2160), .S0 (nx579)
                      ) ;
    MXIT2_X0P5M_A12TS ix2010 (.Y (nx2159), .A (nx2109), .B (nx2104), .S0 (nx556)
                      ) ;
    NAND2_X0P5A_A12TS ix2012 (.Y (nx2160), .A (tmp_mul_7), .B (nx386)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_7 (.Q (tmp_mul_7), .CK (wb_clk_i), .D (
                       mulsrc2_7), .R (wb_rst_i)) ;
    XOR2_X0P5M_A12TS ix311 (.Y (mulsrc2_7), .A (nx468), .B (nx2152)) ;
    XNOR2_X0P5M_A12TS ix580 (.Y (nx579), .A (nx565), .B (nx2160)) ;
    NAND3_X0P5A_A12TS ix582 (.Y (nx581), .A (nx386), .B (tmp_mul_8), .C (nx2110)
                      ) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_9 (.Q (tmp_mul_9), .CK (wb_clk_i), .D (
                       mulsrc1_1), .R (wb_rst_i)) ;
    XOR2_X0P5M_A12TS ix321 (.Y (mulsrc1_1), .A (nx2159), .B (nx579)) ;
    NAND3_X0P5A_A12TS ix2013 (.Y (nx2161), .A (nx386), .B (tmp_mul_11), .C (
                      nx374)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_11 (.Q (tmp_mul_11), .CK (wb_clk_i), .D (
                       mulsrc1_3), .R (wb_rst_i)) ;
    OA21A1OI2_X0P5M_A12TS ix2015 (.Y (mulsrc1_3), .A0 (nx593), .A1 (nx433), .B0 (
                          nx581), .C0 (nx2112)) ;
    INV_X0P5B_A12TS ix594 (.Y (nx593), .A (tmp_mul_9)) ;
    XOR2_X0P5M_A12TS ix419 (.Y (mulsrc1_7), .A (nx2163), .B (nx2167)) ;
    NAND3_X0P5A_A12TS ix2019 (.Y (nx2163), .A (nx386), .B (tmp_mul_12), .C (
                      nx2113)) ;
    INV_X0P5B_A12TS ix602 (.Y (nx601), .A (tmp_mul_11)) ;
    NAND3_X0P5A_A12TS ix2023 (.Y (nx2165), .A (nx386), .B (tmp_mul_10), .C (
                      nx2112)) ;
    NAND2_X0P5A_A12TS ix2026 (.Y (nx2167), .A (tmp_mul_13), .B (nx386)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_mul_13 (.Q (tmp_mul_13), .CK (wb_clk_i), .D (
                       mulsrc1_5), .R (wb_rst_i)) ;
    OA21A1OI2_X0P5M_A12TS ix387 (.Y (mulsrc1_5), .A0 (nx601), .A1 (nx433), .B0 (
                          nx2165), .C0 (nx2113)) ;
    NOR2_X0P5A_A12TS ix610 (.Y (nx609), .A (mulsrc1_0), .B (mulsrc1_1)) ;
    NOR2_X0P5A_A12TS ix612 (.Y (nx611), .A (mulsrc1_2), .B (mulsrc1_3)) ;
    NOR2_X0P5A_A12TS ix614 (.Y (nx613), .A (mulsrc1_4), .B (mulsrc1_5)) ;
    INV_X0P5B_A12TS ix2028 (.Y (nx2115), .A (nx2163)) ;
    INV_X0P5B_A12TS ix2031 (.Y (nx2113), .A (nx2161)) ;
    INV_X0P5B_A12TS ix375 (.Y (nx374), .A (nx2165)) ;
    INV_X0P5B_A12TS ix2035 (.Y (nx2112), .A (nx583)) ;
    INV_X0P5B_A12TS ix562 (.Y (nx561), .A (nx2105)) ;
    INV_X0P5B_A12TS ix2038 (.Y (nx2104), .A (nx2156)) ;
    INV_X0P5B_A12TS ix2040 (.Y (nx2102), .A (nx2149)) ;
    INV_X0P5B_A12TS ix547 (.Y (nx546), .A (nx210)) ;
    INV_X0P5B_A12TS ix179 (.Y (nx178), .A (nx504)) ;
    INV_X0P5B_A12TS ix528 (.Y (nx527), .A (nx2095)) ;
    INV_X0P5B_A12TS ix2042 (.Y (nx2138), .A (nx146)) ;
    INV_X0P5B_A12TS ix481 (.Y (nx480), .A (nx2091)) ;
    INV_X0P5B_A12TS ix2045 (.Y (nx2087), .A (nx444)) ;
    INV_X0P5B_A12TS ix2048 (.Y (nx386), .A (nx433)) ;
    NOR2B_X0P7M_A12TS ix113 (.Y (mulsrc2_1), .AN (nx437), .B (nx449)) ;
    NAND3B_X0P5M_A12TS ix584 (.Y (nx583), .AN (nx581), .B (nx386), .C (tmp_mul_9
                       )) ;
    NOR2_X0P5A_A12TS ix2168 (.Y (divOv), .A (nx2406), .B (nx2408)) ;
    NOR2_X0P5A_A12TS ix2170 (.Y (divsrc2_0), .A (nx801), .B (nx826)) ;
    OA21A1OI2_X0P5M_A12TS ix802 (.Y (nx801), .A0 (nx2355), .A1 (
                          cycle_0__dup_2349), .B0 (cycle_1__dup_2348), .C0 (
                          nx104)) ;
    NOR2_X0P5A_A12TS ix2171 (.Y (nx2355), .A (src2_7), .B (src2_6)) ;
    DFFRPQ_X0P5M_A12TS reg_cycle_0__dup_66619 (.Q (cycle_0__dup_2349), .CK (
                       wb_clk_i), .D (nx759), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix760 (.Y (nx759), .A0 (nx2410), .A1 (enable_div), .B0 (
                      nx808)) ;
    INV_X0P5B_A12TS ix2175 (.Y (nx2410), .A (cycle_0__dup_2349)) ;
    NAND2_X0P5A_A12TS ix809 (.Y (nx808), .A (nx2410), .B (enable_div)) ;
    DFFRPQ_X0P5M_A12TS reg_cycle_1__dup_66623 (.Q (cycle_1__dup_2348), .CK (
                       wb_clk_i), .D (nx769), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix770 (.Y (nx769), .A0 (nx812), .A1 (enable_div), .B0 (
                      nx2411)) ;
    INV_X0P5B_A12TS ix813 (.Y (nx812), .A (cycle_1__dup_2348)) ;
    NAND3_X0P5A_A12TS ix2179 (.Y (nx2411), .A (nx2351), .B (nx730), .C (
                      enable_div)) ;
    NAND2_X0P5A_A12TS ix2181 (.Y (nx730), .A (cycle_0__dup_2349), .B (
                      cycle_1__dup_2348)) ;
    AND4_X0P5M_A12TS ix2182 (.Y (nx104), .A (nx819), .B (nx821), .C (nx823), .D (
                     nx2353)) ;
    MXIT2_X0P5M_A12TS ix820 (.Y (nx819), .A (src2_4), .B (src2_6), .S0 (
                      cycle_0__dup_2349)) ;
    MXIT2_X0P5M_A12TS ix822 (.Y (nx821), .A (src2_3), .B (src2_5), .S0 (
                      cycle_0__dup_2349)) ;
    MXIT2_X0P5M_A12TS ix824 (.Y (nx823), .A (src2_2), .B (src2_4), .S0 (
                      cycle_0__dup_2349)) ;
    OA21A1OI2_X0P5M_A12TS ix2183 (.Y (nx2353), .A0 (src2_5), .A1 (src2_6), .B0 (
                          nx2410), .C0 (src2_7)) ;
    MXIT2_X0P5M_A12TS ix827 (.Y (nx826), .A (nx2400), .B (nx2444), .S0 (nx2437)
                      ) ;
    MXIT2_X0P5M_A12TS ix2186 (.Y (nx2400), .A (nx829), .B (nx2362), .S0 (nx966)
                      ) ;
    MXIT2_X0P5M_A12TS ix830 (.Y (nx829), .A (nx2386), .B (nx950), .S0 (nx2423)
                      ) ;
    MXIT2_X0P5M_A12TS ix2192 (.Y (nx2386), .A (nx832), .B (nx2369), .S0 (nx929)
                      ) ;
    MXIT2_X0P5M_A12TS ix833 (.Y (nx832), .A (nx426), .B (nx2442), .S0 (nx2419)
                      ) ;
    MXIT2_X0P5M_A12TS ix2195 (.Y (nx426), .A (nx835), .B (nx214), .S0 (nx890)) ;
    MXIT2_X0P5M_A12TS ix836 (.Y (nx835), .A (nx739), .B (nx849), .S0 (nx851)) ;
    NAND4B_X0P5M_A12TS ix269 (.Y (nx739), .AN (tmp_rem_0), .B (cycle_0__dup_2349
                       ), .C (cycle_1__dup_2348), .D (src2_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_0 (.Q (tmp_rem_0), .CK (wb_clk_i), .D (
                       divsrc1_0), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix257 (.Y (divsrc1_0), .A0 (divsrc2_0), .A1 (nx238), .B0 (
                          nx841), .C0 (nx843)) ;
    AOI32_X0P5M_A12TS ix2197 (.Y (nx841), .A0 (src1_0), .A1 (nx2410), .A2 (nx812
                      ), .B0 (tmp_rem_0), .B1 (nx2351)) ;
    NAND3_X0P5A_A12TS ix2198 (.Y (nx849), .A (src2_1), .B (cycle_0__dup_2349), .C (
                      cycle_1__dup_2348)) ;
    XOR2_X0P5M_A12TS ix2200 (.Y (nx851), .A (nx849), .B (nx853)) ;
    AOI21_X0P5M_A12TS ix2201 (.Y (nx853), .A0 (nx855), .A1 (divsrc2_1), .B0 (
                      nx2376)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_1 (.Q (tmp_rem_1), .CK (wb_clk_i), .D (
                       divsrc1_1), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2206 (.Y (divsrc1_1), .A0 (nx853), .A1 (divsrc2_0), .B0 (
                      nx861)) ;
    NAND2_X0P5A_A12TS ix2207 (.Y (nx861), .A (divsrc2_0), .B (nx2372)) ;
    XNOR2_X0P5M_A12TS ix2212 (.Y (nx2372), .A (nx739), .B (nx851)) ;
    NOR3_X0P5A_A12TS ix2214 (.Y (divsrc2_1), .A (nx865), .B (nx2358), .C (nx801)
                     ) ;
    CGENI_X1M_A12TS ix2216 (.CON (nx354), .A (nx2413), .B (nx953), .CI (nx2365)
                    ) ;
    CGENI_X1M_A12TS ix2217 (.CON (nx2413), .A (nx2374), .B (nx743), .CI (nx931)
                    ) ;
    CGENI_X1M_A12TS ix2219 (.CON (nx2374), .A (nx871), .B (nx915), .CI (nx2371)
                    ) ;
    CGENI_X1M_A12TS ix2220 (.CON (nx873), .A (nx334), .B (nx746), .CI (nx849)) ;
    NAND4B_X0P5M_A12TS ix335 (.Y (nx334), .AN (tmp_rem_1), .B (src2_0), .C (
                       cycle_0__dup_2349), .D (cycle_1__dup_2348)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_2 (.Q (tmp_rem_2), .CK (wb_clk_i), .D (
                       divsrc1_2), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2222 (.Y (divsrc1_2), .A0 (nx879), .A1 (divsrc2_0), .B0 (
                      nx887)) ;
    AOI21_X0P5M_A12TS ix2224 (.Y (nx879), .A0 (divsrc2_1), .A1 (nx2381), .B0 (
                      nx2379)) ;
    XNOR2_X0P5M_A12TS ix2225 (.Y (nx2381), .A (nx334), .B (nx2415)) ;
    XOR2_X0P5M_A12TS ix2226 (.Y (nx2415), .A (nx884), .B (nx849)) ;
    AOI32_X0P5M_A12TS ix2227 (.Y (nx884), .A0 (src1_2), .A1 (nx2410), .A2 (nx812
                      ), .B0 (tmp_rem_2), .B1 (nx2351)) ;
    NOR2_X0P5A_A12TS ix2229 (.Y (nx2379), .A (nx884), .B (divsrc2_1)) ;
    NAND2_X0P5A_A12TS ix2230 (.Y (nx887), .A (divsrc2_0), .B (nx2377)) ;
    XOR2_X0P5M_A12TS ix2231 (.Y (nx2377), .A (nx835), .B (nx890)) ;
    XNOR2_X0P5M_A12TS ix2234 (.Y (nx890), .A (nx214), .B (nx879)) ;
    NOR2_X0P5A_A12TS ix215 (.Y (nx214), .A (nx812), .B (nx893)) ;
    MXIT2_X0P5M_A12TS ix2236 (.Y (nx893), .A (src2_0), .B (src2_2), .S0 (
                      cycle_0__dup_2349)) ;
    NOR2_X0P5A_A12TS ix2238 (.Y (nx895), .A (cycle_0__dup_2349), .B (
                     cycle_1__dup_2348)) ;
    AOI32_X0P5M_A12TS ix2240 (.Y (nx897), .A0 (src1_3), .A1 (nx2410), .A2 (nx812
                      ), .B0 (tmp_rem_3), .B1 (nx2351)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_3 (.Q (tmp_rem_3), .CK (wb_clk_i), .D (
                       divsrc1_3), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2241 (.Y (divsrc1_3), .A0 (nx901), .A1 (divsrc2_0), .B0 (
                      nx907)) ;
    AOI21_X0P5M_A12TS ix2242 (.Y (nx901), .A0 (divsrc2_1), .A1 (nx446), .B0 (
                      nx2382)) ;
    XOR2_X0P5M_A12TS ix447 (.Y (nx446), .A (nx873), .B (nx2417)) ;
    XNOR2_X0P5M_A12TS ix2243 (.Y (nx2417), .A (nx897), .B (nx214)) ;
    NOR2_X0P5A_A12TS ix2247 (.Y (nx2382), .A (nx897), .B (divsrc2_1)) ;
    NAND2_X0P5A_A12TS ix908 (.Y (nx907), .A (divsrc2_0), .B (nx428)) ;
    XNOR2_X0P5M_A12TS ix429 (.Y (nx428), .A (nx426), .B (nx2419)) ;
    XNOR2_X0P5M_A12TS ix2249 (.Y (nx2419), .A (nx2371), .B (nx901)) ;
    NOR2_X0P5A_A12TS ix2253 (.Y (nx2371), .A (nx812), .B (nx913)) ;
    MXIT2_X0P5M_A12TS ix914 (.Y (nx913), .A (src2_1), .B (src2_3), .S0 (
                      cycle_0__dup_2349)) ;
    AOI32_X0P5M_A12TS ix916 (.Y (nx915), .A0 (src1_4), .A1 (nx2410), .A2 (nx812)
                      , .B0 (tmp_rem_4), .B1 (nx2351)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_4 (.Q (tmp_rem_4), .CK (wb_clk_i), .D (
                       divsrc1_4), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2254 (.Y (divsrc1_4), .A0 (nx919), .A1 (divsrc2_0), .B0 (
                      nx926)) ;
    AOI21_X0P5M_A12TS ix920 (.Y (nx919), .A0 (divsrc2_1), .A1 (nx482), .B0 (
                      nx2384)) ;
    XNOR2_X0P5M_A12TS ix483 (.Y (nx482), .A (nx342), .B (nx923)) ;
    CGENI_X1M_A12TS ix2256 (.CON (nx342), .A (nx873), .B (nx897), .CI (nx214)) ;
    XNOR2_X0P5M_A12TS ix924 (.Y (nx923), .A (nx915), .B (nx2371)) ;
    NOR2_X0P5A_A12TS ix2258 (.Y (nx2384), .A (nx915), .B (divsrc2_1)) ;
    NAND2_X0P5A_A12TS ix927 (.Y (nx926), .A (divsrc2_0), .B (nx464)) ;
    XOR2_X0P5M_A12TS ix2259 (.Y (nx464), .A (nx832), .B (nx929)) ;
    XOR2_X0P5M_A12TS ix930 (.Y (nx929), .A (nx931), .B (nx919)) ;
    AOI31_X0P5M_A12TS ix932 (.Y (nx931), .A0 (cycle_0__dup_2349), .A1 (src2_0), 
                      .A2 (nx812), .B0 (nx2367)) ;
    NOR2_X0P5A_A12TS ix2261 (.Y (nx2367), .A (nx812), .B (nx823)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_5 (.Q (tmp_rem_5), .CK (wb_clk_i), .D (
                       divsrc1_5), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2263 (.Y (divsrc1_5), .A0 (nx937), .A1 (divsrc2_0), .B0 (
                      nx945)) ;
    AOI21_X0P5M_A12TS ix938 (.Y (nx937), .A0 (divsrc2_1), .A1 (nx2393), .B0 (
                      nx2392)) ;
    XNOR2_X0P5M_A12TS ix2265 (.Y (nx2393), .A (nx2374), .B (nx940)) ;
    XOR2_X0P5M_A12TS ix941 (.Y (nx940), .A (nx2421), .B (nx931)) ;
    AOI32_X0P5M_A12TS ix2267 (.Y (nx2421), .A0 (src1_5), .A1 (nx2410), .A2 (
                      nx812), .B0 (tmp_rem_5), .B1 (nx2351)) ;
    NOR2_X0P5A_A12TS ix2268 (.Y (nx2392), .A (nx2421), .B (divsrc2_1)) ;
    NAND2_X0P5A_A12TS ix946 (.Y (nx945), .A (divsrc2_0), .B (nx2390)) ;
    XNOR2_X0P5M_A12TS ix2270 (.Y (nx2390), .A (nx2386), .B (nx2423)) ;
    XOR2_X0P5M_A12TS ix2272 (.Y (nx2423), .A (nx950), .B (nx937)) ;
    AOI31_X0P5M_A12TS ix951 (.Y (nx950), .A0 (cycle_0__dup_2349), .A1 (src2_1), 
                      .A2 (nx812), .B0 (nx2364)) ;
    NOR2_X0P5A_A12TS ix2274 (.Y (nx2364), .A (nx812), .B (nx821)) ;
    AOI32_X0P5M_A12TS ix954 (.Y (nx953), .A0 (src1_6), .A1 (nx2410), .A2 (nx812)
                      , .B0 (tmp_rem_6), .B1 (nx2351)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_6 (.Q (tmp_rem_6), .CK (wb_clk_i), .D (
                       divsrc1_6), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix541 (.Y (divsrc1_6), .A0 (nx957), .A1 (divsrc2_0), .B0 (
                      nx963)) ;
    AOI21_X0P5M_A12TS ix958 (.Y (nx957), .A0 (divsrc2_1), .A1 (nx2399), .B0 (
                      nx2397)) ;
    XOR2_X0P5M_A12TS ix2276 (.Y (nx2399), .A (nx2413), .B (nx2424)) ;
    XOR2_X0P5M_A12TS ix2278 (.Y (nx2424), .A (nx953), .B (nx950)) ;
    NOR2_X0P5A_A12TS ix2279 (.Y (nx2397), .A (nx953), .B (divsrc2_1)) ;
    NAND2_X0P5A_A12TS ix964 (.Y (nx963), .A (divsrc2_0), .B (nx2395)) ;
    XOR2_X0P5M_A12TS ix2281 (.Y (nx2395), .A (nx829), .B (nx966)) ;
    XNOR2_X0P5M_A12TS ix967 (.Y (nx966), .A (nx2362), .B (nx957)) ;
    MXIT2_X0P5M_A12TS ix2282 (.Y (nx2362), .A (nx893), .B (nx819), .S0 (
                      cycle_1__dup_2348)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_rem_7 (.Q (tmp_rem_7), .CK (wb_clk_i), .D (
                       divsrc1_7), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix2284 (.Y (divsrc1_7), .A0 (nx2428), .A1 (divsrc2_0), .B0 (
                      nx2435)) ;
    AOI21_X0P5M_A12TS ix976 (.Y (nx2428), .A0 (nx590), .A1 (divsrc2_1), .B0 (
                      nx2404)) ;
    XNOR2_X0P5M_A12TS ix591 (.Y (nx590), .A (nx354), .B (nx2432)) ;
    XNOR2_X0P5M_A12TS ix2286 (.Y (nx2432), .A (nx2433), .B (nx2362)) ;
    AOI32_X0P5M_A12TS ix2288 (.Y (nx2433), .A0 (src1_7), .A1 (nx2410), .A2 (
                      nx812), .B0 (tmp_rem_7), .B1 (nx2351)) ;
    NOR2_X0P5A_A12TS ix2289 (.Y (nx2404), .A (nx2433), .B (divsrc2_1)) ;
    NAND2_X0P5A_A12TS ix984 (.Y (nx2435), .A (nx2402), .B (divsrc2_0)) ;
    XNOR2_X0P5M_A12TS ix2291 (.Y (nx2402), .A (nx2400), .B (nx2437)) ;
    XNOR2_X0P5M_A12TS ix987 (.Y (nx2437), .A (nx2358), .B (nx2428)) ;
    MXIT2_X0P5M_A12TS ix2292 (.Y (nx2358), .A (nx913), .B (nx2439), .S0 (
                      cycle_1__dup_2348)) ;
    MXIT2_X0P5M_A12TS ix990 (.Y (nx2439), .A (src2_5), .B (src2_7), .S0 (
                      cycle_0__dup_2349)) ;
    AOI21_X0P5M_A12TS ix2296 (.Y (nx2376), .A0 (divsrc2_1), .A1 (nx238), .B0 (
                      nx2440)) ;
    AOI32_X0P5M_A12TS ix999 (.Y (nx2440), .A0 (src1_1), .A1 (nx2410), .A2 (nx812
                      ), .B0 (tmp_rem_1), .B1 (nx2351)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_div_0 (.Q (divsrc2_2), .CK (wb_clk_i), .D (
                       divsrc2_0), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_div_1 (.Q (divsrc2_3), .CK (wb_clk_i), .D (
                       divsrc2_1), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_div_2 (.Q (divsrc2_4), .CK (wb_clk_i), .D (
                       divsrc2_2), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_div_3 (.Q (divsrc2_5), .CK (wb_clk_i), .D (
                       divsrc2_3), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_div_4 (.Q (divsrc2_6), .CK (wb_clk_i), .D (
                       divsrc2_4), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tmp_div_5 (.Q (divsrc2_7), .CK (wb_clk_i), .D (
                       divsrc2_5), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix2298 (.Y (nx871), .A (nx342)) ;
    INV_X0P5B_A12TS ix2299 (.Y (nx855), .A (nx334)) ;
    INV_X0P5B_A12TS ix405 (.Y (nx746), .A (nx884)) ;
    INV_X0P5B_A12TS ix513 (.Y (nx743), .A (nx2421)) ;
    INV_X0P5B_A12TS ix1001 (.Y (nx2442), .A (nx2371)) ;
    INV_X0P5B_A12TS ix2300 (.Y (nx2369), .A (nx931)) ;
    INV_X0P5B_A12TS ix2302 (.Y (nx2365), .A (nx950)) ;
    INV_X0P5B_A12TS ix2303 (.Y (nx2444), .A (nx2358)) ;
    INV_X0P5B_A12TS ix2306 (.Y (nx2351), .A (nx895)) ;
    OR4_X0P5M_A12TS ix2308 (.Y (nx2406), .A (src2_7), .B (src2_6), .C (src2_5), 
                    .D (src2_4)) ;
    OR4_X0P5M_A12TS ix2309 (.Y (nx2408), .A (src2_3), .B (src2_2), .C (src2_1), 
                    .D (src2_0)) ;
    NOR2B_X0P7M_A12TS ix239 (.Y (nx238), .AN (src2_0), .B (nx730)) ;
    NAND2B_X0P7M_A12TS ix2310 (.Y (nx843), .AN (nx739), .B (divsrc2_0)) ;
    CGEN_X1M_A12TS ix2312 (.CO (nx865), .A (nx1025), .B (nx2433), .CI (nx2362)
                   ) ;
    INV_X0P5B_A12TS ix2314 (.Y (nx1025), .A (nx354)) ;
    NAND4_X0P5A_A12TS ix2445 (.Y (nx3225), .A (wr_addr_m_0), .B (wr_addr_m_1), .C (
                      wr_addr_m_2), .D (wr_addr_m_3)) ;
    INV_X4M_A12TS ix2449 (.Y (nx3286), .A (wr_dup_1054)) ;
    NAND4_X0P5A_A12TS ix5443 (.Y (nx5442), .A (wr_addr_m_4), .B (wr_addr_m_5), .C (
                      wr_addr_m_6), .D (wr_addr_7)) ;
    NAND3_X0P5A_A12TS ix2450 (.Y (nx3224), .A (nx3287), .B (wr_addr_m_2), .C (
                      wr_addr_m_3)) ;
    NAND3_X0P5A_A12TS ix391 (.Y (nx390), .A (nx443), .B (wr_addr_m_2), .C (
                      wr_addr_m_3)) ;
    NAND3_X0P5A_A12TS ix2452 (.Y (nx3223), .A (nx3288), .B (wr_addr_m_2), .C (
                      wr_addr_m_3)) ;
    NOR2_X0P5A_A12TS ix2454 (.Y (nx3288), .A (wr_addr_m_0), .B (wr_addr_m_1)) ;
    NAND3_X0P5A_A12TS ix337 (.Y (nx336), .A (nx3289), .B (wr_addr_m_0), .C (
                      wr_addr_m_1)) ;
    NAND2_X0P5A_A12TS ix2457 (.Y (nx316), .A (nx3289), .B (nx3287)) ;
    NAND2_X0P5A_A12TS ix293 (.Y (nx292), .A (nx3289), .B (nx443)) ;
    NAND2_X0P5A_A12TS ix2458 (.Y (nx3220), .A (nx3289), .B (nx3288)) ;
    NAND3_X0P5A_A12TS ix2460 (.Y (nx3218), .A (nx3290), .B (wr_addr_m_0), .C (
                      wr_addr_m_1)) ;
    NAND2_X0P5A_A12TS ix2462 (.Y (nx3217), .A (nx3290), .B (nx3287)) ;
    NAND2_X0P5A_A12TS ix2464 (.Y (nx3216), .A (nx3290), .B (nx443)) ;
    NAND2_X0P5A_A12TS ix2467 (.Y (nx172), .A (nx3290), .B (nx3288)) ;
    NAND3_X0P5A_A12TS ix2469 (.Y (nx140), .A (nx490), .B (wr_addr_m_0), .C (
                      wr_addr_m_1)) ;
    NOR2_X0P5A_A12TS ix491 (.Y (nx490), .A (wr_addr_m_2), .B (wr_addr_m_3)) ;
    NAND2_X0P5A_A12TS ix2470 (.Y (nx3215), .A (nx490), .B (nx3287)) ;
    NAND2_X0P5A_A12TS ix2471 (.Y (nx3214), .A (nx490), .B (nx443)) ;
    NAND2_X0P5A_A12TS ix63 (.Y (nx62), .A (nx490), .B (nx3288)) ;
    NAND3_X0P5A_A12TS ix5093 (.Y (nx5092), .A (nx503), .B (wr_addr_m_6), .C (
                      wr_addr_7)) ;
    NAND3_X0P5A_A12TS ix4739 (.Y (nx4738), .A (nx529), .B (wr_addr_m_6), .C (
                      wr_addr_7)) ;
    NAND3_X0P5A_A12TS ix2473 (.Y (nx3263), .A (nx557), .B (wr_addr_m_6), .C (
                      wr_addr_7)) ;
    NOR2_X0P5A_A12TS ix558 (.Y (nx557), .A (wr_addr_m_4), .B (wr_addr_m_5)) ;
    NAND3_X0P5A_A12TS ix4025 (.Y (nx4024), .A (nx3291), .B (wr_addr_m_4), .C (
                      wr_addr_m_5)) ;
    NAND2_X0P5A_A12TS ix3675 (.Y (nx3674), .A (nx3291), .B (nx503)) ;
    NAND2_X0P5A_A12TS ix3321 (.Y (nx3320), .A (nx3291), .B (nx529)) ;
    NAND2_X0P5A_A12TS ix2971 (.Y (nx2970), .A (nx3291), .B (nx557)) ;
    NAND3_X0P5A_A12TS ix2474 (.Y (nx3257), .A (nx673), .B (wr_addr_m_4), .C (
                      wr_addr_m_5)) ;
    NAND2_X0P5A_A12TS ix2475 (.Y (nx3250), .A (nx673), .B (nx503)) ;
    NAND2_X0P5A_A12TS ix2476 (.Y (nx3247), .A (nx673), .B (nx529)) ;
    NAND2_X0P5A_A12TS ix2477 (.Y (nx1550), .A (nx673), .B (nx557)) ;
    NAND3_X0P5A_A12TS ix2478 (.Y (nx3239), .A (nx763), .B (wr_addr_m_4), .C (
                      wr_addr_m_5)) ;
    NOR2_X0P5A_A12TS ix764 (.Y (nx763), .A (wr_addr_m_6), .B (wr_addr_7)) ;
    NAND2_X0P5A_A12TS ix2480 (.Y (nx3231), .A (nx763), .B (nx503)) ;
    NAND2_X0P5A_A12TS ix2481 (.Y (nx3227), .A (nx763), .B (nx529)) ;
    NAND2_X0P5A_A12TS ix2483 (.Y (nx3213), .A (nx763), .B (nx557)) ;
    TIELO_X1M_A12TS ix2484 (.Y (nx3204)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_0 (.Q (rd_data_m_0), .CK (wb_clk_i), .D (
                        nx5810), .R (wb_rst_i), .SE (NOT_nx50), .SI (rd_data_m_0
                        )) ;
    MXIT2_X0P5M_A12TS ix5811 (.Y (nx5810), .A (nx863), .B (nx3292), .S0 (nx1127)
                      ) ;
    INV_X0P5B_A12TS ix2486 (.Y (nx863), .A (wr_data_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2488 (.Y (nx3292), .A0 (nx5796), .A1 (nx4380), .B0 (
                          rd_addr_7), .C0 (nx2964)) ;
    OA21A1OI2_X0P5M_A12TS ix5797 (.Y (nx5796), .A0 (rd_addr_m_5), .A1 (nx869), .B0 (
                          nx3298), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2490 (.Y (nx869), .A0 (rd_addr_m_4), .A1 (nx5082), .B0 (
                      nx4736)) ;
    MXT4_X0P5M_A12TS ix5083 (.Y (nx5082), .A (nx4818), .B (nx4990), .C (nx4902)
                     , .D (nx5074), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix4819 (.Y (nx4818), .A (modgen_ram_ix167_a_208__dup_2445)
                     , .B (modgen_ram_ix167_a_210__dup_2443), .C (
                     modgen_ram_ix167_a_209__dup_2444), .D (
                     modgen_ram_ix167_a_211__dup_2442), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix4991 (.Y (nx4990), .A (modgen_ram_ix167_a_216__dup_2437)
                     , .B (modgen_ram_ix167_a_218__dup_2435), .C (
                     modgen_ram_ix167_a_217__dup_2436), .D (
                     modgen_ram_ix167_a_219__dup_2434), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix4903 (.Y (nx4902), .A (modgen_ram_ix167_a_212__dup_2441)
                     , .B (modgen_ram_ix167_a_214__dup_2439), .C (
                     modgen_ram_ix167_a_213__dup_2440), .D (
                     modgen_ram_ix167_a_215__dup_2438), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix5075 (.Y (nx5074), .A (modgen_ram_ix167_a_220__dup_2433)
                     , .B (modgen_ram_ix167_a_222__dup_2431), .C (
                     modgen_ram_ix167_a_221__dup_2432), .D (
                     modgen_ram_ix167_a_223__dup_2430), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix4737 (.Y (nx4736), .A0 (rd_addr_m_3), .A1 (nx3293), 
                          .B0 (nx889), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2492 (.Y (nx3293), .A0 (rd_addr_m_2), .A1 (nx4552), .B0 (
                      nx4472)) ;
    MXT4_X0P5M_A12TS ix4553 (.Y (nx4552), .A (modgen_ram_ix167_a_196__dup_2457)
                     , .B (modgen_ram_ix167_a_198__dup_2455), .C (
                     modgen_ram_ix167_a_197__dup_2456), .D (
                     modgen_ram_ix167_a_199__dup_2454), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix4473 (.Y (nx4472), .A0 (rd_addr_m_1), .A1 (nx3294), 
                          .B0 (nx886), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2493 (.Y (nx3294), .A (modgen_ram_ix167_a_192__dup_2461)
                      , .B (modgen_ram_ix167_a_193__dup_2460), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2494 (.Y (nx886), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_2458), .B0 (nx3264), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2495 (.Y (nx3264), .AN (modgen_ram_ix167_a_194__dup_2459
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2497 (.Y (nx889), .A0 (rd_addr_m_2), .A1 (nx4724), .B0 (
                          nx4644), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix4725 (.Y (nx4724), .A (modgen_ram_ix167_a_204__dup_2449)
                     , .B (modgen_ram_ix167_a_206__dup_2447), .C (
                     modgen_ram_ix167_a_205__dup_2448), .D (
                     modgen_ram_ix167_a_207__dup_2446), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix4645 (.Y (nx4644), .A0 (rd_addr_m_1), .A1 (nx3295), 
                          .B0 (nx3297), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2498 (.Y (nx3295), .A (modgen_ram_ix167_a_200__dup_2453)
                      , .B (modgen_ram_ix167_a_201__dup_2452), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2499 (.Y (nx3297), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_2450), .B0 (nx4618), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix4619 (.Y (nx4618), .AN (modgen_ram_ix167_a_202__dup_2451
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2502 (.Y (nx3298), .A0 (rd_addr_m_4), .A1 (nx5786), 
                          .B0 (nx5440), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix5787 (.Y (nx5786), .A (nx5522), .B (nx3265), .C (nx5606)
                     , .D (nx5778), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix5523 (.Y (nx5522), .A (modgen_ram_ix167_a_240__dup_2413)
                     , .B (modgen_ram_ix167_a_242__dup_2411), .C (
                     modgen_ram_ix167_a_241__dup_2412), .D (
                     modgen_ram_ix167_a_243__dup_2410), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2504 (.Y (nx3265), .A (modgen_ram_ix167_a_248__dup_2405)
                     , .B (modgen_ram_ix167_a_250__dup_2403), .C (
                     modgen_ram_ix167_a_249__dup_2404), .D (
                     modgen_ram_ix167_a_251__dup_2402), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix5607 (.Y (nx5606), .A (modgen_ram_ix167_a_244__dup_2409)
                     , .B (modgen_ram_ix167_a_246__dup_2407), .C (
                     modgen_ram_ix167_a_245__dup_2408), .D (
                     modgen_ram_ix167_a_247__dup_2406), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix5779 (.Y (nx5778), .A (modgen_ram_ix167_a_252__dup_2401)
                     , .B (modgen_ram_ix167_a_254__dup_2399), .C (
                     modgen_ram_ix167_a_253__dup_2400), .D (
                     modgen_ram_ix167_a_255__dup_2398), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix5441 (.Y (nx5440), .A0 (rd_addr_m_3), .A1 (nx911), .B0 (
                          nx3300), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix912 (.Y (nx911), .A0 (rd_addr_m_2), .A1 (nx5256), .B0 (
                      nx5176)) ;
    MXT4_X0P5M_A12TS ix5257 (.Y (nx5256), .A (modgen_ram_ix167_a_228__dup_2425)
                     , .B (modgen_ram_ix167_a_230__dup_2423), .C (
                     modgen_ram_ix167_a_229__dup_2424), .D (
                     modgen_ram_ix167_a_231__dup_2422), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix5177 (.Y (nx5176), .A0 (rd_addr_m_1), .A1 (nx917), .B0 (
                          nx3299), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix918 (.Y (nx917), .A (modgen_ram_ix167_a_224__dup_2429), 
                      .B (modgen_ram_ix167_a_225__dup_2428), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2507 (.Y (nx3299), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_2426), .B0 (nx5150), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix5151 (.Y (nx5150), .AN (modgen_ram_ix167_a_226__dup_2427
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2508 (.Y (nx3300), .A0 (rd_addr_m_2), .A1 (nx5428), 
                          .B0 (nx5348), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix5429 (.Y (nx5428), .A (modgen_ram_ix167_a_236__dup_2417)
                     , .B (modgen_ram_ix167_a_238__dup_2415), .C (
                     modgen_ram_ix167_a_237__dup_2416), .D (
                     modgen_ram_ix167_a_239__dup_2414), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix5349 (.Y (nx5348), .A0 (rd_addr_m_1), .A1 (nx928), .B0 (
                          nx3301), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix929 (.Y (nx928), .A (modgen_ram_ix167_a_232__dup_2421), 
                      .B (modgen_ram_ix167_a_233__dup_2420), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2510 (.Y (nx3301), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_2418), .B0 (nx5322), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix5323 (.Y (nx5322), .AN (modgen_ram_ix167_a_234__dup_2419
                      ), .B (rd_addr_m_0)) ;
    INV_X0P5B_A12TS ix934 (.Y (nx933), .A (rd_addr_m_6)) ;
    OA21A1OI2_X0P5M_A12TS ix2511 (.Y (nx4380), .A0 (rd_addr_m_5), .A1 (nx3303), 
                          .B0 (nx967), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2512 (.Y (nx3303), .A0 (rd_addr_m_4), .A1 (nx3664), .B0 (
                      nx3318)) ;
    MXT4_X0P5M_A12TS ix3665 (.Y (nx3664), .A (nx3400), .B (nx3572), .C (nx3260)
                     , .D (nx3261), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix3401 (.Y (nx3400), .A (modgen_ram_ix167_a_144__dup_2509)
                     , .B (modgen_ram_ix167_a_146__dup_2507), .C (
                     modgen_ram_ix167_a_145__dup_2508), .D (
                     modgen_ram_ix167_a_147__dup_2506), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix3573 (.Y (nx3572), .A (modgen_ram_ix167_a_152__dup_2501)
                     , .B (modgen_ram_ix167_a_154__dup_2499), .C (
                     modgen_ram_ix167_a_153__dup_2500), .D (
                     modgen_ram_ix167_a_155__dup_2498), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2514 (.Y (nx3260), .A (modgen_ram_ix167_a_148__dup_2505)
                     , .B (modgen_ram_ix167_a_150__dup_2503), .C (
                     modgen_ram_ix167_a_149__dup_2504), .D (
                     modgen_ram_ix167_a_151__dup_2502), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2515 (.Y (nx3261), .A (modgen_ram_ix167_a_156__dup_2497)
                     , .B (modgen_ram_ix167_a_158__dup_2495), .C (
                     modgen_ram_ix167_a_157__dup_2496), .D (
                     modgen_ram_ix167_a_159__dup_2494), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix3319 (.Y (nx3318), .A0 (rd_addr_m_3), .A1 (nx947), .B0 (
                          nx3305), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix948 (.Y (nx947), .A0 (rd_addr_m_2), .A1 (nx3134), .B0 (
                      nx3054)) ;
    MXT4_X0P5M_A12TS ix3135 (.Y (nx3134), .A (modgen_ram_ix167_a_132__dup_2521)
                     , .B (modgen_ram_ix167_a_134__dup_2519), .C (
                     modgen_ram_ix167_a_133__dup_2520), .D (
                     modgen_ram_ix167_a_135__dup_2518), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix3055 (.Y (nx3054), .A0 (rd_addr_m_1), .A1 (nx951), .B0 (
                          nx3304), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix952 (.Y (nx951), .A (modgen_ram_ix167_a_128__dup_2525), 
                      .B (modgen_ram_ix167_a_129__dup_2524), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2517 (.Y (nx3304), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_2522), .B0 (nx3028), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix3029 (.Y (nx3028), .AN (modgen_ram_ix167_a_130__dup_2523
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2518 (.Y (nx3305), .A0 (rd_addr_m_2), .A1 (nx3306), 
                          .B0 (nx3259), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix3307 (.Y (nx3306), .A (modgen_ram_ix167_a_140__dup_2513)
                     , .B (modgen_ram_ix167_a_142__dup_2511), .C (
                     modgen_ram_ix167_a_141__dup_2512), .D (
                     modgen_ram_ix167_a_143__dup_2510), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix3227 (.Y (nx3259), .A0 (rd_addr_m_1), .A1 (nx961), .B0 (
                          nx3307), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix962 (.Y (nx961), .A (modgen_ram_ix167_a_136__dup_2517), 
                      .B (modgen_ram_ix167_a_137__dup_2516), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2519 (.Y (nx3307), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_2514), .B0 (nx3200), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix3201 (.Y (nx3200), .AN (modgen_ram_ix167_a_138__dup_2515
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix968 (.Y (nx967), .A0 (rd_addr_m_4), .A1 (nx4368), .B0 (
                          nx4022), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix2520 (.Y (nx4368), .A (nx4104), .B (nx4276), .C (nx3262)
                     , .D (nx4360), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix4105 (.Y (nx4104), .A (modgen_ram_ix167_a_176__dup_2477)
                     , .B (modgen_ram_ix167_a_178__dup_2475), .C (
                     modgen_ram_ix167_a_177__dup_2476), .D (
                     modgen_ram_ix167_a_179__dup_2474), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix4277 (.Y (nx4276), .A (modgen_ram_ix167_a_184__dup_2469)
                     , .B (modgen_ram_ix167_a_186__dup_2467), .C (
                     modgen_ram_ix167_a_185__dup_2468), .D (
                     modgen_ram_ix167_a_187__dup_2466), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2521 (.Y (nx3262), .A (modgen_ram_ix167_a_180__dup_2473)
                     , .B (modgen_ram_ix167_a_182__dup_2471), .C (
                     modgen_ram_ix167_a_181__dup_2472), .D (
                     modgen_ram_ix167_a_183__dup_2470), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix4361 (.Y (nx4360), .A (modgen_ram_ix167_a_188__dup_2465)
                     , .B (modgen_ram_ix167_a_190__dup_2463), .C (
                     modgen_ram_ix167_a_189__dup_2464), .D (
                     modgen_ram_ix167_a_191__dup_2462), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix4023 (.Y (nx4022), .A0 (rd_addr_m_3), .A1 (nx3309), 
                          .B0 (nx3312), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2523 (.Y (nx3309), .A0 (rd_addr_m_2), .A1 (nx3838), .B0 (
                      nx3758)) ;
    MXT4_X0P5M_A12TS ix3839 (.Y (nx3838), .A (modgen_ram_ix167_a_164__dup_2489)
                     , .B (modgen_ram_ix167_a_166__dup_2487), .C (
                     modgen_ram_ix167_a_165__dup_2488), .D (
                     modgen_ram_ix167_a_167__dup_2486), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix3759 (.Y (nx3758), .A0 (rd_addr_m_1), .A1 (nx3310), 
                          .B0 (nx3311), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix980 (.Y (nx3310), .A (modgen_ram_ix167_a_160__dup_2493)
                      , .B (modgen_ram_ix167_a_161__dup_2492), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix982 (.Y (nx3311), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_2490), .B0 (nx3732), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix3733 (.Y (nx3732), .AN (modgen_ram_ix167_a_162__dup_2491
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix986 (.Y (nx3312), .A0 (rd_addr_m_2), .A1 (nx4010), .B0 (
                          nx3930), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix4011 (.Y (nx4010), .A (modgen_ram_ix167_a_172__dup_2481)
                     , .B (modgen_ram_ix167_a_174__dup_2479), .C (
                     modgen_ram_ix167_a_173__dup_2480), .D (
                     modgen_ram_ix167_a_175__dup_2478), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix3931 (.Y (nx3930), .A0 (rd_addr_m_1), .A1 (nx3313), 
                          .B0 (nx3314), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2524 (.Y (nx3313), .A (modgen_ram_ix167_a_168__dup_2485)
                      , .B (modgen_ram_ix167_a_169__dup_2484), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix992 (.Y (nx3314), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_2482), .B0 (nx3904), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix3905 (.Y (nx3904), .AN (modgen_ram_ix167_a_170__dup_2483
                      ), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix2965 (.Y (nx2964), .A (rd_addr_7), .B (nx3315)) ;
    AOI21_X0P5M_A12TS ix998 (.Y (nx3315), .A0 (rd_addr_m_6), .A1 (nx2956), .B0 (
                      nx1544)) ;
    OAI21_X0P5M_A12TS ix2957 (.Y (nx2956), .A0 (rd_addr_m_5), .A1 (nx3316), .B0 (
                      nx1033)) ;
    AOI21_X0P5M_A12TS ix1002 (.Y (nx3316), .A0 (rd_addr_m_4), .A1 (nx2244), .B0 (
                      nx3245)) ;
    MXT4_X0P5M_A12TS ix2525 (.Y (nx2244), .A (nx1980), .B (nx3248), .C (nx2064)
                     , .D (nx3249), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix2526 (.Y (nx1980), .A (modgen_ram_ix167_a_80__dup_2573), 
                     .B (modgen_ram_ix167_a_82__dup_2571), .C (
                     modgen_ram_ix167_a_81__dup_2572), .D (
                     modgen_ram_ix167_a_83__dup_2570), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2153 (.Y (nx3248), .A (modgen_ram_ix167_a_88__dup_2565), 
                     .B (modgen_ram_ix167_a_90__dup_2563), .C (
                     modgen_ram_ix167_a_89__dup_2564), .D (
                     modgen_ram_ix167_a_91__dup_2562), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2065 (.Y (nx2064), .A (modgen_ram_ix167_a_84__dup_2569), 
                     .B (modgen_ram_ix167_a_86__dup_2567), .C (
                     modgen_ram_ix167_a_85__dup_2568), .D (
                     modgen_ram_ix167_a_87__dup_2566), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2528 (.Y (nx3249), .A (modgen_ram_ix167_a_92__dup_2561), 
                     .B (modgen_ram_ix167_a_94__dup_2559), .C (
                     modgen_ram_ix167_a_93__dup_2560), .D (
                     modgen_ram_ix167_a_95__dup_2558), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2529 (.Y (nx3245), .A0 (rd_addr_m_3), .A1 (nx1011), 
                          .B0 (nx1021), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2530 (.Y (nx1011), .A0 (rd_addr_m_2), .A1 (nx3241), .B0 (
                      nx1634)) ;
    MXT4_X0P5M_A12TS ix2531 (.Y (nx3241), .A (modgen_ram_ix167_a_68__dup_2585), 
                     .B (modgen_ram_ix167_a_70__dup_2583), .C (
                     modgen_ram_ix167_a_69__dup_2584), .D (
                     modgen_ram_ix167_a_71__dup_2582), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2532 (.Y (nx1634), .A0 (rd_addr_m_1), .A1 (nx3317), 
                          .B0 (nx1018), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2534 (.Y (nx3317), .A (modgen_ram_ix167_a_64__dup_2589)
                      , .B (modgen_ram_ix167_a_65__dup_2588), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2535 (.Y (nx1018), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_2586), .B0 (nx1608), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2536 (.Y (nx1608), .AN (modgen_ram_ix167_a_66__dup_2587)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2538 (.Y (nx1021), .A0 (rd_addr_m_2), .A1 (nx3244), 
                          .B0 (nx3243), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix1887 (.Y (nx3244), .A (modgen_ram_ix167_a_76__dup_2577), 
                     .B (modgen_ram_ix167_a_78__dup_2575), .C (
                     modgen_ram_ix167_a_77__dup_2576), .D (
                     modgen_ram_ix167_a_79__dup_2574), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix1807 (.Y (nx3243), .A0 (rd_addr_m_1), .A1 (nx1027), 
                          .B0 (nx1029), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2539 (.Y (nx1027), .A (modgen_ram_ix167_a_72__dup_2581)
                      , .B (modgen_ram_ix167_a_73__dup_2580), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2540 (.Y (nx1029), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_2578), .B0 (nx3242), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2541 (.Y (nx3242), .AN (modgen_ram_ix167_a_74__dup_2579)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2542 (.Y (nx1033), .A0 (rd_addr_m_4), .A1 (nx2948), 
                          .B0 (nx3256), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix2949 (.Y (nx2948), .A (nx3258), .B (nx2856), .C (nx2768)
                     , .D (nx2940), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix2544 (.Y (nx3258), .A (modgen_ram_ix167_a_112__dup_2541)
                     , .B (modgen_ram_ix167_a_114__dup_2539), .C (
                     modgen_ram_ix167_a_113__dup_2540), .D (
                     modgen_ram_ix167_a_115__dup_2538), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2857 (.Y (nx2856), .A (modgen_ram_ix167_a_120__dup_2533)
                     , .B (modgen_ram_ix167_a_122__dup_2531), .C (
                     modgen_ram_ix167_a_121__dup_2532), .D (
                     modgen_ram_ix167_a_123__dup_2530), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2769 (.Y (nx2768), .A (modgen_ram_ix167_a_116__dup_2537)
                     , .B (modgen_ram_ix167_a_118__dup_2535), .C (
                     modgen_ram_ix167_a_117__dup_2536), .D (
                     modgen_ram_ix167_a_119__dup_2534), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2941 (.Y (nx2940), .A (modgen_ram_ix167_a_124__dup_2529)
                     , .B (modgen_ram_ix167_a_126__dup_2527), .C (
                     modgen_ram_ix167_a_125__dup_2528), .D (
                     modgen_ram_ix167_a_127__dup_2526), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2546 (.Y (nx3256), .A0 (rd_addr_m_3), .A1 (nx1043), 
                          .B0 (nx3319), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1044 (.Y (nx1043), .A0 (rd_addr_m_2), .A1 (nx3253), .B0 (
                      nx3252)) ;
    MXT4_X0P5M_A12TS ix2548 (.Y (nx3253), .A (modgen_ram_ix167_a_100__dup_2553)
                     , .B (modgen_ram_ix167_a_102__dup_2551), .C (
                     modgen_ram_ix167_a_101__dup_2552), .D (
                     modgen_ram_ix167_a_103__dup_2550), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2550 (.Y (nx3252), .A0 (rd_addr_m_1), .A1 (nx1049), 
                          .B0 (nx1051), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1050 (.Y (nx1049), .A (modgen_ram_ix167_a_96__dup_2557)
                      , .B (modgen_ram_ix167_a_97__dup_2556), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1052 (.Y (nx1051), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_2554), .B0 (nx3251), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2552 (.Y (nx3251), .AN (modgen_ram_ix167_a_98__dup_2555)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1056 (.Y (nx3319), .A0 (rd_addr_m_2), .A1 (nx2590), 
                          .B0 (nx2510), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix2554 (.Y (nx2590), .A (modgen_ram_ix167_a_108__dup_2545)
                     , .B (modgen_ram_ix167_a_110__dup_2543), .C (
                     modgen_ram_ix167_a_109__dup_2544), .D (
                     modgen_ram_ix167_a_111__dup_2542), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2556 (.Y (nx2510), .A0 (rd_addr_m_1), .A1 (nx3321), 
                          .B0 (nx3322), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1060 (.Y (nx3321), .A (modgen_ram_ix167_a_104__dup_2549)
                      , .B (modgen_ram_ix167_a_105__dup_2548), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1062 (.Y (nx3322), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_2546), .B0 (nx3255), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2557 (.Y (nx3255), .AN (modgen_ram_ix167_a_106__dup_2547
                      ), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2561 (.Y (nx1544), .A0 (rd_addr_m_5), .A1 (nx1067), 
                          .B0 (nx1099), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2564 (.Y (nx1067), .A0 (rd_addr_m_4), .A1 (nx818), .B0 (
                      nx3226)) ;
    MXT4_X0P5M_A12TS ix819 (.Y (nx818), .A (nx3229), .B (nx726), .C (nx638), .D (
                     nx3230), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix2566 (.Y (nx3229), .A (modgen_ram_ix167_a_16__dup_2637), 
                     .B (modgen_ram_ix167_a_18__dup_2635), .C (
                     modgen_ram_ix167_a_17__dup_2636), .D (
                     modgen_ram_ix167_a_19__dup_2634), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix727 (.Y (nx726), .A (modgen_ram_ix167_a_24__dup_2629), .B (
                     modgen_ram_ix167_a_26__dup_2627), .C (
                     modgen_ram_ix167_a_25__dup_2628), .D (
                     modgen_ram_ix167_a_27__dup_2626), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix639 (.Y (nx638), .A (modgen_ram_ix167_a_20__dup_2633), .B (
                     modgen_ram_ix167_a_22__dup_2631), .C (
                     modgen_ram_ix167_a_21__dup_2632), .D (
                     modgen_ram_ix167_a_23__dup_2630), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2568 (.Y (nx3230), .A (modgen_ram_ix167_a_28__dup_2625), 
                     .B (modgen_ram_ix167_a_30__dup_2623), .C (
                     modgen_ram_ix167_a_29__dup_2624), .D (
                     modgen_ram_ix167_a_31__dup_2622), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2570 (.Y (nx3226), .A0 (rd_addr_m_3), .A1 (nx3323), 
                          .B0 (nx1087), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2571 (.Y (nx3323), .A0 (rd_addr_m_2), .A1 (nx3219), .B0 (
                      nx166)) ;
    MXT4_X0P5M_A12TS ix2572 (.Y (nx3219), .A (modgen_ram_ix167_a_4__dup_2649), .B (
                     modgen_ram_ix167_a_6__dup_2647), .C (
                     modgen_ram_ix167_a_5__dup_2648), .D (
                     modgen_ram_ix167_a_7__dup_2646), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix167 (.Y (nx166), .A0 (rd_addr_m_1), .A1 (nx1081), .B0 (
                          nx1083), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2574 (.Y (nx1081), .A (modgen_ram_ix167_a_0__dup_2653), 
                      .B (modgen_ram_ix167_a_1__dup_2652), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2576 (.Y (nx1083), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_2650), .B0 (nx132), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix133 (.Y (nx132), .AN (modgen_ram_ix167_a_2__dup_2651), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2578 (.Y (nx1087), .A0 (rd_addr_m_2), .A1 (nx456), .B0 (
                          nx362), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix457 (.Y (nx456), .A (modgen_ram_ix167_a_12__dup_2641), .B (
                     modgen_ram_ix167_a_14__dup_2639), .C (
                     modgen_ram_ix167_a_13__dup_2640), .D (
                     modgen_ram_ix167_a_15__dup_2638), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix363 (.Y (nx362), .A0 (rd_addr_m_1), .A1 (nx1093), .B0 (
                          nx1095), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2580 (.Y (nx1093), .A (modgen_ram_ix167_a_8__dup_2645), 
                      .B (modgen_ram_ix167_a_9__dup_2644), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1096 (.Y (nx1095), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_2642), .B0 (nx3221), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2582 (.Y (nx3221), .AN (modgen_ram_ix167_a_10__dup_2643)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1100 (.Y (nx1099), .A0 (rd_addr_m_4), .A1 (nx1532), 
                          .B0 (nx3238), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix2584 (.Y (nx1532), .A (nx1268), .B (nx1440), .C (nx3240)
                     , .D (nx1524), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix2586 (.Y (nx1268), .A (modgen_ram_ix167_a_48__dup_2605), 
                     .B (modgen_ram_ix167_a_50__dup_2603), .C (
                     modgen_ram_ix167_a_49__dup_2604), .D (
                     modgen_ram_ix167_a_51__dup_2602), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2587 (.Y (nx1440), .A (modgen_ram_ix167_a_56__dup_2597), 
                     .B (modgen_ram_ix167_a_58__dup_2595), .C (
                     modgen_ram_ix167_a_57__dup_2596), .D (
                     modgen_ram_ix167_a_59__dup_2594), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2593 (.Y (nx3240), .A (modgen_ram_ix167_a_52__dup_2601), 
                     .B (modgen_ram_ix167_a_54__dup_2599), .C (
                     modgen_ram_ix167_a_53__dup_2600), .D (
                     modgen_ram_ix167_a_55__dup_2598), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2594 (.Y (nx1524), .A (modgen_ram_ix167_a_60__dup_2593), 
                     .B (modgen_ram_ix167_a_62__dup_2591), .C (
                     modgen_ram_ix167_a_61__dup_2592), .D (
                     modgen_ram_ix167_a_63__dup_2590), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2596 (.Y (nx3238), .A0 (rd_addr_m_3), .A1 (nx1107), 
                          .B0 (nx1117), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1108 (.Y (nx1107), .A0 (rd_addr_m_2), .A1 (nx3235), .B0 (
                      nx3233)) ;
    MXT4_X0P5M_A12TS ix2598 (.Y (nx3235), .A (modgen_ram_ix167_a_36__dup_2617), 
                     .B (modgen_ram_ix167_a_38__dup_2615), .C (
                     modgen_ram_ix167_a_37__dup_2616), .D (
                     modgen_ram_ix167_a_39__dup_2614), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2600 (.Y (nx3233), .A0 (rd_addr_m_1), .A1 (nx1111), 
                          .B0 (nx1113), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1112 (.Y (nx1111), .A (modgen_ram_ix167_a_32__dup_2621)
                      , .B (modgen_ram_ix167_a_33__dup_2620), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1114 (.Y (nx1113), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_2618), .B0 (nx3232), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2601 (.Y (nx3232), .AN (modgen_ram_ix167_a_34__dup_2619)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1118 (.Y (nx1117), .A0 (rd_addr_m_2), .A1 (nx3237), 
                          .B0 (nx1088), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix2602 (.Y (nx3237), .A (modgen_ram_ix167_a_44__dup_2609), 
                     .B (modgen_ram_ix167_a_46__dup_2607), .C (
                     modgen_ram_ix167_a_45__dup_2608), .D (
                     modgen_ram_ix167_a_47__dup_2606), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2604 (.Y (nx1088), .A0 (rd_addr_m_1), .A1 (nx1121), 
                          .B0 (nx1123), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1122 (.Y (nx1121), .A (modgen_ram_ix167_a_40__dup_2613)
                      , .B (modgen_ram_ix167_a_41__dup_2612), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1124 (.Y (nx1123), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_2610), .B0 (nx3236), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix1063 (.Y (nx3236), .AN (modgen_ram_ix167_a_42__dup_2611)
                      , .B (rd_addr_m_0)) ;
    NAND4_X0P5A_A12TS ix1128 (.Y (nx1127), .A (nx3208), .B (nx3212), .C (nx1142)
                      , .D (nx3325)) ;
    NOR3_X0P5A_A12TS ix2606 (.Y (nx3208), .A (nx1131), .B (nx3205), .C (nx3207)
                     ) ;
    NAND3_X0P5A_A12TS ix1132 (.Y (nx1131), .A (nx1133), .B (NOT_rd_en), .C (
                      wr_dup_1054)) ;
    XNOR2_X0P5M_A12TS ix1134 (.Y (nx1133), .A (wr_addr_m_0), .B (rd_addr_m_0)) ;
    XOR2_X0P5M_A12TS ix2608 (.Y (nx3205), .A (wr_addr_m_1), .B (rd_addr_m_1)) ;
    XOR2_X0P5M_A12TS ix2610 (.Y (nx3207), .A (wr_addr_m_2), .B (rd_addr_m_2)) ;
    NOR3_X0P5A_A12TS ix2612 (.Y (nx3212), .A (nx3209), .B (nx3210), .C (nx3211)
                     ) ;
    XOR2_X0P5M_A12TS ix2614 (.Y (nx3209), .A (wr_addr_m_5), .B (rd_addr_m_5)) ;
    XOR2_X0P5M_A12TS ix2616 (.Y (nx3210), .A (wr_addr_m_3), .B (rd_addr_m_3)) ;
    XOR2_X0P5M_A12TS ix2617 (.Y (nx3211), .A (wr_addr_m_4), .B (rd_addr_m_4)) ;
    XNOR2_X0P5M_A12TS ix1143 (.Y (nx1142), .A (wr_addr_m_6), .B (rd_addr_m_6)) ;
    XNOR2_X0P5M_A12TS ix1145 (.Y (nx3325), .A (wr_addr_7), .B (rd_addr_7)) ;
    INV_X0P5B_A12TS ix2619 (.Y (NOT_nx50), .A (NOT_rd_en)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_1 (.Q (rd_data_m_1), .CK (wb_clk_i), .D (
                        nx9398), .R (wb_rst_i), .SE (NOT_nx50), .SI (rd_data_m_1
                        )) ;
    MXIT2_X0P5M_A12TS ix9399 (.Y (nx9398), .A (nx3326), .B (nx3327), .S0 (nx1127
                      )) ;
    INV_X0P5B_A12TS ix1154 (.Y (nx3326), .A (wr_data_m_1)) ;
    OA21A1OI2_X0P5M_A12TS ix1156 (.Y (nx3327), .A0 (nx9384), .A1 (nx3281), .B0 (
                          rd_addr_7), .C0 (nx7602)) ;
    OA21A1OI2_X0P5M_A12TS ix9385 (.Y (nx9384), .A0 (rd_addr_m_5), .A1 (nx1158), 
                          .B0 (nx1191), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2621 (.Y (nx1158), .A0 (rd_addr_m_4), .A1 (nx3284), .B0 (
                      nx8714)) ;
    MXT4_X0P5M_A12TS ix2623 (.Y (nx3284), .A (nx8762), .B (nx8870), .C (nx8814)
                     , .D (nx8922), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix8763 (.Y (nx8762), .A (modgen_ram_ix167_a_208__dup_2181)
                     , .B (modgen_ram_ix167_a_210__dup_2179), .C (
                     modgen_ram_ix167_a_209__dup_2180), .D (
                     modgen_ram_ix167_a_211__dup_2178), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix8871 (.Y (nx8870), .A (modgen_ram_ix167_a_216__dup_2173)
                     , .B (modgen_ram_ix167_a_218__dup_2171), .C (
                     modgen_ram_ix167_a_217__dup_2172), .D (
                     modgen_ram_ix167_a_219__dup_2170), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix8815 (.Y (nx8814), .A (modgen_ram_ix167_a_212__dup_2177)
                     , .B (modgen_ram_ix167_a_214__dup_2175), .C (
                     modgen_ram_ix167_a_213__dup_2176), .D (
                     modgen_ram_ix167_a_215__dup_2174), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix8923 (.Y (nx8922), .A (modgen_ram_ix167_a_220__dup_2169)
                     , .B (modgen_ram_ix167_a_222__dup_2167), .C (
                     modgen_ram_ix167_a_221__dup_2168), .D (
                     modgen_ram_ix167_a_223__dup_2166), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix8715 (.Y (nx8714), .A0 (rd_addr_m_3), .A1 (nx1169), 
                          .B0 (nx1181), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1170 (.Y (nx1169), .A0 (rd_addr_m_2), .A1 (nx8594), .B0 (
                      nx3283)) ;
    MXT4_X0P5M_A12TS ix8595 (.Y (nx8594), .A (modgen_ram_ix167_a_196__dup_2193)
                     , .B (modgen_ram_ix167_a_198__dup_2191), .C (
                     modgen_ram_ix167_a_197__dup_2192), .D (
                     modgen_ram_ix167_a_199__dup_2190), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2624 (.Y (nx3283), .A0 (rd_addr_m_1), .A1 (nx3328), 
                          .B0 (nx3329), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1176 (.Y (nx3328), .A (modgen_ram_ix167_a_192__dup_2197)
                      , .B (modgen_ram_ix167_a_193__dup_2196), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1178 (.Y (nx3329), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_2194), .B0 (nx3282), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2626 (.Y (nx3282), .AN (modgen_ram_ix167_a_194__dup_2195
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1182 (.Y (nx1181), .A0 (rd_addr_m_2), .A1 (nx8702), 
                          .B0 (nx8654), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix8703 (.Y (nx8702), .A (modgen_ram_ix167_a_204__dup_2185)
                     , .B (modgen_ram_ix167_a_206__dup_2183), .C (
                     modgen_ram_ix167_a_205__dup_2184), .D (
                     modgen_ram_ix167_a_207__dup_2182), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix8655 (.Y (nx8654), .A0 (rd_addr_m_1), .A1 (nx1185), 
                          .B0 (nx1187), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2628 (.Y (nx1185), .A (modgen_ram_ix167_a_200__dup_2189)
                      , .B (modgen_ram_ix167_a_201__dup_2188), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2630 (.Y (nx1187), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_2186), .B0 (nx8636), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix8637 (.Y (nx8636), .AN (modgen_ram_ix167_a_202__dup_2187
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2631 (.Y (nx1191), .A0 (rd_addr_m_4), .A1 (nx9374), 
                          .B0 (nx9158), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix9375 (.Y (nx9374), .A (nx9206), .B (nx9314), .C (nx9258)
                     , .D (nx9366), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix9207 (.Y (nx9206), .A (modgen_ram_ix167_a_240__dup_2149)
                     , .B (modgen_ram_ix167_a_242__dup_2147), .C (
                     modgen_ram_ix167_a_241__dup_2148), .D (
                     modgen_ram_ix167_a_243__dup_2146), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix9315 (.Y (nx9314), .A (modgen_ram_ix167_a_248__dup_2141)
                     , .B (modgen_ram_ix167_a_250__dup_2139), .C (
                     modgen_ram_ix167_a_249__dup_2140), .D (
                     modgen_ram_ix167_a_251__dup_2138), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix9259 (.Y (nx9258), .A (modgen_ram_ix167_a_244__dup_2145)
                     , .B (modgen_ram_ix167_a_246__dup_2143), .C (
                     modgen_ram_ix167_a_245__dup_2144), .D (
                     modgen_ram_ix167_a_247__dup_2142), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix9367 (.Y (nx9366), .A (modgen_ram_ix167_a_252__dup_2137)
                     , .B (modgen_ram_ix167_a_254__dup_2135), .C (
                     modgen_ram_ix167_a_253__dup_2136), .D (
                     modgen_ram_ix167_a_255__dup_2134), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix9159 (.Y (nx9158), .A0 (rd_addr_m_3), .A1 (nx1202), 
                          .B0 (nx1213), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2632 (.Y (nx1202), .A0 (rd_addr_m_2), .A1 (nx3285), .B0 (
                      nx8990)) ;
    MXT4_X0P5M_A12TS ix2634 (.Y (nx3285), .A (modgen_ram_ix167_a_228__dup_2161)
                     , .B (modgen_ram_ix167_a_230__dup_2159), .C (
                     modgen_ram_ix167_a_229__dup_2160), .D (
                     modgen_ram_ix167_a_231__dup_2158), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix8991 (.Y (nx8990), .A0 (rd_addr_m_1), .A1 (nx1207), 
                          .B0 (nx1209), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2636 (.Y (nx1207), .A (modgen_ram_ix167_a_224__dup_2165)
                      , .B (modgen_ram_ix167_a_225__dup_2164), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2638 (.Y (nx1209), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_2162), .B0 (nx8972), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix8973 (.Y (nx8972), .AN (modgen_ram_ix167_a_226__dup_2163
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2640 (.Y (nx1213), .A0 (rd_addr_m_2), .A1 (nx9146), 
                          .B0 (nx9098), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix9147 (.Y (nx9146), .A (modgen_ram_ix167_a_236__dup_2153)
                     , .B (modgen_ram_ix167_a_238__dup_2151), .C (
                     modgen_ram_ix167_a_237__dup_2152), .D (
                     modgen_ram_ix167_a_239__dup_2150), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix9099 (.Y (nx9098), .A0 (rd_addr_m_1), .A1 (nx1218), 
                          .B0 (nx1220), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2642 (.Y (nx1218), .A (modgen_ram_ix167_a_232__dup_2157)
                      , .B (modgen_ram_ix167_a_233__dup_2156), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2644 (.Y (nx1220), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_2154), .B0 (nx9080), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix9081 (.Y (nx9080), .AN (modgen_ram_ix167_a_234__dup_2155
                      ), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2646 (.Y (nx3281), .A0 (rd_addr_m_5), .A1 (nx1225), 
                          .B0 (nx3336), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix1226 (.Y (nx1225), .A0 (rd_addr_m_4), .A1 (nx8038), .B0 (
                      nx7822)) ;
    MXT4_X0P5M_A12TS ix8039 (.Y (nx8038), .A (nx7870), .B (nx7978), .C (nx7922)
                     , .D (nx8030), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix7871 (.Y (nx7870), .A (modgen_ram_ix167_a_144__dup_2245)
                     , .B (modgen_ram_ix167_a_146__dup_2243), .C (
                     modgen_ram_ix167_a_145__dup_2244), .D (
                     modgen_ram_ix167_a_147__dup_2242), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2647 (.Y (nx7978), .A (modgen_ram_ix167_a_152__dup_2237)
                     , .B (modgen_ram_ix167_a_154__dup_2235), .C (
                     modgen_ram_ix167_a_153__dup_2236), .D (
                     modgen_ram_ix167_a_155__dup_2234), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix7923 (.Y (nx7922), .A (modgen_ram_ix167_a_148__dup_2241)
                     , .B (modgen_ram_ix167_a_150__dup_2239), .C (
                     modgen_ram_ix167_a_149__dup_2240), .D (
                     modgen_ram_ix167_a_151__dup_2238), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix8031 (.Y (nx8030), .A (modgen_ram_ix167_a_156__dup_2233)
                     , .B (modgen_ram_ix167_a_158__dup_2231), .C (
                     modgen_ram_ix167_a_157__dup_2232), .D (
                     modgen_ram_ix167_a_159__dup_2230), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix7823 (.Y (nx7822), .A0 (rd_addr_m_3), .A1 (nx3330), 
                          .B0 (nx3333), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1236 (.Y (nx3330), .A0 (rd_addr_m_2), .A1 (nx7702), .B0 (
                      nx3276)) ;
    MXT4_X0P5M_A12TS ix7703 (.Y (nx7702), .A (modgen_ram_ix167_a_132__dup_2257)
                     , .B (modgen_ram_ix167_a_134__dup_2255), .C (
                     modgen_ram_ix167_a_133__dup_2256), .D (
                     modgen_ram_ix167_a_135__dup_2254), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2651 (.Y (nx3276), .A0 (rd_addr_m_1), .A1 (nx3331), 
                          .B0 (nx3332), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2653 (.Y (nx3331), .A (modgen_ram_ix167_a_128__dup_2261)
                      , .B (modgen_ram_ix167_a_129__dup_2260), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2654 (.Y (nx3332), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_2258), .B0 (nx7636), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix7637 (.Y (nx7636), .AN (modgen_ram_ix167_a_130__dup_2259
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1246 (.Y (nx3333), .A0 (rd_addr_m_2), .A1 (nx7810), 
                          .B0 (nx7762), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix7811 (.Y (nx7810), .A (modgen_ram_ix167_a_140__dup_2249)
                     , .B (modgen_ram_ix167_a_142__dup_2247), .C (
                     modgen_ram_ix167_a_141__dup_2248), .D (
                     modgen_ram_ix167_a_143__dup_2246), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix7763 (.Y (nx7762), .A0 (rd_addr_m_1), .A1 (nx3334), 
                          .B0 (nx3335), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1252 (.Y (nx3334), .A (modgen_ram_ix167_a_136__dup_2253)
                      , .B (modgen_ram_ix167_a_137__dup_2252), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1254 (.Y (nx3335), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_2250), .B0 (nx3277), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix2656 (.Y (nx3277), .AN (modgen_ram_ix167_a_138__dup_2251
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1258 (.Y (nx3336), .A0 (rd_addr_m_4), .A1 (nx8482), 
                          .B0 (nx8266), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix8483 (.Y (nx8482), .A (nx8314), .B (nx3279), .C (nx8366)
                     , .D (nx3280), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix8315 (.Y (nx8314), .A (modgen_ram_ix167_a_176__dup_2213)
                     , .B (modgen_ram_ix167_a_178__dup_2211), .C (
                     modgen_ram_ix167_a_177__dup_2212), .D (
                     modgen_ram_ix167_a_179__dup_2210), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2658 (.Y (nx3279), .A (modgen_ram_ix167_a_184__dup_2205)
                     , .B (modgen_ram_ix167_a_186__dup_2203), .C (
                     modgen_ram_ix167_a_185__dup_2204), .D (
                     modgen_ram_ix167_a_187__dup_2202), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix8367 (.Y (nx8366), .A (modgen_ram_ix167_a_180__dup_2209)
                     , .B (modgen_ram_ix167_a_182__dup_2207), .C (
                     modgen_ram_ix167_a_181__dup_2208), .D (
                     modgen_ram_ix167_a_183__dup_2206), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2660 (.Y (nx3280), .A (modgen_ram_ix167_a_188__dup_2201)
                     , .B (modgen_ram_ix167_a_190__dup_2199), .C (
                     modgen_ram_ix167_a_189__dup_2200), .D (
                     modgen_ram_ix167_a_191__dup_2198), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix8267 (.Y (nx8266), .A0 (rd_addr_m_3), .A1 (nx1267), 
                          .B0 (nx1279), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2661 (.Y (nx1267), .A0 (rd_addr_m_2), .A1 (nx8146), .B0 (
                      nx3278)) ;
    MXT4_X0P5M_A12TS ix8147 (.Y (nx8146), .A (modgen_ram_ix167_a_164__dup_2225)
                     , .B (modgen_ram_ix167_a_166__dup_2223), .C (
                     modgen_ram_ix167_a_165__dup_2224), .D (
                     modgen_ram_ix167_a_167__dup_2222), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2662 (.Y (nx3278), .A0 (rd_addr_m_1), .A1 (nx1273), 
                          .B0 (nx1275), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2664 (.Y (nx1273), .A (modgen_ram_ix167_a_160__dup_2229)
                      , .B (modgen_ram_ix167_a_161__dup_2228), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2666 (.Y (nx1275), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_2226), .B0 (nx8080), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix8081 (.Y (nx8080), .AN (modgen_ram_ix167_a_162__dup_2227
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2668 (.Y (nx1279), .A0 (rd_addr_m_2), .A1 (nx8254), 
                          .B0 (nx8206), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix8255 (.Y (nx8254), .A (modgen_ram_ix167_a_172__dup_2217)
                     , .B (modgen_ram_ix167_a_174__dup_2215), .C (
                     modgen_ram_ix167_a_173__dup_2216), .D (
                     modgen_ram_ix167_a_175__dup_2214), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix8207 (.Y (nx8206), .A0 (rd_addr_m_1), .A1 (nx1284), 
                          .B0 (nx1286), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2670 (.Y (nx1284), .A (modgen_ram_ix167_a_168__dup_2221)
                      , .B (modgen_ram_ix167_a_169__dup_2220), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2672 (.Y (nx1286), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_2218), .B0 (nx8188), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix8189 (.Y (nx8188), .AN (modgen_ram_ix167_a_170__dup_2219
                      ), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix7603 (.Y (nx7602), .A (rd_addr_7), .B (nx1291)) ;
    AOI21_X0P5M_A12TS ix2674 (.Y (nx1291), .A0 (rd_addr_m_6), .A1 (nx7594), .B0 (
                      nx6706)) ;
    OAI21_X0P5M_A12TS ix7595 (.Y (nx7594), .A0 (rd_addr_m_5), .A1 (nx1295), .B0 (
                      nx1326)) ;
    AOI21_X0P5M_A12TS ix2676 (.Y (nx1295), .A0 (rd_addr_m_4), .A1 (nx7142), .B0 (
                      nx6926)) ;
    MXT4_X0P5M_A12TS ix7143 (.Y (nx7142), .A (nx6974), .B (nx7082), .C (nx7026)
                     , .D (nx3272), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix6975 (.Y (nx6974), .A (modgen_ram_ix167_a_80__dup_2309), 
                     .B (modgen_ram_ix167_a_82__dup_2307), .C (
                     modgen_ram_ix167_a_81__dup_2308), .D (
                     modgen_ram_ix167_a_83__dup_2306), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix7083 (.Y (nx7082), .A (modgen_ram_ix167_a_88__dup_2301), 
                     .B (modgen_ram_ix167_a_90__dup_2299), .C (
                     modgen_ram_ix167_a_89__dup_2300), .D (
                     modgen_ram_ix167_a_91__dup_2298), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix7027 (.Y (nx7026), .A (modgen_ram_ix167_a_84__dup_2305), 
                     .B (modgen_ram_ix167_a_86__dup_2303), .C (
                     modgen_ram_ix167_a_85__dup_2304), .D (
                     modgen_ram_ix167_a_87__dup_2302), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2677 (.Y (nx3272), .A (modgen_ram_ix167_a_92__dup_2297), 
                     .B (modgen_ram_ix167_a_94__dup_2295), .C (
                     modgen_ram_ix167_a_93__dup_2296), .D (
                     modgen_ram_ix167_a_95__dup_2294), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6927 (.Y (nx6926), .A0 (rd_addr_m_3), .A1 (nx3337), 
                          .B0 (nx1315), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2679 (.Y (nx3337), .A0 (rd_addr_m_2), .A1 (nx6806), .B0 (
                      nx6758)) ;
    MXT4_X0P5M_A12TS ix6807 (.Y (nx6806), .A (modgen_ram_ix167_a_68__dup_2321), 
                     .B (modgen_ram_ix167_a_70__dup_2319), .C (
                     modgen_ram_ix167_a_69__dup_2320), .D (
                     modgen_ram_ix167_a_71__dup_2318), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6759 (.Y (nx6758), .A0 (rd_addr_m_1), .A1 (nx1309), 
                          .B0 (nx1311), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2681 (.Y (nx1309), .A (modgen_ram_ix167_a_64__dup_2325)
                      , .B (modgen_ram_ix167_a_65__dup_2324), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2683 (.Y (nx1311), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_2322), .B0 (nx6740), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix6741 (.Y (nx6740), .AN (modgen_ram_ix167_a_66__dup_2323)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2684 (.Y (nx1315), .A0 (rd_addr_m_2), .A1 (nx3271), 
                          .B0 (nx6866), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix2686 (.Y (nx3271), .A (modgen_ram_ix167_a_76__dup_2313), 
                     .B (modgen_ram_ix167_a_78__dup_2311), .C (
                     modgen_ram_ix167_a_77__dup_2312), .D (
                     modgen_ram_ix167_a_79__dup_2310), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6867 (.Y (nx6866), .A0 (rd_addr_m_1), .A1 (nx1321), 
                          .B0 (nx1323), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2688 (.Y (nx1321), .A (modgen_ram_ix167_a_72__dup_2317)
                      , .B (modgen_ram_ix167_a_73__dup_2316), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2690 (.Y (nx1323), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_2314), .B0 (nx6848), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix6849 (.Y (nx6848), .AN (modgen_ram_ix167_a_74__dup_2315)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2691 (.Y (nx1326), .A0 (rd_addr_m_4), .A1 (nx3275), 
                          .B0 (nx7370), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix2692 (.Y (nx3275), .A (nx7418), .B (nx3273), .C (nx7470)
                     , .D (nx7578), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix7419 (.Y (nx7418), .A (modgen_ram_ix167_a_112__dup_2277)
                     , .B (modgen_ram_ix167_a_114__dup_2275), .C (
                     modgen_ram_ix167_a_113__dup_2276), .D (
                     modgen_ram_ix167_a_115__dup_2274), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2694 (.Y (nx3273), .A (modgen_ram_ix167_a_120__dup_2269)
                     , .B (modgen_ram_ix167_a_122__dup_2267), .C (
                     modgen_ram_ix167_a_121__dup_2268), .D (
                     modgen_ram_ix167_a_123__dup_2266), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix7471 (.Y (nx7470), .A (modgen_ram_ix167_a_116__dup_2273)
                     , .B (modgen_ram_ix167_a_118__dup_2271), .C (
                     modgen_ram_ix167_a_117__dup_2272), .D (
                     modgen_ram_ix167_a_119__dup_2270), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix7579 (.Y (nx7578), .A (modgen_ram_ix167_a_124__dup_2265)
                     , .B (modgen_ram_ix167_a_126__dup_2263), .C (
                     modgen_ram_ix167_a_125__dup_2264), .D (
                     modgen_ram_ix167_a_127__dup_2262), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix7371 (.Y (nx7370), .A0 (rd_addr_m_3), .A1 (nx1335), 
                          .B0 (nx1344), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2696 (.Y (nx1335), .A0 (rd_addr_m_2), .A1 (nx7250), .B0 (
                      nx7202)) ;
    MXT4_X0P5M_A12TS ix7251 (.Y (nx7250), .A (modgen_ram_ix167_a_100__dup_2289)
                     , .B (modgen_ram_ix167_a_102__dup_2287), .C (
                     modgen_ram_ix167_a_101__dup_2288), .D (
                     modgen_ram_ix167_a_103__dup_2286), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix7203 (.Y (nx7202), .A0 (rd_addr_m_1), .A1 (nx1339), 
                          .B0 (nx1341), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2698 (.Y (nx1339), .A (modgen_ram_ix167_a_96__dup_2293)
                      , .B (modgen_ram_ix167_a_97__dup_2292), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2700 (.Y (nx1341), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_2290), .B0 (nx7184), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix7185 (.Y (nx7184), .AN (modgen_ram_ix167_a_98__dup_2291)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2702 (.Y (nx1344), .A0 (rd_addr_m_2), .A1 (nx7358), 
                          .B0 (nx7310), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix7359 (.Y (nx7358), .A (modgen_ram_ix167_a_108__dup_2281)
                     , .B (modgen_ram_ix167_a_110__dup_2279), .C (
                     modgen_ram_ix167_a_109__dup_2280), .D (
                     modgen_ram_ix167_a_111__dup_2278), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix7311 (.Y (nx7310), .A0 (rd_addr_m_1), .A1 (nx1349), 
                          .B0 (nx1351), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2704 (.Y (nx1349), .A (modgen_ram_ix167_a_104__dup_2285)
                      , .B (modgen_ram_ix167_a_105__dup_2284), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2706 (.Y (nx1351), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_2282), .B0 (nx7292), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix7293 (.Y (nx7292), .AN (modgen_ram_ix167_a_106__dup_2283
                      ), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6707 (.Y (nx6706), .A0 (rd_addr_m_5), .A1 (nx1357), 
                          .B0 (nx1389), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2707 (.Y (nx1357), .A0 (rd_addr_m_4), .A1 (nx6250), .B0 (
                      nx3269)) ;
    MXT4_X0P5M_A12TS ix6251 (.Y (nx6250), .A (nx6082), .B (nx6190), .C (nx3270)
                     , .D (nx6242), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix6083 (.Y (nx6082), .A (modgen_ram_ix167_a_16__dup_2373), 
                     .B (modgen_ram_ix167_a_18__dup_2371), .C (
                     modgen_ram_ix167_a_17__dup_2372), .D (
                     modgen_ram_ix167_a_19__dup_2370), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix6191 (.Y (nx6190), .A (modgen_ram_ix167_a_24__dup_2365), 
                     .B (modgen_ram_ix167_a_26__dup_2363), .C (
                     modgen_ram_ix167_a_25__dup_2364), .D (
                     modgen_ram_ix167_a_27__dup_2362), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix2709 (.Y (nx3270), .A (modgen_ram_ix167_a_20__dup_2369), 
                     .B (modgen_ram_ix167_a_22__dup_2367), .C (
                     modgen_ram_ix167_a_21__dup_2368), .D (
                     modgen_ram_ix167_a_23__dup_2366), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix6243 (.Y (nx6242), .A (modgen_ram_ix167_a_28__dup_2361), 
                     .B (modgen_ram_ix167_a_30__dup_2359), .C (
                     modgen_ram_ix167_a_29__dup_2360), .D (
                     modgen_ram_ix167_a_31__dup_2358), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2713 (.Y (nx3269), .A0 (rd_addr_m_3), .A1 (nx1367), 
                          .B0 (nx1377), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1368 (.Y (nx1367), .A0 (rd_addr_m_2), .A1 (nx3267), .B0 (
                      nx5866)) ;
    MXT4_X0P5M_A12TS ix2714 (.Y (nx3267), .A (modgen_ram_ix167_a_4__dup_2385), .B (
                     modgen_ram_ix167_a_6__dup_2383), .C (
                     modgen_ram_ix167_a_5__dup_2384), .D (
                     modgen_ram_ix167_a_7__dup_2382), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix5867 (.Y (nx5866), .A0 (rd_addr_m_1), .A1 (nx3339), 
                          .B0 (nx1374), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2716 (.Y (nx3339), .A (modgen_ram_ix167_a_0__dup_2389), 
                      .B (modgen_ram_ix167_a_1__dup_2388), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2718 (.Y (nx1374), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_2386), .B0 (nx5848), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix5849 (.Y (nx5848), .AN (modgen_ram_ix167_a_2__dup_2387)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1378 (.Y (nx1377), .A0 (rd_addr_m_2), .A1 (nx6022), 
                          .B0 (nx3268), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix6023 (.Y (nx6022), .A (modgen_ram_ix167_a_12__dup_2377), 
                     .B (modgen_ram_ix167_a_14__dup_2375), .C (
                     modgen_ram_ix167_a_13__dup_2376), .D (
                     modgen_ram_ix167_a_15__dup_2374), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix2720 (.Y (nx3268), .A0 (rd_addr_m_1), .A1 (nx1383), 
                          .B0 (nx1385), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1384 (.Y (nx1383), .A (modgen_ram_ix167_a_8__dup_2381), 
                      .B (modgen_ram_ix167_a_9__dup_2380), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1386 (.Y (nx1385), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_2378), .B0 (nx5956), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix5957 (.Y (nx5956), .AN (modgen_ram_ix167_a_10__dup_2379)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1390 (.Y (nx1389), .A0 (rd_addr_m_4), .A1 (nx6694), 
                          .B0 (nx6478), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix6695 (.Y (nx6694), .A (nx6526), .B (nx6634), .C (nx6578)
                     , .D (nx6686), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix6527 (.Y (nx6526), .A (modgen_ram_ix167_a_48__dup_2341), 
                     .B (modgen_ram_ix167_a_50__dup_2339), .C (
                     modgen_ram_ix167_a_49__dup_2340), .D (
                     modgen_ram_ix167_a_51__dup_2338), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix6635 (.Y (nx6634), .A (modgen_ram_ix167_a_56__dup_2333), 
                     .B (modgen_ram_ix167_a_58__dup_2331), .C (
                     modgen_ram_ix167_a_57__dup_2332), .D (
                     modgen_ram_ix167_a_59__dup_2330), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix6579 (.Y (nx6578), .A (modgen_ram_ix167_a_52__dup_2337), 
                     .B (modgen_ram_ix167_a_54__dup_2335), .C (
                     modgen_ram_ix167_a_53__dup_2336), .D (
                     modgen_ram_ix167_a_55__dup_2334), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix6687 (.Y (nx6686), .A (modgen_ram_ix167_a_60__dup_2329), 
                     .B (modgen_ram_ix167_a_62__dup_2327), .C (
                     modgen_ram_ix167_a_61__dup_2328), .D (
                     modgen_ram_ix167_a_63__dup_2326), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6479 (.Y (nx6478), .A0 (rd_addr_m_3), .A1 (nx1399), 
                          .B0 (nx1411), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1400 (.Y (nx1399), .A0 (rd_addr_m_2), .A1 (nx6358), .B0 (
                      nx6310)) ;
    MXT4_X0P5M_A12TS ix6359 (.Y (nx6358), .A (modgen_ram_ix167_a_36__dup_2353), 
                     .B (modgen_ram_ix167_a_38__dup_2351), .C (
                     modgen_ram_ix167_a_37__dup_2352), .D (
                     modgen_ram_ix167_a_39__dup_2350), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6311 (.Y (nx6310), .A0 (rd_addr_m_1), .A1 (nx1405), 
                          .B0 (nx1407), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2721 (.Y (nx1405), .A (modgen_ram_ix167_a_32__dup_2357)
                      , .B (modgen_ram_ix167_a_33__dup_2356), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1408 (.Y (nx1407), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_2354), .B0 (nx6292), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix6293 (.Y (nx6292), .AN (modgen_ram_ix167_a_34__dup_2355)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1412 (.Y (nx1411), .A0 (rd_addr_m_2), .A1 (nx6466), 
                          .B0 (nx6418), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix6467 (.Y (nx6466), .A (modgen_ram_ix167_a_44__dup_2345), 
                     .B (modgen_ram_ix167_a_46__dup_2343), .C (
                     modgen_ram_ix167_a_45__dup_2344), .D (
                     modgen_ram_ix167_a_47__dup_2342), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix6419 (.Y (nx6418), .A0 (rd_addr_m_1), .A1 (nx1415), 
                          .B0 (nx1417), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1416 (.Y (nx1415), .A (modgen_ram_ix167_a_40__dup_2349)
                      , .B (modgen_ram_ix167_a_41__dup_2348), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1418 (.Y (nx1417), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_2346), .B0 (nx6400), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix6401 (.Y (nx6400), .AN (modgen_ram_ix167_a_42__dup_2347)
                      , .B (rd_addr_m_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_2 (.Q (rd_data_m_2), .CK (wb_clk_i), .D (
                        nx12986), .R (wb_rst_i), .SE (NOT_nx50), .SI (
                        rd_data_m_2)) ;
    MXIT2_X0P5M_A12TS ix12987 (.Y (nx12986), .A (nx1423), .B (nx1425), .S0 (
                      nx1127)) ;
    INV_X0P5B_A12TS ix1424 (.Y (nx1423), .A (wr_data_m_2)) ;
    OA21A1OI2_X0P5M_A12TS ix1426 (.Y (nx1425), .A0 (nx12972), .A1 (nx12082), .B0 (
                          rd_addr_7), .C0 (nx11190)) ;
    OA21A1OI2_X0P5M_A12TS ix12973 (.Y (nx12972), .A0 (rd_addr_m_5), .A1 (nx1429)
                          , .B0 (nx1461), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix1430 (.Y (nx1429), .A0 (rd_addr_m_4), .A1 (nx12518), .B0 (
                      nx12302)) ;
    MXT4_X0P5M_A12TS ix12519 (.Y (nx12518), .A (nx12350), .B (nx12458), .C (
                     nx12402), .D (nx12510), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix12351 (.Y (nx12350), .A (modgen_ram_ix167_a_208__dup_1917
                     ), .B (modgen_ram_ix167_a_210__dup_1915), .C (
                     modgen_ram_ix167_a_209__dup_1916), .D (
                     modgen_ram_ix167_a_211__dup_1914), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12459 (.Y (nx12458), .A (modgen_ram_ix167_a_216__dup_1909
                     ), .B (modgen_ram_ix167_a_218__dup_1907), .C (
                     modgen_ram_ix167_a_217__dup_1908), .D (
                     modgen_ram_ix167_a_219__dup_1906), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12403 (.Y (nx12402), .A (modgen_ram_ix167_a_212__dup_1913
                     ), .B (modgen_ram_ix167_a_214__dup_1911), .C (
                     modgen_ram_ix167_a_213__dup_1912), .D (
                     modgen_ram_ix167_a_215__dup_1910), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12511 (.Y (nx12510), .A (modgen_ram_ix167_a_220__dup_1905
                     ), .B (modgen_ram_ix167_a_222__dup_1903), .C (
                     modgen_ram_ix167_a_221__dup_1904), .D (
                     modgen_ram_ix167_a_223__dup_1902), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12303 (.Y (nx12302), .A0 (rd_addr_m_3), .A1 (nx1439)
                          , .B0 (nx1451), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1440 (.Y (nx1439), .A0 (rd_addr_m_2), .A1 (nx12182), .B0 (
                      nx12134)) ;
    MXT4_X0P5M_A12TS ix12183 (.Y (nx12182), .A (modgen_ram_ix167_a_196__dup_1929
                     ), .B (modgen_ram_ix167_a_198__dup_1927), .C (
                     modgen_ram_ix167_a_197__dup_1928), .D (
                     modgen_ram_ix167_a_199__dup_1926), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12135 (.Y (nx12134), .A0 (rd_addr_m_1), .A1 (nx1445)
                          , .B0 (nx1447), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1446 (.Y (nx1445), .A (modgen_ram_ix167_a_192__dup_1933)
                      , .B (modgen_ram_ix167_a_193__dup_1932), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1448 (.Y (nx1447), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_1930), .B0 (nx12116), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix12117 (.Y (nx12116), .AN (
                      modgen_ram_ix167_a_194__dup_1931), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1452 (.Y (nx1451), .A0 (rd_addr_m_2), .A1 (nx12290)
                          , .B0 (nx12242), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix12291 (.Y (nx12290), .A (modgen_ram_ix167_a_204__dup_1921
                     ), .B (modgen_ram_ix167_a_206__dup_1919), .C (
                     modgen_ram_ix167_a_205__dup_1920), .D (
                     modgen_ram_ix167_a_207__dup_1918), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12243 (.Y (nx12242), .A0 (rd_addr_m_1), .A1 (nx3340)
                          , .B0 (nx1458), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2722 (.Y (nx3340), .A (modgen_ram_ix167_a_200__dup_1925)
                      , .B (modgen_ram_ix167_a_201__dup_1924), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1459 (.Y (nx1458), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_1922), .B0 (nx12224), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix12225 (.Y (nx12224), .AN (
                      modgen_ram_ix167_a_202__dup_1923), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1462 (.Y (nx1461), .A0 (rd_addr_m_4), .A1 (nx12962)
                          , .B0 (nx12746), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix12963 (.Y (nx12962), .A (nx12794), .B (nx12902), .C (
                     nx12846), .D (nx12954), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix12795 (.Y (nx12794), .A (modgen_ram_ix167_a_240__dup_1885
                     ), .B (modgen_ram_ix167_a_242__dup_1883), .C (
                     modgen_ram_ix167_a_241__dup_1884), .D (
                     modgen_ram_ix167_a_243__dup_1882), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12903 (.Y (nx12902), .A (modgen_ram_ix167_a_248__dup_1877
                     ), .B (modgen_ram_ix167_a_250__dup_1875), .C (
                     modgen_ram_ix167_a_249__dup_1876), .D (
                     modgen_ram_ix167_a_251__dup_1874), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12847 (.Y (nx12846), .A (modgen_ram_ix167_a_244__dup_1881
                     ), .B (modgen_ram_ix167_a_246__dup_1879), .C (
                     modgen_ram_ix167_a_245__dup_1880), .D (
                     modgen_ram_ix167_a_247__dup_1878), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12955 (.Y (nx12954), .A (modgen_ram_ix167_a_252__dup_1873
                     ), .B (modgen_ram_ix167_a_254__dup_1871), .C (
                     modgen_ram_ix167_a_253__dup_1872), .D (
                     modgen_ram_ix167_a_255__dup_1870), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12747 (.Y (nx12746), .A0 (rd_addr_m_3), .A1 (nx3341)
                          , .B0 (nx3345), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1472 (.Y (nx3341), .A0 (rd_addr_m_2), .A1 (nx12626), .B0 (
                      nx12578)) ;
    MXT4_X0P5M_A12TS ix12627 (.Y (nx12626), .A (modgen_ram_ix167_a_228__dup_1897
                     ), .B (modgen_ram_ix167_a_230__dup_1895), .C (
                     modgen_ram_ix167_a_229__dup_1896), .D (
                     modgen_ram_ix167_a_231__dup_1894), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12579 (.Y (nx12578), .A0 (rd_addr_m_1), .A1 (nx3342)
                          , .B0 (nx3343), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1476 (.Y (nx3342), .A (modgen_ram_ix167_a_224__dup_1901)
                      , .B (modgen_ram_ix167_a_225__dup_1900), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1478 (.Y (nx3343), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_1898), .B0 (nx12560), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix12561 (.Y (nx12560), .AN (
                      modgen_ram_ix167_a_226__dup_1899), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1482 (.Y (nx3345), .A0 (rd_addr_m_2), .A1 (nx12734)
                          , .B0 (nx12686), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix12735 (.Y (nx12734), .A (modgen_ram_ix167_a_236__dup_1889
                     ), .B (modgen_ram_ix167_a_238__dup_1887), .C (
                     modgen_ram_ix167_a_237__dup_1888), .D (
                     modgen_ram_ix167_a_239__dup_1886), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12687 (.Y (nx12686), .A0 (rd_addr_m_1), .A1 (nx3346)
                          , .B0 (nx3347), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1486 (.Y (nx3346), .A (modgen_ram_ix167_a_232__dup_1893)
                      , .B (modgen_ram_ix167_a_233__dup_1892), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1488 (.Y (nx3347), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_1890), .B0 (nx12668), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix12669 (.Y (nx12668), .AN (
                      modgen_ram_ix167_a_234__dup_1891), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix12083 (.Y (nx12082), .A0 (rd_addr_m_5), .A1 (nx3348)
                          , .B0 (nx3355), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix1494 (.Y (nx3348), .A0 (rd_addr_m_4), .A1 (nx11626), .B0 (
                      nx11410)) ;
    MXT4_X0P5M_A12TS ix11627 (.Y (nx11626), .A (nx11458), .B (nx11566), .C (
                     nx11510), .D (nx11618), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix11459 (.Y (nx11458), .A (modgen_ram_ix167_a_144__dup_1981
                     ), .B (modgen_ram_ix167_a_146__dup_1979), .C (
                     modgen_ram_ix167_a_145__dup_1980), .D (
                     modgen_ram_ix167_a_147__dup_1978), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11567 (.Y (nx11566), .A (modgen_ram_ix167_a_152__dup_1973
                     ), .B (modgen_ram_ix167_a_154__dup_1971), .C (
                     modgen_ram_ix167_a_153__dup_1972), .D (
                     modgen_ram_ix167_a_155__dup_1970), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11511 (.Y (nx11510), .A (modgen_ram_ix167_a_148__dup_1977
                     ), .B (modgen_ram_ix167_a_150__dup_1975), .C (
                     modgen_ram_ix167_a_149__dup_1976), .D (
                     modgen_ram_ix167_a_151__dup_1974), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11619 (.Y (nx11618), .A (modgen_ram_ix167_a_156__dup_1969
                     ), .B (modgen_ram_ix167_a_158__dup_1967), .C (
                     modgen_ram_ix167_a_157__dup_1968), .D (
                     modgen_ram_ix167_a_159__dup_1966), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix11411 (.Y (nx11410), .A0 (rd_addr_m_3), .A1 (nx3349)
                          , .B0 (nx3352), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2724 (.Y (nx3349), .A0 (rd_addr_m_2), .A1 (nx11290), .B0 (
                      nx11242)) ;
    MXT4_X0P5M_A12TS ix11291 (.Y (nx11290), .A (modgen_ram_ix167_a_132__dup_1993
                     ), .B (modgen_ram_ix167_a_134__dup_1991), .C (
                     modgen_ram_ix167_a_133__dup_1992), .D (
                     modgen_ram_ix167_a_135__dup_1990), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix11243 (.Y (nx11242), .A0 (rd_addr_m_1), .A1 (nx3350)
                          , .B0 (nx3351), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1508 (.Y (nx3350), .A (modgen_ram_ix167_a_128__dup_1997)
                      , .B (modgen_ram_ix167_a_129__dup_1996), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2726 (.Y (nx3351), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_1994), .B0 (nx11224), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix11225 (.Y (nx11224), .AN (
                      modgen_ram_ix167_a_130__dup_1995), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2728 (.Y (nx3352), .A0 (rd_addr_m_2), .A1 (nx11398)
                          , .B0 (nx11350), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix11399 (.Y (nx11398), .A (modgen_ram_ix167_a_140__dup_1985
                     ), .B (modgen_ram_ix167_a_142__dup_1983), .C (
                     modgen_ram_ix167_a_141__dup_1984), .D (
                     modgen_ram_ix167_a_143__dup_1982), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix11351 (.Y (nx11350), .A0 (rd_addr_m_1), .A1 (nx3353)
                          , .B0 (nx3354), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1518 (.Y (nx3353), .A (modgen_ram_ix167_a_136__dup_1989)
                      , .B (modgen_ram_ix167_a_137__dup_1988), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2730 (.Y (nx3354), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_1986), .B0 (nx11332), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix11333 (.Y (nx11332), .AN (
                      modgen_ram_ix167_a_138__dup_1987), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2732 (.Y (nx3355), .A0 (rd_addr_m_4), .A1 (nx12070)
                          , .B0 (nx11854), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix12071 (.Y (nx12070), .A (nx11902), .B (nx12010), .C (
                     nx11954), .D (nx12062), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix11903 (.Y (nx11902), .A (modgen_ram_ix167_a_176__dup_1949
                     ), .B (modgen_ram_ix167_a_178__dup_1947), .C (
                     modgen_ram_ix167_a_177__dup_1948), .D (
                     modgen_ram_ix167_a_179__dup_1946), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12011 (.Y (nx12010), .A (modgen_ram_ix167_a_184__dup_1941
                     ), .B (modgen_ram_ix167_a_186__dup_1939), .C (
                     modgen_ram_ix167_a_185__dup_1940), .D (
                     modgen_ram_ix167_a_187__dup_1938), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11955 (.Y (nx11954), .A (modgen_ram_ix167_a_180__dup_1945
                     ), .B (modgen_ram_ix167_a_182__dup_1943), .C (
                     modgen_ram_ix167_a_181__dup_1944), .D (
                     modgen_ram_ix167_a_183__dup_1942), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix12063 (.Y (nx12062), .A (modgen_ram_ix167_a_188__dup_1937
                     ), .B (modgen_ram_ix167_a_190__dup_1935), .C (
                     modgen_ram_ix167_a_189__dup_1936), .D (
                     modgen_ram_ix167_a_191__dup_1934), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix11855 (.Y (nx11854), .A0 (rd_addr_m_3), .A1 (nx3356)
                          , .B0 (nx1549), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2734 (.Y (nx3356), .A0 (rd_addr_m_2), .A1 (nx11734), .B0 (
                      nx11686)) ;
    MXT4_X0P5M_A12TS ix11735 (.Y (nx11734), .A (modgen_ram_ix167_a_164__dup_1961
                     ), .B (modgen_ram_ix167_a_166__dup_1959), .C (
                     modgen_ram_ix167_a_165__dup_1960), .D (
                     modgen_ram_ix167_a_167__dup_1958), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix11687 (.Y (nx11686), .A0 (rd_addr_m_1), .A1 (nx3357)
                          , .B0 (nx1545), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2736 (.Y (nx3357), .A (modgen_ram_ix167_a_160__dup_1965)
                      , .B (modgen_ram_ix167_a_161__dup_1964), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2737 (.Y (nx1545), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_1962), .B0 (nx11668), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix11669 (.Y (nx11668), .AN (
                      modgen_ram_ix167_a_162__dup_1963), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2739 (.Y (nx1549), .A0 (rd_addr_m_2), .A1 (nx11842)
                          , .B0 (nx11794), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix11843 (.Y (nx11842), .A (modgen_ram_ix167_a_172__dup_1953
                     ), .B (modgen_ram_ix167_a_174__dup_1951), .C (
                     modgen_ram_ix167_a_173__dup_1952), .D (
                     modgen_ram_ix167_a_175__dup_1950), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix11795 (.Y (nx11794), .A0 (rd_addr_m_1), .A1 (nx1555)
                          , .B0 (nx3358), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2741 (.Y (nx1555), .A (modgen_ram_ix167_a_168__dup_1957)
                      , .B (modgen_ram_ix167_a_169__dup_1956), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2743 (.Y (nx3358), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_1954), .B0 (nx11776), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix11777 (.Y (nx11776), .AN (
                      modgen_ram_ix167_a_170__dup_1955), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix11191 (.Y (nx11190), .A (rd_addr_7), .B (nx1562)) ;
    AOI21_X0P5M_A12TS ix2744 (.Y (nx1562), .A0 (rd_addr_m_6), .A1 (nx11182), .B0 (
                      nx10294)) ;
    OAI21_X0P5M_A12TS ix11183 (.Y (nx11182), .A0 (rd_addr_m_5), .A1 (nx3359), .B0 (
                      nx1597)) ;
    AOI21_X0P5M_A12TS ix2746 (.Y (nx3359), .A0 (rd_addr_m_4), .A1 (nx10730), .B0 (
                      nx10514)) ;
    MXT4_X0P5M_A12TS ix10731 (.Y (nx10730), .A (nx10562), .B (nx10670), .C (
                     nx10614), .D (nx10722), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix10563 (.Y (nx10562), .A (modgen_ram_ix167_a_80__dup_2045)
                     , .B (modgen_ram_ix167_a_82__dup_2043), .C (
                     modgen_ram_ix167_a_81__dup_2044), .D (
                     modgen_ram_ix167_a_83__dup_2042), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix10671 (.Y (nx10670), .A (modgen_ram_ix167_a_88__dup_2037)
                     , .B (modgen_ram_ix167_a_90__dup_2035), .C (
                     modgen_ram_ix167_a_89__dup_2036), .D (
                     modgen_ram_ix167_a_91__dup_2034), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix10615 (.Y (nx10614), .A (modgen_ram_ix167_a_84__dup_2041)
                     , .B (modgen_ram_ix167_a_86__dup_2039), .C (
                     modgen_ram_ix167_a_85__dup_2040), .D (
                     modgen_ram_ix167_a_87__dup_2038), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix10723 (.Y (nx10722), .A (modgen_ram_ix167_a_92__dup_2033)
                     , .B (modgen_ram_ix167_a_94__dup_2031), .C (
                     modgen_ram_ix167_a_93__dup_2032), .D (
                     modgen_ram_ix167_a_95__dup_2030), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10515 (.Y (nx10514), .A0 (rd_addr_m_3), .A1 (nx1575)
                          , .B0 (nx3362), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2748 (.Y (nx1575), .A0 (rd_addr_m_2), .A1 (nx10394), .B0 (
                      nx10346)) ;
    MXT4_X0P5M_A12TS ix10395 (.Y (nx10394), .A (modgen_ram_ix167_a_68__dup_2057)
                     , .B (modgen_ram_ix167_a_70__dup_2055), .C (
                     modgen_ram_ix167_a_69__dup_2056), .D (
                     modgen_ram_ix167_a_71__dup_2054), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10347 (.Y (nx10346), .A0 (rd_addr_m_1), .A1 (nx3361)
                          , .B0 (nx1582), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2750 (.Y (nx3361), .A (modgen_ram_ix167_a_64__dup_2061)
                      , .B (modgen_ram_ix167_a_65__dup_2060), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2751 (.Y (nx1582), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_2058), .B0 (nx10328), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix10329 (.Y (nx10328), .AN (
                      modgen_ram_ix167_a_66__dup_2059), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2752 (.Y (nx3362), .A0 (rd_addr_m_2), .A1 (nx10502)
                          , .B0 (nx10454), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix10503 (.Y (nx10502), .A (modgen_ram_ix167_a_76__dup_2049)
                     , .B (modgen_ram_ix167_a_78__dup_2047), .C (
                     modgen_ram_ix167_a_77__dup_2048), .D (
                     modgen_ram_ix167_a_79__dup_2046), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10455 (.Y (nx10454), .A0 (rd_addr_m_1), .A1 (nx3363)
                          , .B0 (nx3364), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2753 (.Y (nx3363), .A (modgen_ram_ix167_a_72__dup_2053)
                      , .B (modgen_ram_ix167_a_73__dup_2052), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2754 (.Y (nx3364), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_2050), .B0 (nx10436), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix10437 (.Y (nx10436), .AN (
                      modgen_ram_ix167_a_74__dup_2051), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2756 (.Y (nx1597), .A0 (rd_addr_m_4), .A1 (nx11174)
                          , .B0 (nx10958), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix11175 (.Y (nx11174), .A (nx11006), .B (nx11114), .C (
                     nx11058), .D (nx11166), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix11007 (.Y (nx11006), .A (modgen_ram_ix167_a_112__dup_2013
                     ), .B (modgen_ram_ix167_a_114__dup_2011), .C (
                     modgen_ram_ix167_a_113__dup_2012), .D (
                     modgen_ram_ix167_a_115__dup_2010), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11115 (.Y (nx11114), .A (modgen_ram_ix167_a_120__dup_2005
                     ), .B (modgen_ram_ix167_a_122__dup_2003), .C (
                     modgen_ram_ix167_a_121__dup_2004), .D (
                     modgen_ram_ix167_a_123__dup_2002), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11059 (.Y (nx11058), .A (modgen_ram_ix167_a_116__dup_2009
                     ), .B (modgen_ram_ix167_a_118__dup_2007), .C (
                     modgen_ram_ix167_a_117__dup_2008), .D (
                     modgen_ram_ix167_a_119__dup_2006), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix11167 (.Y (nx11166), .A (modgen_ram_ix167_a_124__dup_2001
                     ), .B (modgen_ram_ix167_a_126__dup_1999), .C (
                     modgen_ram_ix167_a_125__dup_2000), .D (
                     modgen_ram_ix167_a_127__dup_1998), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10959 (.Y (nx10958), .A0 (rd_addr_m_3), .A1 (nx1606)
                          , .B0 (nx1617), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2757 (.Y (nx1606), .A0 (rd_addr_m_2), .A1 (nx10838), .B0 (
                      nx10790)) ;
    MXT4_X0P5M_A12TS ix10839 (.Y (nx10838), .A (modgen_ram_ix167_a_100__dup_2025
                     ), .B (modgen_ram_ix167_a_102__dup_2023), .C (
                     modgen_ram_ix167_a_101__dup_2024), .D (
                     modgen_ram_ix167_a_103__dup_2022), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10791 (.Y (nx10790), .A0 (rd_addr_m_1), .A1 (nx3365)
                          , .B0 (nx1613), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2758 (.Y (nx3365), .A (modgen_ram_ix167_a_96__dup_2029)
                      , .B (modgen_ram_ix167_a_97__dup_2028), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2759 (.Y (nx1613), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_2026), .B0 (nx10772), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix10773 (.Y (nx10772), .AN (
                      modgen_ram_ix167_a_98__dup_2027), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2760 (.Y (nx1617), .A0 (rd_addr_m_2), .A1 (nx10946)
                          , .B0 (nx10898), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix10947 (.Y (nx10946), .A (modgen_ram_ix167_a_108__dup_2017
                     ), .B (modgen_ram_ix167_a_110__dup_2015), .C (
                     modgen_ram_ix167_a_109__dup_2016), .D (
                     modgen_ram_ix167_a_111__dup_2014), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10899 (.Y (nx10898), .A0 (rd_addr_m_1), .A1 (nx1621)
                          , .B0 (nx3366), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2761 (.Y (nx1621), .A (modgen_ram_ix167_a_104__dup_2021)
                      , .B (modgen_ram_ix167_a_105__dup_2020), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2762 (.Y (nx3366), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_2018), .B0 (nx10880), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix10881 (.Y (nx10880), .AN (
                      modgen_ram_ix167_a_106__dup_2019), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10295 (.Y (nx10294), .A0 (rd_addr_m_5), .A1 (nx3367)
                          , .B0 (nx1659), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2763 (.Y (nx3367), .A0 (rd_addr_m_4), .A1 (nx9838), .B0 (
                      nx9622)) ;
    MXT4_X0P5M_A12TS ix9839 (.Y (nx9838), .A (nx9670), .B (nx9778), .C (nx9722)
                     , .D (nx9830), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2)) ;
    MXT4_X0P5M_A12TS ix9671 (.Y (nx9670), .A (modgen_ram_ix167_a_16__dup_2109), 
                     .B (modgen_ram_ix167_a_18__dup_2107), .C (
                     modgen_ram_ix167_a_17__dup_2108), .D (
                     modgen_ram_ix167_a_19__dup_2106), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix9779 (.Y (nx9778), .A (modgen_ram_ix167_a_24__dup_2101), 
                     .B (modgen_ram_ix167_a_26__dup_2099), .C (
                     modgen_ram_ix167_a_25__dup_2100), .D (
                     modgen_ram_ix167_a_27__dup_2098), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix9723 (.Y (nx9722), .A (modgen_ram_ix167_a_20__dup_2105), 
                     .B (modgen_ram_ix167_a_22__dup_2103), .C (
                     modgen_ram_ix167_a_21__dup_2104), .D (
                     modgen_ram_ix167_a_23__dup_2102), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix9831 (.Y (nx9830), .A (modgen_ram_ix167_a_28__dup_2097), 
                     .B (modgen_ram_ix167_a_30__dup_2095), .C (
                     modgen_ram_ix167_a_29__dup_2096), .D (
                     modgen_ram_ix167_a_31__dup_2094), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix9623 (.Y (nx9622), .A0 (rd_addr_m_3), .A1 (nx3369), 
                          .B0 (nx1648), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2764 (.Y (nx3369), .A0 (rd_addr_m_2), .A1 (nx9502), .B0 (
                      nx9454)) ;
    MXT4_X0P5M_A12TS ix9503 (.Y (nx9502), .A (modgen_ram_ix167_a_4__dup_2121), .B (
                     modgen_ram_ix167_a_6__dup_2119), .C (
                     modgen_ram_ix167_a_5__dup_2120), .D (
                     modgen_ram_ix167_a_7__dup_2118), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix9455 (.Y (nx9454), .A0 (rd_addr_m_1), .A1 (nx3370), 
                          .B0 (nx3371), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2765 (.Y (nx3370), .A (modgen_ram_ix167_a_0__dup_2125), 
                      .B (modgen_ram_ix167_a_1__dup_2124), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2766 (.Y (nx3371), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_2122), .B0 (nx9436), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix9437 (.Y (nx9436), .AN (modgen_ram_ix167_a_2__dup_2123)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2767 (.Y (nx1648), .A0 (rd_addr_m_2), .A1 (nx9610), 
                          .B0 (nx9562), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix9611 (.Y (nx9610), .A (modgen_ram_ix167_a_12__dup_2113), 
                     .B (modgen_ram_ix167_a_14__dup_2111), .C (
                     modgen_ram_ix167_a_13__dup_2112), .D (
                     modgen_ram_ix167_a_15__dup_2110), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix9563 (.Y (nx9562), .A0 (rd_addr_m_1), .A1 (nx3372), 
                          .B0 (nx1655), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2768 (.Y (nx3372), .A (modgen_ram_ix167_a_8__dup_2117), 
                      .B (modgen_ram_ix167_a_9__dup_2116), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2770 (.Y (nx1655), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_2114), .B0 (nx9544), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix9545 (.Y (nx9544), .AN (modgen_ram_ix167_a_10__dup_2115)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2772 (.Y (nx1659), .A0 (rd_addr_m_4), .A1 (nx10282)
                          , .B0 (nx10066), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix10283 (.Y (nx10282), .A (nx10114), .B (nx10222), .C (
                     nx10166), .D (nx10274), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix10115 (.Y (nx10114), .A (modgen_ram_ix167_a_48__dup_2077)
                     , .B (modgen_ram_ix167_a_50__dup_2075), .C (
                     modgen_ram_ix167_a_49__dup_2076), .D (
                     modgen_ram_ix167_a_51__dup_2074), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix10223 (.Y (nx10222), .A (modgen_ram_ix167_a_56__dup_2069)
                     , .B (modgen_ram_ix167_a_58__dup_2067), .C (
                     modgen_ram_ix167_a_57__dup_2068), .D (
                     modgen_ram_ix167_a_59__dup_2066), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix10167 (.Y (nx10166), .A (modgen_ram_ix167_a_52__dup_2073)
                     , .B (modgen_ram_ix167_a_54__dup_2071), .C (
                     modgen_ram_ix167_a_53__dup_2072), .D (
                     modgen_ram_ix167_a_55__dup_2070), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix10275 (.Y (nx10274), .A (modgen_ram_ix167_a_60__dup_2065)
                     , .B (modgen_ram_ix167_a_62__dup_2063), .C (
                     modgen_ram_ix167_a_61__dup_2064), .D (
                     modgen_ram_ix167_a_63__dup_2062), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10067 (.Y (nx10066), .A0 (rd_addr_m_3), .A1 (nx1669)
                          , .B0 (nx3373), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2773 (.Y (nx1669), .A0 (rd_addr_m_2), .A1 (nx9946), .B0 (
                      nx9898)) ;
    MXT4_X0P5M_A12TS ix9947 (.Y (nx9946), .A (modgen_ram_ix167_a_36__dup_2089), 
                     .B (modgen_ram_ix167_a_38__dup_2087), .C (
                     modgen_ram_ix167_a_37__dup_2088), .D (
                     modgen_ram_ix167_a_39__dup_2086), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix9899 (.Y (nx9898), .A0 (rd_addr_m_1), .A1 (nx1675), 
                          .B0 (nx1677), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2774 (.Y (nx1675), .A (modgen_ram_ix167_a_32__dup_2093)
                      , .B (modgen_ram_ix167_a_33__dup_2092), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2775 (.Y (nx1677), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_2090), .B0 (nx9880), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix9881 (.Y (nx9880), .AN (modgen_ram_ix167_a_34__dup_2091)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2776 (.Y (nx3373), .A0 (rd_addr_m_2), .A1 (nx10054)
                          , .B0 (nx10006), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix10055 (.Y (nx10054), .A (modgen_ram_ix167_a_44__dup_2081)
                     , .B (modgen_ram_ix167_a_46__dup_2079), .C (
                     modgen_ram_ix167_a_45__dup_2080), .D (
                     modgen_ram_ix167_a_47__dup_2078), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix10007 (.Y (nx10006), .A0 (rd_addr_m_1), .A1 (nx1686)
                          , .B0 (nx1688), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2777 (.Y (nx1686), .A (modgen_ram_ix167_a_40__dup_2085)
                      , .B (modgen_ram_ix167_a_41__dup_2084), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2778 (.Y (nx1688), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_2082), .B0 (nx9988), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix9989 (.Y (nx9988), .AN (modgen_ram_ix167_a_42__dup_2083)
                      , .B (rd_addr_m_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_3 (.Q (rd_data_m_3), .CK (wb_clk_i), .D (
                        nx16574), .R (wb_rst_i), .SE (NOT_nx50), .SI (
                        rd_data_m_3)) ;
    MXIT2_X0P5M_A12TS ix16575 (.Y (nx16574), .A (nx3374), .B (nx1695), .S0 (
                      nx1127)) ;
    INV_X0P5B_A12TS ix2779 (.Y (nx3374), .A (wr_data_m_3)) ;
    OA21A1OI2_X0P5M_A12TS ix2780 (.Y (nx1695), .A0 (nx16560), .A1 (nx15670), .B0 (
                          rd_addr_7), .C0 (nx14778)) ;
    OA21A1OI2_X0P5M_A12TS ix16561 (.Y (nx16560), .A0 (rd_addr_m_5), .A1 (nx1699)
                          , .B0 (nx3377), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2781 (.Y (nx1699), .A0 (rd_addr_m_4), .A1 (nx16106), .B0 (
                      nx15890)) ;
    MXT4_X0P5M_A12TS ix16107 (.Y (nx16106), .A (nx15938), .B (nx16046), .C (
                     nx15990), .D (nx16098), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix15939 (.Y (nx15938), .A (modgen_ram_ix167_a_208__dup_1653
                     ), .B (modgen_ram_ix167_a_210__dup_1651), .C (
                     modgen_ram_ix167_a_209__dup_1652), .D (
                     modgen_ram_ix167_a_211__dup_1650), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16047 (.Y (nx16046), .A (modgen_ram_ix167_a_216__dup_1645
                     ), .B (modgen_ram_ix167_a_218__dup_1643), .C (
                     modgen_ram_ix167_a_217__dup_1644), .D (
                     modgen_ram_ix167_a_219__dup_1642), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15991 (.Y (nx15990), .A (modgen_ram_ix167_a_212__dup_1649
                     ), .B (modgen_ram_ix167_a_214__dup_1647), .C (
                     modgen_ram_ix167_a_213__dup_1648), .D (
                     modgen_ram_ix167_a_215__dup_1646), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16099 (.Y (nx16098), .A (modgen_ram_ix167_a_220__dup_1641
                     ), .B (modgen_ram_ix167_a_222__dup_1639), .C (
                     modgen_ram_ix167_a_221__dup_1640), .D (
                     modgen_ram_ix167_a_223__dup_1638), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15891 (.Y (nx15890), .A0 (rd_addr_m_3), .A1 (nx1709)
                          , .B0 (nx1721), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2782 (.Y (nx1709), .A0 (rd_addr_m_2), .A1 (nx15770), .B0 (
                      nx15722)) ;
    MXT4_X0P5M_A12TS ix15771 (.Y (nx15770), .A (modgen_ram_ix167_a_196__dup_1665
                     ), .B (modgen_ram_ix167_a_198__dup_1663), .C (
                     modgen_ram_ix167_a_197__dup_1664), .D (
                     modgen_ram_ix167_a_199__dup_1662), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15723 (.Y (nx15722), .A0 (rd_addr_m_1), .A1 (nx1715)
                          , .B0 (nx1717), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1716 (.Y (nx1715), .A (modgen_ram_ix167_a_192__dup_1669)
                      , .B (modgen_ram_ix167_a_193__dup_1668), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1718 (.Y (nx1717), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_1666), .B0 (nx15704), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix15705 (.Y (nx15704), .AN (
                      modgen_ram_ix167_a_194__dup_1667), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1722 (.Y (nx1721), .A0 (rd_addr_m_2), .A1 (nx15878)
                          , .B0 (nx15830), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix15879 (.Y (nx15878), .A (modgen_ram_ix167_a_204__dup_1657
                     ), .B (modgen_ram_ix167_a_206__dup_1655), .C (
                     modgen_ram_ix167_a_205__dup_1656), .D (
                     modgen_ram_ix167_a_207__dup_1654), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15831 (.Y (nx15830), .A0 (rd_addr_m_1), .A1 (nx3375)
                          , .B0 (nx1729), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2783 (.Y (nx3375), .A (modgen_ram_ix167_a_200__dup_1661)
                      , .B (modgen_ram_ix167_a_201__dup_1660), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1730 (.Y (nx1729), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_1658), .B0 (nx15812), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix15813 (.Y (nx15812), .AN (
                      modgen_ram_ix167_a_202__dup_1659), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2784 (.Y (nx3377), .A0 (rd_addr_m_4), .A1 (nx16550)
                          , .B0 (nx16334), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix16551 (.Y (nx16550), .A (nx16382), .B (nx16490), .C (
                     nx16434), .D (nx16542), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix16383 (.Y (nx16382), .A (modgen_ram_ix167_a_240__dup_1621
                     ), .B (modgen_ram_ix167_a_242__dup_1619), .C (
                     modgen_ram_ix167_a_241__dup_1620), .D (
                     modgen_ram_ix167_a_243__dup_1618), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16491 (.Y (nx16490), .A (modgen_ram_ix167_a_248__dup_1613
                     ), .B (modgen_ram_ix167_a_250__dup_1611), .C (
                     modgen_ram_ix167_a_249__dup_1612), .D (
                     modgen_ram_ix167_a_251__dup_1610), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16435 (.Y (nx16434), .A (modgen_ram_ix167_a_244__dup_1617
                     ), .B (modgen_ram_ix167_a_246__dup_1615), .C (
                     modgen_ram_ix167_a_245__dup_1616), .D (
                     modgen_ram_ix167_a_247__dup_1614), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16543 (.Y (nx16542), .A (modgen_ram_ix167_a_252__dup_1609
                     ), .B (modgen_ram_ix167_a_254__dup_1607), .C (
                     modgen_ram_ix167_a_253__dup_1608), .D (
                     modgen_ram_ix167_a_255__dup_1606), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix16335 (.Y (nx16334), .A0 (rd_addr_m_3), .A1 (nx1741)
                          , .B0 (nx1751), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1742 (.Y (nx1741), .A0 (rd_addr_m_2), .A1 (nx16214), .B0 (
                      nx16166)) ;
    MXT4_X0P5M_A12TS ix16215 (.Y (nx16214), .A (modgen_ram_ix167_a_228__dup_1633
                     ), .B (modgen_ram_ix167_a_230__dup_1631), .C (
                     modgen_ram_ix167_a_229__dup_1632), .D (
                     modgen_ram_ix167_a_231__dup_1630), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix16167 (.Y (nx16166), .A0 (rd_addr_m_1), .A1 (nx1745)
                          , .B0 (nx1747), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1746 (.Y (nx1745), .A (modgen_ram_ix167_a_224__dup_1637)
                      , .B (modgen_ram_ix167_a_225__dup_1636), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1748 (.Y (nx1747), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_1634), .B0 (nx16148), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix16149 (.Y (nx16148), .AN (
                      modgen_ram_ix167_a_226__dup_1635), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1752 (.Y (nx1751), .A0 (rd_addr_m_2), .A1 (nx16322)
                          , .B0 (nx16274), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix16323 (.Y (nx16322), .A (modgen_ram_ix167_a_236__dup_1625
                     ), .B (modgen_ram_ix167_a_238__dup_1623), .C (
                     modgen_ram_ix167_a_237__dup_1624), .D (
                     modgen_ram_ix167_a_239__dup_1622), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix16275 (.Y (nx16274), .A0 (rd_addr_m_1), .A1 (nx1755)
                          , .B0 (nx3378), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1756 (.Y (nx1755), .A (modgen_ram_ix167_a_232__dup_1629)
                      , .B (modgen_ram_ix167_a_233__dup_1628), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2785 (.Y (nx3378), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_1626), .B0 (nx16256), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix16257 (.Y (nx16256), .AN (
                      modgen_ram_ix167_a_234__dup_1627), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15671 (.Y (nx15670), .A0 (rd_addr_m_5), .A1 (nx3379)
                          , .B0 (nx3382), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2787 (.Y (nx3379), .A0 (rd_addr_m_4), .A1 (nx15214), .B0 (
                      nx14998)) ;
    MXT4_X0P5M_A12TS ix15215 (.Y (nx15214), .A (nx15046), .B (nx15154), .C (
                     nx15098), .D (nx15206), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix15047 (.Y (nx15046), .A (modgen_ram_ix167_a_144__dup_1717
                     ), .B (modgen_ram_ix167_a_146__dup_1715), .C (
                     modgen_ram_ix167_a_145__dup_1716), .D (
                     modgen_ram_ix167_a_147__dup_1714), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15155 (.Y (nx15154), .A (modgen_ram_ix167_a_152__dup_1709
                     ), .B (modgen_ram_ix167_a_154__dup_1707), .C (
                     modgen_ram_ix167_a_153__dup_1708), .D (
                     modgen_ram_ix167_a_155__dup_1706), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15099 (.Y (nx15098), .A (modgen_ram_ix167_a_148__dup_1713
                     ), .B (modgen_ram_ix167_a_150__dup_1711), .C (
                     modgen_ram_ix167_a_149__dup_1712), .D (
                     modgen_ram_ix167_a_151__dup_1710), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15207 (.Y (nx15206), .A (modgen_ram_ix167_a_156__dup_1705
                     ), .B (modgen_ram_ix167_a_158__dup_1703), .C (
                     modgen_ram_ix167_a_157__dup_1704), .D (
                     modgen_ram_ix167_a_159__dup_1702), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14999 (.Y (nx14998), .A0 (rd_addr_m_3), .A1 (nx3380)
                          , .B0 (nx1783), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2788 (.Y (nx3380), .A0 (rd_addr_m_2), .A1 (nx14878), .B0 (
                      nx14830)) ;
    MXT4_X0P5M_A12TS ix14879 (.Y (nx14878), .A (modgen_ram_ix167_a_132__dup_1729
                     ), .B (modgen_ram_ix167_a_134__dup_1727), .C (
                     modgen_ram_ix167_a_133__dup_1728), .D (
                     modgen_ram_ix167_a_135__dup_1726), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14831 (.Y (nx14830), .A0 (rd_addr_m_1), .A1 (nx1777)
                          , .B0 (nx1779), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1778 (.Y (nx1777), .A (modgen_ram_ix167_a_128__dup_1733)
                      , .B (modgen_ram_ix167_a_129__dup_1732), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1780 (.Y (nx1779), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_1730), .B0 (nx14812), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix14813 (.Y (nx14812), .AN (
                      modgen_ram_ix167_a_130__dup_1731), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1784 (.Y (nx1783), .A0 (rd_addr_m_2), .A1 (nx14986)
                          , .B0 (nx14938), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix14987 (.Y (nx14986), .A (modgen_ram_ix167_a_140__dup_1721
                     ), .B (modgen_ram_ix167_a_142__dup_1719), .C (
                     modgen_ram_ix167_a_141__dup_1720), .D (
                     modgen_ram_ix167_a_143__dup_1718), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14939 (.Y (nx14938), .A0 (rd_addr_m_1), .A1 (nx1789)
                          , .B0 (nx3381), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1790 (.Y (nx1789), .A (modgen_ram_ix167_a_136__dup_1725)
                      , .B (modgen_ram_ix167_a_137__dup_1724), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1792 (.Y (nx3381), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_1722), .B0 (nx14920), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix14921 (.Y (nx14920), .AN (
                      modgen_ram_ix167_a_138__dup_1723), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1795 (.Y (nx3382), .A0 (rd_addr_m_4), .A1 (nx15658)
                          , .B0 (nx15442), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix15659 (.Y (nx15658), .A (nx15490), .B (nx15598), .C (
                     nx15542), .D (nx15650), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix15491 (.Y (nx15490), .A (modgen_ram_ix167_a_176__dup_1685
                     ), .B (modgen_ram_ix167_a_178__dup_1683), .C (
                     modgen_ram_ix167_a_177__dup_1684), .D (
                     modgen_ram_ix167_a_179__dup_1682), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15599 (.Y (nx15598), .A (modgen_ram_ix167_a_184__dup_1677
                     ), .B (modgen_ram_ix167_a_186__dup_1675), .C (
                     modgen_ram_ix167_a_185__dup_1676), .D (
                     modgen_ram_ix167_a_187__dup_1674), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15543 (.Y (nx15542), .A (modgen_ram_ix167_a_180__dup_1681
                     ), .B (modgen_ram_ix167_a_182__dup_1679), .C (
                     modgen_ram_ix167_a_181__dup_1680), .D (
                     modgen_ram_ix167_a_183__dup_1678), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix15651 (.Y (nx15650), .A (modgen_ram_ix167_a_188__dup_1673
                     ), .B (modgen_ram_ix167_a_190__dup_1671), .C (
                     modgen_ram_ix167_a_189__dup_1672), .D (
                     modgen_ram_ix167_a_191__dup_1670), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15443 (.Y (nx15442), .A0 (rd_addr_m_3), .A1 (nx3383)
                          , .B0 (nx3386), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1808 (.Y (nx3383), .A0 (rd_addr_m_2), .A1 (nx15322), .B0 (
                      nx15274)) ;
    MXT4_X0P5M_A12TS ix15323 (.Y (nx15322), .A (modgen_ram_ix167_a_164__dup_1697
                     ), .B (modgen_ram_ix167_a_166__dup_1695), .C (
                     modgen_ram_ix167_a_165__dup_1696), .D (
                     modgen_ram_ix167_a_167__dup_1694), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15275 (.Y (nx15274), .A0 (rd_addr_m_1), .A1 (nx3384)
                          , .B0 (nx3385), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2789 (.Y (nx3384), .A (modgen_ram_ix167_a_160__dup_1701)
                      , .B (modgen_ram_ix167_a_161__dup_1700), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1814 (.Y (nx3385), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_1698), .B0 (nx15256), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix15257 (.Y (nx15256), .AN (
                      modgen_ram_ix167_a_162__dup_1699), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1818 (.Y (nx3386), .A0 (rd_addr_m_2), .A1 (nx15430)
                          , .B0 (nx15382), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix15431 (.Y (nx15430), .A (modgen_ram_ix167_a_172__dup_1689
                     ), .B (modgen_ram_ix167_a_174__dup_1687), .C (
                     modgen_ram_ix167_a_173__dup_1688), .D (
                     modgen_ram_ix167_a_175__dup_1686), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix15383 (.Y (nx15382), .A0 (rd_addr_m_1), .A1 (nx3387)
                          , .B0 (nx3388), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1822 (.Y (nx3387), .A (modgen_ram_ix167_a_168__dup_1693)
                      , .B (modgen_ram_ix167_a_169__dup_1692), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1824 (.Y (nx3388), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_1690), .B0 (nx15364), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix15365 (.Y (nx15364), .AN (
                      modgen_ram_ix167_a_170__dup_1691), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix14779 (.Y (nx14778), .A (rd_addr_7), .B (nx3389)) ;
    AOI21_X0P5M_A12TS ix1830 (.Y (nx3389), .A0 (rd_addr_m_6), .A1 (nx14770), .B0 (
                      nx13882)) ;
    OAI21_X0P5M_A12TS ix14771 (.Y (nx14770), .A0 (rd_addr_m_5), .A1 (nx3390), .B0 (
                      nx3397)) ;
    AOI21_X0P5M_A12TS ix1834 (.Y (nx3390), .A0 (rd_addr_m_4), .A1 (nx14318), .B0 (
                      nx14102)) ;
    MXT4_X0P5M_A12TS ix14319 (.Y (nx14318), .A (nx14150), .B (nx14258), .C (
                     nx14202), .D (nx14310), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix14151 (.Y (nx14150), .A (modgen_ram_ix167_a_80__dup_1781)
                     , .B (modgen_ram_ix167_a_82__dup_1779), .C (
                     modgen_ram_ix167_a_81__dup_1780), .D (
                     modgen_ram_ix167_a_83__dup_1778), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix14259 (.Y (nx14258), .A (modgen_ram_ix167_a_88__dup_1773)
                     , .B (modgen_ram_ix167_a_90__dup_1771), .C (
                     modgen_ram_ix167_a_89__dup_1772), .D (
                     modgen_ram_ix167_a_91__dup_1770), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix14203 (.Y (nx14202), .A (modgen_ram_ix167_a_84__dup_1777)
                     , .B (modgen_ram_ix167_a_86__dup_1775), .C (
                     modgen_ram_ix167_a_85__dup_1776), .D (
                     modgen_ram_ix167_a_87__dup_1774), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix14311 (.Y (nx14310), .A (modgen_ram_ix167_a_92__dup_1769)
                     , .B (modgen_ram_ix167_a_94__dup_1767), .C (
                     modgen_ram_ix167_a_93__dup_1768), .D (
                     modgen_ram_ix167_a_95__dup_1766), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14103 (.Y (nx14102), .A0 (rd_addr_m_3), .A1 (nx3391)
                          , .B0 (nx3394), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1842 (.Y (nx3391), .A0 (rd_addr_m_2), .A1 (nx13982), .B0 (
                      nx13934)) ;
    MXT4_X0P5M_A12TS ix13983 (.Y (nx13982), .A (modgen_ram_ix167_a_68__dup_1793)
                     , .B (modgen_ram_ix167_a_70__dup_1791), .C (
                     modgen_ram_ix167_a_69__dup_1792), .D (
                     modgen_ram_ix167_a_71__dup_1790), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13935 (.Y (nx13934), .A0 (rd_addr_m_1), .A1 (nx3392)
                          , .B0 (nx3393), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2790 (.Y (nx3392), .A (modgen_ram_ix167_a_64__dup_1797)
                      , .B (modgen_ram_ix167_a_65__dup_1796), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2791 (.Y (nx3393), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_1794), .B0 (nx13916), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix13917 (.Y (nx13916), .AN (
                      modgen_ram_ix167_a_66__dup_1795), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1854 (.Y (nx3394), .A0 (rd_addr_m_2), .A1 (nx14090)
                          , .B0 (nx14042), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix14091 (.Y (nx14090), .A (modgen_ram_ix167_a_76__dup_1785)
                     , .B (modgen_ram_ix167_a_78__dup_1783), .C (
                     modgen_ram_ix167_a_77__dup_1784), .D (
                     modgen_ram_ix167_a_79__dup_1782), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14043 (.Y (nx14042), .A0 (rd_addr_m_1), .A1 (nx3395)
                          , .B0 (nx3396), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1859 (.Y (nx3395), .A (modgen_ram_ix167_a_72__dup_1789)
                      , .B (modgen_ram_ix167_a_73__dup_1788), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2792 (.Y (nx3396), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_1786), .B0 (nx14024), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix14025 (.Y (nx14024), .AN (
                      modgen_ram_ix167_a_74__dup_1787), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1864 (.Y (nx3397), .A0 (rd_addr_m_4), .A1 (nx14762)
                          , .B0 (nx14546), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix14763 (.Y (nx14762), .A (nx14594), .B (nx14702), .C (
                     nx14646), .D (nx14754), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix14595 (.Y (nx14594), .A (modgen_ram_ix167_a_112__dup_1749
                     ), .B (modgen_ram_ix167_a_114__dup_1747), .C (
                     modgen_ram_ix167_a_113__dup_1748), .D (
                     modgen_ram_ix167_a_115__dup_1746), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix14703 (.Y (nx14702), .A (modgen_ram_ix167_a_120__dup_1741
                     ), .B (modgen_ram_ix167_a_122__dup_1739), .C (
                     modgen_ram_ix167_a_121__dup_1740), .D (
                     modgen_ram_ix167_a_123__dup_1738), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix14647 (.Y (nx14646), .A (modgen_ram_ix167_a_116__dup_1745
                     ), .B (modgen_ram_ix167_a_118__dup_1743), .C (
                     modgen_ram_ix167_a_117__dup_1744), .D (
                     modgen_ram_ix167_a_119__dup_1742), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix14755 (.Y (nx14754), .A (modgen_ram_ix167_a_124__dup_1737
                     ), .B (modgen_ram_ix167_a_126__dup_1735), .C (
                     modgen_ram_ix167_a_125__dup_1736), .D (
                     modgen_ram_ix167_a_127__dup_1734), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14547 (.Y (nx14546), .A0 (rd_addr_m_3), .A1 (nx3398)
                          , .B0 (nx3402), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2793 (.Y (nx3398), .A0 (rd_addr_m_2), .A1 (nx14426), .B0 (
                      nx14378)) ;
    MXT4_X0P5M_A12TS ix14427 (.Y (nx14426), .A (modgen_ram_ix167_a_100__dup_1761
                     ), .B (modgen_ram_ix167_a_102__dup_1759), .C (
                     modgen_ram_ix167_a_101__dup_1760), .D (
                     modgen_ram_ix167_a_103__dup_1758), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14379 (.Y (nx14378), .A0 (rd_addr_m_1), .A1 (nx3399)
                          , .B0 (nx3401), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2794 (.Y (nx3399), .A (modgen_ram_ix167_a_96__dup_1765)
                      , .B (modgen_ram_ix167_a_97__dup_1764), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1880 (.Y (nx3401), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_1762), .B0 (nx14360), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix14361 (.Y (nx14360), .AN (
                      modgen_ram_ix167_a_98__dup_1763), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1884 (.Y (nx3402), .A0 (rd_addr_m_2), .A1 (nx14534)
                          , .B0 (nx14486), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix14535 (.Y (nx14534), .A (modgen_ram_ix167_a_108__dup_1753
                     ), .B (modgen_ram_ix167_a_110__dup_1751), .C (
                     modgen_ram_ix167_a_109__dup_1752), .D (
                     modgen_ram_ix167_a_111__dup_1750), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix14487 (.Y (nx14486), .A0 (rd_addr_m_1), .A1 (nx3403)
                          , .B0 (nx3404), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1890 (.Y (nx3403), .A (modgen_ram_ix167_a_104__dup_1757)
                      , .B (modgen_ram_ix167_a_105__dup_1756), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix1892 (.Y (nx3404), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_1754), .B0 (nx14468), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix14469 (.Y (nx14468), .AN (
                      modgen_ram_ix167_a_106__dup_1755), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13883 (.Y (nx13882), .A0 (rd_addr_m_5), .A1 (nx3405)
                          , .B0 (nx1929), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix1898 (.Y (nx3405), .A0 (rd_addr_m_4), .A1 (nx13426), .B0 (
                      nx13210)) ;
    MXT4_X0P5M_A12TS ix13427 (.Y (nx13426), .A (nx13258), .B (nx13366), .C (
                     nx13310), .D (nx13418), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix13259 (.Y (nx13258), .A (modgen_ram_ix167_a_16__dup_1845)
                     , .B (modgen_ram_ix167_a_18__dup_1843), .C (
                     modgen_ram_ix167_a_17__dup_1844), .D (
                     modgen_ram_ix167_a_19__dup_1842), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix13367 (.Y (nx13366), .A (modgen_ram_ix167_a_24__dup_1837)
                     , .B (modgen_ram_ix167_a_26__dup_1835), .C (
                     modgen_ram_ix167_a_25__dup_1836), .D (
                     modgen_ram_ix167_a_27__dup_1834), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix13311 (.Y (nx13310), .A (modgen_ram_ix167_a_20__dup_1841)
                     , .B (modgen_ram_ix167_a_22__dup_1839), .C (
                     modgen_ram_ix167_a_21__dup_1840), .D (
                     modgen_ram_ix167_a_23__dup_1838), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix13419 (.Y (nx13418), .A (modgen_ram_ix167_a_28__dup_1833)
                     , .B (modgen_ram_ix167_a_30__dup_1831), .C (
                     modgen_ram_ix167_a_29__dup_1832), .D (
                     modgen_ram_ix167_a_31__dup_1830), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13211 (.Y (nx13210), .A0 (rd_addr_m_3), .A1 (nx3406)
                          , .B0 (nx3409), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix1910 (.Y (nx3406), .A0 (rd_addr_m_2), .A1 (nx13090), .B0 (
                      nx13042)) ;
    MXT4_X0P5M_A12TS ix13091 (.Y (nx13090), .A (modgen_ram_ix167_a_4__dup_1857)
                     , .B (modgen_ram_ix167_a_6__dup_1855), .C (
                     modgen_ram_ix167_a_5__dup_1856), .D (
                     modgen_ram_ix167_a_7__dup_1854), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13043 (.Y (nx13042), .A0 (rd_addr_m_1), .A1 (nx3407)
                          , .B0 (nx3408), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1914 (.Y (nx3407), .A (modgen_ram_ix167_a_0__dup_1861), 
                      .B (modgen_ram_ix167_a_1__dup_1860), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1916 (.Y (nx3408), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_1858), .B0 (nx13024), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix13025 (.Y (nx13024), .AN (modgen_ram_ix167_a_2__dup_1859
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1920 (.Y (nx3409), .A0 (rd_addr_m_2), .A1 (nx13198)
                          , .B0 (nx13150), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix13199 (.Y (nx13198), .A (modgen_ram_ix167_a_12__dup_1849)
                     , .B (modgen_ram_ix167_a_14__dup_1847), .C (
                     modgen_ram_ix167_a_13__dup_1848), .D (
                     modgen_ram_ix167_a_15__dup_1846), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13151 (.Y (nx13150), .A0 (rd_addr_m_1), .A1 (nx3411)
                          , .B0 (nx3412), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix1924 (.Y (nx3411), .A (modgen_ram_ix167_a_8__dup_1853), 
                      .B (modgen_ram_ix167_a_9__dup_1852), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix1926 (.Y (nx3412), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_1850), .B0 (nx13132), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix13133 (.Y (nx13132), .AN (
                      modgen_ram_ix167_a_10__dup_1851), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2795 (.Y (nx1929), .A0 (rd_addr_m_4), .A1 (nx13870)
                          , .B0 (nx13654), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix13871 (.Y (nx13870), .A (nx13702), .B (nx13810), .C (
                     nx13754), .D (nx13862), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix13703 (.Y (nx13702), .A (modgen_ram_ix167_a_48__dup_1813)
                     , .B (modgen_ram_ix167_a_50__dup_1811), .C (
                     modgen_ram_ix167_a_49__dup_1812), .D (
                     modgen_ram_ix167_a_51__dup_1810), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix13811 (.Y (nx13810), .A (modgen_ram_ix167_a_56__dup_1805)
                     , .B (modgen_ram_ix167_a_58__dup_1803), .C (
                     modgen_ram_ix167_a_57__dup_1804), .D (
                     modgen_ram_ix167_a_59__dup_1802), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix13755 (.Y (nx13754), .A (modgen_ram_ix167_a_52__dup_1809)
                     , .B (modgen_ram_ix167_a_54__dup_1807), .C (
                     modgen_ram_ix167_a_53__dup_1808), .D (
                     modgen_ram_ix167_a_55__dup_1806), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix13863 (.Y (nx13862), .A (modgen_ram_ix167_a_60__dup_1801)
                     , .B (modgen_ram_ix167_a_62__dup_1799), .C (
                     modgen_ram_ix167_a_61__dup_1800), .D (
                     modgen_ram_ix167_a_63__dup_1798), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13655 (.Y (nx13654), .A0 (rd_addr_m_3), .A1 (nx1939)
                          , .B0 (nx1951), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2796 (.Y (nx1939), .A0 (rd_addr_m_2), .A1 (nx13534), .B0 (
                      nx13486)) ;
    MXT4_X0P5M_A12TS ix13535 (.Y (nx13534), .A (modgen_ram_ix167_a_36__dup_1825)
                     , .B (modgen_ram_ix167_a_38__dup_1823), .C (
                     modgen_ram_ix167_a_37__dup_1824), .D (
                     modgen_ram_ix167_a_39__dup_1822), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13487 (.Y (nx13486), .A0 (rd_addr_m_1), .A1 (nx3413)
                          , .B0 (nx3414), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2797 (.Y (nx3413), .A (modgen_ram_ix167_a_32__dup_1829)
                      , .B (modgen_ram_ix167_a_33__dup_1828), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2798 (.Y (nx3414), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_1826), .B0 (nx13468), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix13469 (.Y (nx13468), .AN (
                      modgen_ram_ix167_a_34__dup_1827), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2799 (.Y (nx1951), .A0 (rd_addr_m_2), .A1 (nx13642)
                          , .B0 (nx13594), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix13643 (.Y (nx13642), .A (modgen_ram_ix167_a_44__dup_1817)
                     , .B (modgen_ram_ix167_a_46__dup_1815), .C (
                     modgen_ram_ix167_a_45__dup_1816), .D (
                     modgen_ram_ix167_a_47__dup_1814), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix13595 (.Y (nx13594), .A0 (rd_addr_m_1), .A1 (nx1955)
                          , .B0 (nx1957), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2800 (.Y (nx1955), .A (modgen_ram_ix167_a_40__dup_1821)
                      , .B (modgen_ram_ix167_a_41__dup_1820), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2801 (.Y (nx1957), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_1818), .B0 (nx13576), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix13577 (.Y (nx13576), .AN (
                      modgen_ram_ix167_a_42__dup_1819), .B (rd_addr_m_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_4 (.Q (rd_data_m_4), .CK (wb_clk_i), .D (
                        nx20162), .R (wb_rst_i), .SE (NOT_nx50), .SI (
                        rd_data_m_4)) ;
    MXIT2_X0P5M_A12TS ix20163 (.Y (nx20162), .A (nx3415), .B (nx1965), .S0 (
                      nx1127)) ;
    INV_X0P5B_A12TS ix2802 (.Y (nx3415), .A (wr_data_m_4)) ;
    OA21A1OI2_X0P5M_A12TS ix2803 (.Y (nx1965), .A0 (nx20148), .A1 (nx19258), .B0 (
                          rd_addr_7), .C0 (nx18366)) ;
    OA21A1OI2_X0P5M_A12TS ix20149 (.Y (nx20148), .A0 (rd_addr_m_5), .A1 (nx1969)
                          , .B0 (nx3417), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2804 (.Y (nx1969), .A0 (rd_addr_m_4), .A1 (nx19694), .B0 (
                      nx19478)) ;
    MXT4_X0P5M_A12TS ix19695 (.Y (nx19694), .A (nx19526), .B (nx19634), .C (
                     nx19578), .D (nx19686), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix19527 (.Y (nx19526), .A (modgen_ram_ix167_a_208__dup_1389
                     ), .B (modgen_ram_ix167_a_210__dup_1387), .C (
                     modgen_ram_ix167_a_209__dup_1388), .D (
                     modgen_ram_ix167_a_211__dup_1386), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix19635 (.Y (nx19634), .A (modgen_ram_ix167_a_216__dup_1381
                     ), .B (modgen_ram_ix167_a_218__dup_1379), .C (
                     modgen_ram_ix167_a_217__dup_1380), .D (
                     modgen_ram_ix167_a_219__dup_1378), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix19579 (.Y (nx19578), .A (modgen_ram_ix167_a_212__dup_1385
                     ), .B (modgen_ram_ix167_a_214__dup_1383), .C (
                     modgen_ram_ix167_a_213__dup_1384), .D (
                     modgen_ram_ix167_a_215__dup_1382), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix19687 (.Y (nx19686), .A (modgen_ram_ix167_a_220__dup_1377
                     ), .B (modgen_ram_ix167_a_222__dup_1375), .C (
                     modgen_ram_ix167_a_221__dup_1376), .D (
                     modgen_ram_ix167_a_223__dup_1374), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19479 (.Y (nx19478), .A0 (rd_addr_m_3), .A1 (nx1979)
                          , .B0 (nx3416), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2805 (.Y (nx1979), .A0 (rd_addr_m_2), .A1 (nx19358), .B0 (
                      nx19310)) ;
    MXT4_X0P5M_A12TS ix19359 (.Y (nx19358), .A (modgen_ram_ix167_a_196__dup_1401
                     ), .B (modgen_ram_ix167_a_198__dup_1399), .C (
                     modgen_ram_ix167_a_197__dup_1400), .D (
                     modgen_ram_ix167_a_199__dup_1398), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19311 (.Y (nx19310), .A0 (rd_addr_m_1), .A1 (nx1985)
                          , .B0 (nx1987), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2806 (.Y (nx1985), .A (modgen_ram_ix167_a_192__dup_1405)
                      , .B (modgen_ram_ix167_a_193__dup_1404), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2807 (.Y (nx1987), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_1402), .B0 (nx19292), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix19293 (.Y (nx19292), .AN (
                      modgen_ram_ix167_a_194__dup_1403), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2808 (.Y (nx3416), .A0 (rd_addr_m_2), .A1 (nx19466)
                          , .B0 (nx19418), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix19467 (.Y (nx19466), .A (modgen_ram_ix167_a_204__dup_1393
                     ), .B (modgen_ram_ix167_a_206__dup_1391), .C (
                     modgen_ram_ix167_a_205__dup_1392), .D (
                     modgen_ram_ix167_a_207__dup_1390), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19419 (.Y (nx19418), .A0 (rd_addr_m_1), .A1 (nx1996)
                          , .B0 (nx1998), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2809 (.Y (nx1996), .A (modgen_ram_ix167_a_200__dup_1397)
                      , .B (modgen_ram_ix167_a_201__dup_1396), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2810 (.Y (nx1998), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_1394), .B0 (nx19400), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix19401 (.Y (nx19400), .AN (
                      modgen_ram_ix167_a_202__dup_1395), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2811 (.Y (nx3417), .A0 (rd_addr_m_4), .A1 (nx20138)
                          , .B0 (nx19922), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix20139 (.Y (nx20138), .A (nx19970), .B (nx20078), .C (
                     nx20022), .D (nx20130), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix19971 (.Y (nx19970), .A (modgen_ram_ix167_a_240__dup_1357
                     ), .B (modgen_ram_ix167_a_242__dup_1355), .C (
                     modgen_ram_ix167_a_241__dup_1356), .D (
                     modgen_ram_ix167_a_243__dup_1354), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20079 (.Y (nx20078), .A (modgen_ram_ix167_a_248__dup_1349
                     ), .B (modgen_ram_ix167_a_250__dup_1347), .C (
                     modgen_ram_ix167_a_249__dup_1348), .D (
                     modgen_ram_ix167_a_251__dup_1346), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20023 (.Y (nx20022), .A (modgen_ram_ix167_a_244__dup_1353
                     ), .B (modgen_ram_ix167_a_246__dup_1351), .C (
                     modgen_ram_ix167_a_245__dup_1352), .D (
                     modgen_ram_ix167_a_247__dup_1350), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20131 (.Y (nx20130), .A (modgen_ram_ix167_a_252__dup_1345
                     ), .B (modgen_ram_ix167_a_254__dup_1343), .C (
                     modgen_ram_ix167_a_253__dup_1344), .D (
                     modgen_ram_ix167_a_255__dup_1342), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19923 (.Y (nx19922), .A0 (rd_addr_m_3), .A1 (nx2011)
                          , .B0 (nx3420), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2812 (.Y (nx2011), .A0 (rd_addr_m_2), .A1 (nx19802), .B0 (
                      nx19754)) ;
    MXT4_X0P5M_A12TS ix19803 (.Y (nx19802), .A (modgen_ram_ix167_a_228__dup_1369
                     ), .B (modgen_ram_ix167_a_230__dup_1367), .C (
                     modgen_ram_ix167_a_229__dup_1368), .D (
                     modgen_ram_ix167_a_231__dup_1366), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19755 (.Y (nx19754), .A0 (rd_addr_m_1), .A1 (nx3418)
                          , .B0 (nx3419), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2813 (.Y (nx3418), .A (modgen_ram_ix167_a_224__dup_1373)
                      , .B (modgen_ram_ix167_a_225__dup_1372), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2814 (.Y (nx3419), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_1370), .B0 (nx19736), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix19737 (.Y (nx19736), .AN (
                      modgen_ram_ix167_a_226__dup_1371), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2815 (.Y (nx3420), .A0 (rd_addr_m_2), .A1 (nx19910)
                          , .B0 (nx19862), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix19911 (.Y (nx19910), .A (modgen_ram_ix167_a_236__dup_1361
                     ), .B (modgen_ram_ix167_a_238__dup_1359), .C (
                     modgen_ram_ix167_a_237__dup_1360), .D (
                     modgen_ram_ix167_a_239__dup_1358), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19863 (.Y (nx19862), .A0 (rd_addr_m_1), .A1 (nx2025)
                          , .B0 (nx2027), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2816 (.Y (nx2025), .A (modgen_ram_ix167_a_232__dup_1365)
                      , .B (modgen_ram_ix167_a_233__dup_1364), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2817 (.Y (nx2027), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_1362), .B0 (nx19844), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix19845 (.Y (nx19844), .AN (
                      modgen_ram_ix167_a_234__dup_1363), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19259 (.Y (nx19258), .A0 (rd_addr_m_5), .A1 (nx3421)
                          , .B0 (nx3423), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2818 (.Y (nx3421), .A0 (rd_addr_m_4), .A1 (nx18802), .B0 (
                      nx18586)) ;
    MXT4_X0P5M_A12TS ix18803 (.Y (nx18802), .A (nx18634), .B (nx18742), .C (
                     nx18686), .D (nx18794), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix18635 (.Y (nx18634), .A (modgen_ram_ix167_a_144__dup_1453
                     ), .B (modgen_ram_ix167_a_146__dup_1451), .C (
                     modgen_ram_ix167_a_145__dup_1452), .D (
                     modgen_ram_ix167_a_147__dup_1450), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix18743 (.Y (nx18742), .A (modgen_ram_ix167_a_152__dup_1445
                     ), .B (modgen_ram_ix167_a_154__dup_1443), .C (
                     modgen_ram_ix167_a_153__dup_1444), .D (
                     modgen_ram_ix167_a_155__dup_1442), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix18687 (.Y (nx18686), .A (modgen_ram_ix167_a_148__dup_1449
                     ), .B (modgen_ram_ix167_a_150__dup_1447), .C (
                     modgen_ram_ix167_a_149__dup_1448), .D (
                     modgen_ram_ix167_a_151__dup_1446), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix18795 (.Y (nx18794), .A (modgen_ram_ix167_a_156__dup_1441
                     ), .B (modgen_ram_ix167_a_158__dup_1439), .C (
                     modgen_ram_ix167_a_157__dup_1440), .D (
                     modgen_ram_ix167_a_159__dup_1438), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18587 (.Y (nx18586), .A0 (rd_addr_m_3), .A1 (nx2041)
                          , .B0 (nx2053), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2820 (.Y (nx2041), .A0 (rd_addr_m_2), .A1 (nx18466), .B0 (
                      nx18418)) ;
    MXT4_X0P5M_A12TS ix18467 (.Y (nx18466), .A (modgen_ram_ix167_a_132__dup_1465
                     ), .B (modgen_ram_ix167_a_134__dup_1463), .C (
                     modgen_ram_ix167_a_133__dup_1464), .D (
                     modgen_ram_ix167_a_135__dup_1462), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18419 (.Y (nx18418), .A0 (rd_addr_m_1), .A1 (nx2047)
                          , .B0 (nx2049), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2821 (.Y (nx2047), .A (modgen_ram_ix167_a_128__dup_1469)
                      , .B (modgen_ram_ix167_a_129__dup_1468), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2050 (.Y (nx2049), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_1466), .B0 (nx18400), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix18401 (.Y (nx18400), .AN (
                      modgen_ram_ix167_a_130__dup_1467), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2054 (.Y (nx2053), .A0 (rd_addr_m_2), .A1 (nx18574)
                          , .B0 (nx18526), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix18575 (.Y (nx18574), .A (modgen_ram_ix167_a_140__dup_1457
                     ), .B (modgen_ram_ix167_a_142__dup_1455), .C (
                     modgen_ram_ix167_a_141__dup_1456), .D (
                     modgen_ram_ix167_a_143__dup_1454), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18527 (.Y (nx18526), .A0 (rd_addr_m_1), .A1 (nx2057)
                          , .B0 (nx3422), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2058 (.Y (nx2057), .A (modgen_ram_ix167_a_136__dup_1461)
                      , .B (modgen_ram_ix167_a_137__dup_1460), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2822 (.Y (nx3422), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_1458), .B0 (nx18508), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix18509 (.Y (nx18508), .AN (
                      modgen_ram_ix167_a_138__dup_1459), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2823 (.Y (nx3423), .A0 (rd_addr_m_4), .A1 (nx19246)
                          , .B0 (nx19030), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix19247 (.Y (nx19246), .A (nx19078), .B (nx19186), .C (
                     nx19130), .D (nx19238), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix19079 (.Y (nx19078), .A (modgen_ram_ix167_a_176__dup_1421
                     ), .B (modgen_ram_ix167_a_178__dup_1419), .C (
                     modgen_ram_ix167_a_177__dup_1420), .D (
                     modgen_ram_ix167_a_179__dup_1418), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix19187 (.Y (nx19186), .A (modgen_ram_ix167_a_184__dup_1413
                     ), .B (modgen_ram_ix167_a_186__dup_1411), .C (
                     modgen_ram_ix167_a_185__dup_1412), .D (
                     modgen_ram_ix167_a_187__dup_1410), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix19131 (.Y (nx19130), .A (modgen_ram_ix167_a_180__dup_1417
                     ), .B (modgen_ram_ix167_a_182__dup_1415), .C (
                     modgen_ram_ix167_a_181__dup_1416), .D (
                     modgen_ram_ix167_a_183__dup_1414), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix19239 (.Y (nx19238), .A (modgen_ram_ix167_a_188__dup_1409
                     ), .B (modgen_ram_ix167_a_190__dup_1407), .C (
                     modgen_ram_ix167_a_189__dup_1408), .D (
                     modgen_ram_ix167_a_191__dup_1406), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix19031 (.Y (nx19030), .A0 (rd_addr_m_3), .A1 (nx2075)
                          , .B0 (nx3427), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2076 (.Y (nx2075), .A0 (rd_addr_m_2), .A1 (nx18910), .B0 (
                      nx18862)) ;
    MXT4_X0P5M_A12TS ix18911 (.Y (nx18910), .A (modgen_ram_ix167_a_164__dup_1433
                     ), .B (modgen_ram_ix167_a_166__dup_1431), .C (
                     modgen_ram_ix167_a_165__dup_1432), .D (
                     modgen_ram_ix167_a_167__dup_1430), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18863 (.Y (nx18862), .A0 (rd_addr_m_1), .A1 (nx3424)
                          , .B0 (nx3425), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2824 (.Y (nx3424), .A (modgen_ram_ix167_a_160__dup_1437)
                      , .B (modgen_ram_ix167_a_161__dup_1436), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2825 (.Y (nx3425), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_1434), .B0 (nx18844), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix18845 (.Y (nx18844), .AN (
                      modgen_ram_ix167_a_162__dup_1435), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2826 (.Y (nx3427), .A0 (rd_addr_m_2), .A1 (nx19018)
                          , .B0 (nx18970), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix19019 (.Y (nx19018), .A (modgen_ram_ix167_a_172__dup_1425
                     ), .B (modgen_ram_ix167_a_174__dup_1423), .C (
                     modgen_ram_ix167_a_173__dup_1424), .D (
                     modgen_ram_ix167_a_175__dup_1422), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18971 (.Y (nx18970), .A0 (rd_addr_m_1), .A1 (nx3428)
                          , .B0 (nx3429), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2092 (.Y (nx3428), .A (modgen_ram_ix167_a_168__dup_1429)
                      , .B (modgen_ram_ix167_a_169__dup_1428), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2094 (.Y (nx3429), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_1426), .B0 (nx18952), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix18953 (.Y (nx18952), .AN (
                      modgen_ram_ix167_a_170__dup_1427), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix18367 (.Y (nx18366), .A (rd_addr_7), .B (nx3430)) ;
    AOI21_X0P5M_A12TS ix2828 (.Y (nx3430), .A0 (rd_addr_m_6), .A1 (nx18358), .B0 (
                      nx17470)) ;
    OAI21_X0P5M_A12TS ix18359 (.Y (nx18358), .A0 (rd_addr_m_5), .A1 (nx3431), .B0 (
                      nx3440)) ;
    AOI21_X0P5M_A12TS ix2103 (.Y (nx3431), .A0 (rd_addr_m_4), .A1 (nx17906), .B0 (
                      nx17690)) ;
    MXT4_X0P5M_A12TS ix17907 (.Y (nx17906), .A (nx17738), .B (nx17846), .C (
                     nx17790), .D (nx17898), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix17739 (.Y (nx17738), .A (modgen_ram_ix167_a_80__dup_1517)
                     , .B (modgen_ram_ix167_a_82__dup_1515), .C (
                     modgen_ram_ix167_a_81__dup_1516), .D (
                     modgen_ram_ix167_a_83__dup_1514), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17847 (.Y (nx17846), .A (modgen_ram_ix167_a_88__dup_1509)
                     , .B (modgen_ram_ix167_a_90__dup_1507), .C (
                     modgen_ram_ix167_a_89__dup_1508), .D (
                     modgen_ram_ix167_a_91__dup_1506), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17791 (.Y (nx17790), .A (modgen_ram_ix167_a_84__dup_1513)
                     , .B (modgen_ram_ix167_a_86__dup_1511), .C (
                     modgen_ram_ix167_a_85__dup_1512), .D (
                     modgen_ram_ix167_a_87__dup_1510), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17899 (.Y (nx17898), .A (modgen_ram_ix167_a_92__dup_1505)
                     , .B (modgen_ram_ix167_a_94__dup_1503), .C (
                     modgen_ram_ix167_a_93__dup_1504), .D (
                     modgen_ram_ix167_a_95__dup_1502), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17691 (.Y (nx17690), .A0 (rd_addr_m_3), .A1 (nx3433)
                          , .B0 (nx3436), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2114 (.Y (nx3433), .A0 (rd_addr_m_2), .A1 (nx17570), .B0 (
                      nx17522)) ;
    MXT4_X0P5M_A12TS ix17571 (.Y (nx17570), .A (modgen_ram_ix167_a_68__dup_1529)
                     , .B (modgen_ram_ix167_a_70__dup_1527), .C (
                     modgen_ram_ix167_a_69__dup_1528), .D (
                     modgen_ram_ix167_a_71__dup_1526), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17523 (.Y (nx17522), .A0 (rd_addr_m_1), .A1 (nx3434)
                          , .B0 (nx3435), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2829 (.Y (nx3434), .A (modgen_ram_ix167_a_64__dup_1533)
                      , .B (modgen_ram_ix167_a_65__dup_1532), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2830 (.Y (nx3435), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_1530), .B0 (nx17504), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix17505 (.Y (nx17504), .AN (
                      modgen_ram_ix167_a_66__dup_1531), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2831 (.Y (nx3436), .A0 (rd_addr_m_2), .A1 (nx17678)
                          , .B0 (nx17630), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix17679 (.Y (nx17678), .A (modgen_ram_ix167_a_76__dup_1521)
                     , .B (modgen_ram_ix167_a_78__dup_1519), .C (
                     modgen_ram_ix167_a_77__dup_1520), .D (
                     modgen_ram_ix167_a_79__dup_1518), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17631 (.Y (nx17630), .A0 (rd_addr_m_1), .A1 (nx3437)
                          , .B0 (nx3439), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2128 (.Y (nx3437), .A (modgen_ram_ix167_a_72__dup_1525)
                      , .B (modgen_ram_ix167_a_73__dup_1524), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2130 (.Y (nx3439), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_1522), .B0 (nx17612), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix17613 (.Y (nx17612), .AN (
                      modgen_ram_ix167_a_74__dup_1523), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2832 (.Y (nx3440), .A0 (rd_addr_m_4), .A1 (nx18350)
                          , .B0 (nx18134), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix18351 (.Y (nx18350), .A (nx18182), .B (nx18290), .C (
                     nx18234), .D (nx18342), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix18183 (.Y (nx18182), .A (modgen_ram_ix167_a_112__dup_1485
                     ), .B (modgen_ram_ix167_a_114__dup_1483), .C (
                     modgen_ram_ix167_a_113__dup_1484), .D (
                     modgen_ram_ix167_a_115__dup_1482), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix18291 (.Y (nx18290), .A (modgen_ram_ix167_a_120__dup_1477
                     ), .B (modgen_ram_ix167_a_122__dup_1475), .C (
                     modgen_ram_ix167_a_121__dup_1476), .D (
                     modgen_ram_ix167_a_123__dup_1474), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix18235 (.Y (nx18234), .A (modgen_ram_ix167_a_116__dup_1481
                     ), .B (modgen_ram_ix167_a_118__dup_1479), .C (
                     modgen_ram_ix167_a_117__dup_1480), .D (
                     modgen_ram_ix167_a_119__dup_1478), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix18343 (.Y (nx18342), .A (modgen_ram_ix167_a_124__dup_1473
                     ), .B (modgen_ram_ix167_a_126__dup_1471), .C (
                     modgen_ram_ix167_a_125__dup_1472), .D (
                     modgen_ram_ix167_a_127__dup_1470), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18135 (.Y (nx18134), .A0 (rd_addr_m_3), .A1 (nx3441)
                          , .B0 (nx3444), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2144 (.Y (nx3441), .A0 (rd_addr_m_2), .A1 (nx18014), .B0 (
                      nx17966)) ;
    MXT4_X0P5M_A12TS ix18015 (.Y (nx18014), .A (modgen_ram_ix167_a_100__dup_1497
                     ), .B (modgen_ram_ix167_a_102__dup_1495), .C (
                     modgen_ram_ix167_a_101__dup_1496), .D (
                     modgen_ram_ix167_a_103__dup_1494), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17967 (.Y (nx17966), .A0 (rd_addr_m_1), .A1 (nx3442)
                          , .B0 (nx3443), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2148 (.Y (nx3442), .A (modgen_ram_ix167_a_96__dup_1501)
                      , .B (modgen_ram_ix167_a_97__dup_1500), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2150 (.Y (nx3443), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_1498), .B0 (nx17948), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix17949 (.Y (nx17948), .AN (
                      modgen_ram_ix167_a_98__dup_1499), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2154 (.Y (nx3444), .A0 (rd_addr_m_2), .A1 (nx18122)
                          , .B0 (nx18074), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix18123 (.Y (nx18122), .A (modgen_ram_ix167_a_108__dup_1489
                     ), .B (modgen_ram_ix167_a_110__dup_1487), .C (
                     modgen_ram_ix167_a_109__dup_1488), .D (
                     modgen_ram_ix167_a_111__dup_1486), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix18075 (.Y (nx18074), .A0 (rd_addr_m_1), .A1 (nx3445)
                          , .B0 (nx3446), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2833 (.Y (nx3445), .A (modgen_ram_ix167_a_104__dup_1493)
                      , .B (modgen_ram_ix167_a_105__dup_1492), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2160 (.Y (nx3446), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_1490), .B0 (nx18056), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix18057 (.Y (nx18056), .AN (
                      modgen_ram_ix167_a_106__dup_1491), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17471 (.Y (nx17470), .A0 (rd_addr_m_5), .A1 (nx3447)
                          , .B0 (nx3452), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2166 (.Y (nx3447), .A0 (rd_addr_m_4), .A1 (nx17014), .B0 (
                      nx16798)) ;
    MXT4_X0P5M_A12TS ix17015 (.Y (nx17014), .A (nx16846), .B (nx16954), .C (
                     nx16898), .D (nx17006), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix16847 (.Y (nx16846), .A (modgen_ram_ix167_a_16__dup_1581)
                     , .B (modgen_ram_ix167_a_18__dup_1579), .C (
                     modgen_ram_ix167_a_17__dup_1580), .D (
                     modgen_ram_ix167_a_19__dup_1578), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16955 (.Y (nx16954), .A (modgen_ram_ix167_a_24__dup_1573)
                     , .B (modgen_ram_ix167_a_26__dup_1571), .C (
                     modgen_ram_ix167_a_25__dup_1572), .D (
                     modgen_ram_ix167_a_27__dup_1570), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix16899 (.Y (nx16898), .A (modgen_ram_ix167_a_20__dup_1577)
                     , .B (modgen_ram_ix167_a_22__dup_1575), .C (
                     modgen_ram_ix167_a_21__dup_1576), .D (
                     modgen_ram_ix167_a_23__dup_1574), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17007 (.Y (nx17006), .A (modgen_ram_ix167_a_28__dup_1569)
                     , .B (modgen_ram_ix167_a_30__dup_1567), .C (
                     modgen_ram_ix167_a_29__dup_1568), .D (
                     modgen_ram_ix167_a_31__dup_1566), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix16799 (.Y (nx16798), .A0 (rd_addr_m_3), .A1 (nx3448)
                          , .B0 (nx2185), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2834 (.Y (nx3448), .A0 (rd_addr_m_2), .A1 (nx16678), .B0 (
                      nx16630)) ;
    MXT4_X0P5M_A12TS ix16679 (.Y (nx16678), .A (modgen_ram_ix167_a_4__dup_1593)
                     , .B (modgen_ram_ix167_a_6__dup_1591), .C (
                     modgen_ram_ix167_a_5__dup_1592), .D (
                     modgen_ram_ix167_a_7__dup_1590), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix16631 (.Y (nx16630), .A0 (rd_addr_m_1), .A1 (nx3449)
                          , .B0 (nx2181), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2835 (.Y (nx3449), .A (modgen_ram_ix167_a_0__dup_1597), 
                      .B (modgen_ram_ix167_a_1__dup_1596), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2836 (.Y (nx2181), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_1594), .B0 (nx16612), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix16613 (.Y (nx16612), .AN (modgen_ram_ix167_a_2__dup_1595
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2837 (.Y (nx2185), .A0 (rd_addr_m_2), .A1 (nx16786)
                          , .B0 (nx16738), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix16787 (.Y (nx16786), .A (modgen_ram_ix167_a_12__dup_1585)
                     , .B (modgen_ram_ix167_a_14__dup_1583), .C (
                     modgen_ram_ix167_a_13__dup_1584), .D (
                     modgen_ram_ix167_a_15__dup_1582), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix16739 (.Y (nx16738), .A0 (rd_addr_m_1), .A1 (nx3451)
                          , .B0 (nx2191), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2838 (.Y (nx3451), .A (modgen_ram_ix167_a_8__dup_1589), 
                      .B (modgen_ram_ix167_a_9__dup_1588), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2840 (.Y (nx2191), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_1586), .B0 (nx16720), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix16721 (.Y (nx16720), .AN (
                      modgen_ram_ix167_a_10__dup_1587), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2841 (.Y (nx3452), .A0 (rd_addr_m_4), .A1 (nx17458)
                          , .B0 (nx17242), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix17459 (.Y (nx17458), .A (nx17290), .B (nx17398), .C (
                     nx17342), .D (nx17450), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix17291 (.Y (nx17290), .A (modgen_ram_ix167_a_48__dup_1549)
                     , .B (modgen_ram_ix167_a_50__dup_1547), .C (
                     modgen_ram_ix167_a_49__dup_1548), .D (
                     modgen_ram_ix167_a_51__dup_1546), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17399 (.Y (nx17398), .A (modgen_ram_ix167_a_56__dup_1541)
                     , .B (modgen_ram_ix167_a_58__dup_1539), .C (
                     modgen_ram_ix167_a_57__dup_1540), .D (
                     modgen_ram_ix167_a_59__dup_1538), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17343 (.Y (nx17342), .A (modgen_ram_ix167_a_52__dup_1545)
                     , .B (modgen_ram_ix167_a_54__dup_1543), .C (
                     modgen_ram_ix167_a_53__dup_1544), .D (
                     modgen_ram_ix167_a_55__dup_1542), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix17451 (.Y (nx17450), .A (modgen_ram_ix167_a_60__dup_1537)
                     , .B (modgen_ram_ix167_a_62__dup_1535), .C (
                     modgen_ram_ix167_a_61__dup_1536), .D (
                     modgen_ram_ix167_a_63__dup_1534), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17243 (.Y (nx17242), .A0 (rd_addr_m_3), .A1 (nx2205)
                          , .B0 (nx2215), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2842 (.Y (nx2205), .A0 (rd_addr_m_2), .A1 (nx17122), .B0 (
                      nx17074)) ;
    MXT4_X0P5M_A12TS ix17123 (.Y (nx17122), .A (modgen_ram_ix167_a_36__dup_1561)
                     , .B (modgen_ram_ix167_a_38__dup_1559), .C (
                     modgen_ram_ix167_a_37__dup_1560), .D (
                     modgen_ram_ix167_a_39__dup_1558), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17075 (.Y (nx17074), .A0 (rd_addr_m_1), .A1 (nx3453)
                          , .B0 (nx2211), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2843 (.Y (nx3453), .A (modgen_ram_ix167_a_32__dup_1565)
                      , .B (modgen_ram_ix167_a_33__dup_1564), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2844 (.Y (nx2211), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_1562), .B0 (nx17056), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix17057 (.Y (nx17056), .AN (
                      modgen_ram_ix167_a_34__dup_1563), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2845 (.Y (nx2215), .A0 (rd_addr_m_2), .A1 (nx17230)
                          , .B0 (nx17182), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix17231 (.Y (nx17230), .A (modgen_ram_ix167_a_44__dup_1553)
                     , .B (modgen_ram_ix167_a_46__dup_1551), .C (
                     modgen_ram_ix167_a_45__dup_1552), .D (
                     modgen_ram_ix167_a_47__dup_1550), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix17183 (.Y (nx17182), .A0 (rd_addr_m_1), .A1 (nx2219)
                          , .B0 (nx2221), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2846 (.Y (nx2219), .A (modgen_ram_ix167_a_40__dup_1557)
                      , .B (modgen_ram_ix167_a_41__dup_1556), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2847 (.Y (nx2221), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_1554), .B0 (nx17164), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix17165 (.Y (nx17164), .AN (
                      modgen_ram_ix167_a_42__dup_1555), .B (rd_addr_m_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_5 (.Q (rd_data_m_5), .CK (wb_clk_i), .D (
                        nx23750), .R (wb_rst_i), .SE (NOT_nx50), .SI (
                        rd_data_m_5)) ;
    MXIT2_X0P5M_A12TS ix23751 (.Y (nx23750), .A (nx3454), .B (nx2229), .S0 (
                      nx1127)) ;
    INV_X0P5B_A12TS ix2848 (.Y (nx3454), .A (wr_data_m_5)) ;
    OA21A1OI2_X0P5M_A12TS ix2849 (.Y (nx2229), .A0 (nx23736), .A1 (nx22846), .B0 (
                          rd_addr_7), .C0 (nx21954)) ;
    OA21A1OI2_X0P5M_A12TS ix23737 (.Y (nx23736), .A0 (rd_addr_m_5), .A1 (nx2233)
                          , .B0 (nx3459), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2850 (.Y (nx2233), .A0 (rd_addr_m_4), .A1 (nx23282), .B0 (
                      nx23066)) ;
    MXT4_X0P5M_A12TS ix23283 (.Y (nx23282), .A (nx23114), .B (nx23222), .C (
                     nx23166), .D (nx23274), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix23115 (.Y (nx23114), .A (modgen_ram_ix167_a_208__dup_1125
                     ), .B (modgen_ram_ix167_a_210__dup_1123), .C (
                     modgen_ram_ix167_a_209__dup_1124), .D (
                     modgen_ram_ix167_a_211__dup_1122), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix23223 (.Y (nx23222), .A (modgen_ram_ix167_a_216__dup_1117
                     ), .B (modgen_ram_ix167_a_218__dup_1115), .C (
                     modgen_ram_ix167_a_217__dup_1116), .D (
                     modgen_ram_ix167_a_219__dup_1114), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix23167 (.Y (nx23166), .A (modgen_ram_ix167_a_212__dup_1121
                     ), .B (modgen_ram_ix167_a_214__dup_1119), .C (
                     modgen_ram_ix167_a_213__dup_1120), .D (
                     modgen_ram_ix167_a_215__dup_1118), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix23275 (.Y (nx23274), .A (modgen_ram_ix167_a_220__dup_1113
                     ), .B (modgen_ram_ix167_a_222__dup_1111), .C (
                     modgen_ram_ix167_a_221__dup_1112), .D (
                     modgen_ram_ix167_a_223__dup_1110), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23067 (.Y (nx23066), .A0 (rd_addr_m_3), .A1 (nx3455)
                          , .B0 (nx3456), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2852 (.Y (nx3455), .A0 (rd_addr_m_2), .A1 (nx22946), .B0 (
                      nx22898)) ;
    MXT4_X0P5M_A12TS ix22947 (.Y (nx22946), .A (modgen_ram_ix167_a_196__dup_1137
                     ), .B (modgen_ram_ix167_a_198__dup_1135), .C (
                     modgen_ram_ix167_a_197__dup_1136), .D (
                     modgen_ram_ix167_a_199__dup_1134), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22899 (.Y (nx22898), .A0 (rd_addr_m_1), .A1 (nx2253)
                          , .B0 (nx2255), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2853 (.Y (nx2253), .A (modgen_ram_ix167_a_192__dup_1141)
                      , .B (modgen_ram_ix167_a_193__dup_1140), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2854 (.Y (nx2255), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_1138), .B0 (nx22880), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix22881 (.Y (nx22880), .AN (
                      modgen_ram_ix167_a_194__dup_1139), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2855 (.Y (nx3456), .A0 (rd_addr_m_2), .A1 (nx23054)
                          , .B0 (nx23006), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix23055 (.Y (nx23054), .A (modgen_ram_ix167_a_204__dup_1129
                     ), .B (modgen_ram_ix167_a_206__dup_1127), .C (
                     modgen_ram_ix167_a_205__dup_1128), .D (
                     modgen_ram_ix167_a_207__dup_1126), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23007 (.Y (nx23006), .A0 (rd_addr_m_1), .A1 (nx3457)
                          , .B0 (nx2267), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2856 (.Y (nx3457), .A (modgen_ram_ix167_a_200__dup_1133)
                      , .B (modgen_ram_ix167_a_201__dup_1132), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2858 (.Y (nx2267), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_1130), .B0 (nx22988), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix22989 (.Y (nx22988), .AN (
                      modgen_ram_ix167_a_202__dup_1131), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2860 (.Y (nx3459), .A0 (rd_addr_m_4), .A1 (nx23726)
                          , .B0 (nx23510), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix23727 (.Y (nx23726), .A (nx23558), .B (nx23666), .C (
                     nx23610), .D (nx23718), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix23559 (.Y (nx23558), .A (modgen_ram_ix167_a_240__dup_1093
                     ), .B (modgen_ram_ix167_a_242__dup_1091), .C (
                     modgen_ram_ix167_a_241__dup_1092), .D (
                     modgen_ram_ix167_a_243__dup_1090), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix23667 (.Y (nx23666), .A (modgen_ram_ix167_a_248__dup_1085
                     ), .B (modgen_ram_ix167_a_250__dup_1083), .C (
                     modgen_ram_ix167_a_249__dup_1084), .D (
                     modgen_ram_ix167_a_251__dup_1082), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix23611 (.Y (nx23610), .A (modgen_ram_ix167_a_244__dup_1089
                     ), .B (modgen_ram_ix167_a_246__dup_1087), .C (
                     modgen_ram_ix167_a_245__dup_1088), .D (
                     modgen_ram_ix167_a_247__dup_1086), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix23719 (.Y (nx23718), .A (modgen_ram_ix167_a_252__dup_1081
                     ), .B (modgen_ram_ix167_a_254__dup_1079), .C (
                     modgen_ram_ix167_a_253__dup_1080), .D (
                     modgen_ram_ix167_a_255__dup_1078), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23511 (.Y (nx23510), .A0 (rd_addr_m_3), .A1 (nx2281)
                          , .B0 (nx2291), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2861 (.Y (nx2281), .A0 (rd_addr_m_2), .A1 (nx23390), .B0 (
                      nx23342)) ;
    MXT4_X0P5M_A12TS ix23391 (.Y (nx23390), .A (modgen_ram_ix167_a_228__dup_1105
                     ), .B (modgen_ram_ix167_a_230__dup_1103), .C (
                     modgen_ram_ix167_a_229__dup_1104), .D (
                     modgen_ram_ix167_a_231__dup_1102), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23343 (.Y (nx23342), .A0 (rd_addr_m_1), .A1 (nx2285)
                          , .B0 (nx2287), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2862 (.Y (nx2285), .A (modgen_ram_ix167_a_224__dup_1109)
                      , .B (modgen_ram_ix167_a_225__dup_1108), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2863 (.Y (nx2287), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_1106), .B0 (nx23324), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix23325 (.Y (nx23324), .AN (
                      modgen_ram_ix167_a_226__dup_1107), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2864 (.Y (nx2291), .A0 (rd_addr_m_2), .A1 (nx23498)
                          , .B0 (nx23450), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix23499 (.Y (nx23498), .A (modgen_ram_ix167_a_236__dup_1097
                     ), .B (modgen_ram_ix167_a_238__dup_1095), .C (
                     modgen_ram_ix167_a_237__dup_1096), .D (
                     modgen_ram_ix167_a_239__dup_1094), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23451 (.Y (nx23450), .A0 (rd_addr_m_1), .A1 (nx2295)
                          , .B0 (nx2297), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2865 (.Y (nx2295), .A (modgen_ram_ix167_a_232__dup_1101)
                      , .B (modgen_ram_ix167_a_233__dup_1100), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2866 (.Y (nx2297), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_1098), .B0 (nx23432), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix23433 (.Y (nx23432), .AN (
                      modgen_ram_ix167_a_234__dup_1099), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22847 (.Y (nx22846), .A0 (rd_addr_m_5), .A1 (nx3460)
                          , .B0 (nx3462), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2867 (.Y (nx3460), .A0 (rd_addr_m_4), .A1 (nx22390), .B0 (
                      nx22174)) ;
    MXT4_X0P5M_A12TS ix22391 (.Y (nx22390), .A (nx22222), .B (nx22330), .C (
                     nx22274), .D (nx22382), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix22223 (.Y (nx22222), .A (modgen_ram_ix167_a_144__dup_1189
                     ), .B (modgen_ram_ix167_a_146__dup_1187), .C (
                     modgen_ram_ix167_a_145__dup_1188), .D (
                     modgen_ram_ix167_a_147__dup_1186), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix22331 (.Y (nx22330), .A (modgen_ram_ix167_a_152__dup_1181
                     ), .B (modgen_ram_ix167_a_154__dup_1179), .C (
                     modgen_ram_ix167_a_153__dup_1180), .D (
                     modgen_ram_ix167_a_155__dup_1178), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix22275 (.Y (nx22274), .A (modgen_ram_ix167_a_148__dup_1185
                     ), .B (modgen_ram_ix167_a_150__dup_1183), .C (
                     modgen_ram_ix167_a_149__dup_1184), .D (
                     modgen_ram_ix167_a_151__dup_1182), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix22383 (.Y (nx22382), .A (modgen_ram_ix167_a_156__dup_1177
                     ), .B (modgen_ram_ix167_a_158__dup_1175), .C (
                     modgen_ram_ix167_a_157__dup_1176), .D (
                     modgen_ram_ix167_a_159__dup_1174), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22175 (.Y (nx22174), .A0 (rd_addr_m_3), .A1 (nx2311)
                          , .B0 (nx2323), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2868 (.Y (nx2311), .A0 (rd_addr_m_2), .A1 (nx22054), .B0 (
                      nx22006)) ;
    MXT4_X0P5M_A12TS ix22055 (.Y (nx22054), .A (modgen_ram_ix167_a_132__dup_1201
                     ), .B (modgen_ram_ix167_a_134__dup_1199), .C (
                     modgen_ram_ix167_a_133__dup_1200), .D (
                     modgen_ram_ix167_a_135__dup_1198), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22007 (.Y (nx22006), .A0 (rd_addr_m_1), .A1 (nx3461)
                          , .B0 (nx2319), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2869 (.Y (nx3461), .A (modgen_ram_ix167_a_128__dup_1205)
                      , .B (modgen_ram_ix167_a_129__dup_1204), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2320 (.Y (nx2319), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_1202), .B0 (nx21988), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix21989 (.Y (nx21988), .AN (
                      modgen_ram_ix167_a_130__dup_1203), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2324 (.Y (nx2323), .A0 (rd_addr_m_2), .A1 (nx22162)
                          , .B0 (nx22114), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix22163 (.Y (nx22162), .A (modgen_ram_ix167_a_140__dup_1193
                     ), .B (modgen_ram_ix167_a_142__dup_1191), .C (
                     modgen_ram_ix167_a_141__dup_1192), .D (
                     modgen_ram_ix167_a_143__dup_1190), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22115 (.Y (nx22114), .A0 (rd_addr_m_1), .A1 (nx2327)
                          , .B0 (nx2329), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2328 (.Y (nx2327), .A (modgen_ram_ix167_a_136__dup_1197)
                      , .B (modgen_ram_ix167_a_137__dup_1196), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2330 (.Y (nx2329), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_1194), .B0 (nx22096), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix22097 (.Y (nx22096), .AN (
                      modgen_ram_ix167_a_138__dup_1195), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2870 (.Y (nx3462), .A0 (rd_addr_m_4), .A1 (nx22834)
                          , .B0 (nx22618), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix22835 (.Y (nx22834), .A (nx22666), .B (nx22774), .C (
                     nx22718), .D (nx22826), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix22667 (.Y (nx22666), .A (modgen_ram_ix167_a_176__dup_1157
                     ), .B (modgen_ram_ix167_a_178__dup_1155), .C (
                     modgen_ram_ix167_a_177__dup_1156), .D (
                     modgen_ram_ix167_a_179__dup_1154), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix22775 (.Y (nx22774), .A (modgen_ram_ix167_a_184__dup_1149
                     ), .B (modgen_ram_ix167_a_186__dup_1147), .C (
                     modgen_ram_ix167_a_185__dup_1148), .D (
                     modgen_ram_ix167_a_187__dup_1146), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix22719 (.Y (nx22718), .A (modgen_ram_ix167_a_180__dup_1153
                     ), .B (modgen_ram_ix167_a_182__dup_1151), .C (
                     modgen_ram_ix167_a_181__dup_1152), .D (
                     modgen_ram_ix167_a_183__dup_1150), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix22827 (.Y (nx22826), .A (modgen_ram_ix167_a_188__dup_1145
                     ), .B (modgen_ram_ix167_a_190__dup_1143), .C (
                     modgen_ram_ix167_a_189__dup_1144), .D (
                     modgen_ram_ix167_a_191__dup_1142), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22619 (.Y (nx22618), .A0 (rd_addr_m_3), .A1 (nx3463)
                          , .B0 (nx3465), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2871 (.Y (nx3463), .A0 (rd_addr_m_2), .A1 (nx22498), .B0 (
                      nx22450)) ;
    MXT4_X0P5M_A12TS ix22499 (.Y (nx22498), .A (modgen_ram_ix167_a_164__dup_1169
                     ), .B (modgen_ram_ix167_a_166__dup_1167), .C (
                     modgen_ram_ix167_a_165__dup_1168), .D (
                     modgen_ram_ix167_a_167__dup_1166), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22451 (.Y (nx22450), .A0 (rd_addr_m_1), .A1 (nx3464)
                          , .B0 (nx2349), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2872 (.Y (nx3464), .A (modgen_ram_ix167_a_160__dup_1173)
                      , .B (modgen_ram_ix167_a_161__dup_1172), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2350 (.Y (nx2349), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_1170), .B0 (nx22432), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix22433 (.Y (nx22432), .AN (
                      modgen_ram_ix167_a_162__dup_1171), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2873 (.Y (nx3465), .A0 (rd_addr_m_2), .A1 (nx22606)
                          , .B0 (nx22558), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix22607 (.Y (nx22606), .A (modgen_ram_ix167_a_172__dup_1161
                     ), .B (modgen_ram_ix167_a_174__dup_1159), .C (
                     modgen_ram_ix167_a_173__dup_1160), .D (
                     modgen_ram_ix167_a_175__dup_1158), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix22559 (.Y (nx22558), .A0 (rd_addr_m_1), .A1 (nx3466)
                          , .B0 (nx3467), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2874 (.Y (nx3466), .A (modgen_ram_ix167_a_168__dup_1165)
                      , .B (modgen_ram_ix167_a_169__dup_1164), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2876 (.Y (nx3467), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_1162), .B0 (nx22540), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix22541 (.Y (nx22540), .AN (
                      modgen_ram_ix167_a_170__dup_1163), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix21955 (.Y (nx21954), .A (rd_addr_7), .B (nx3468)) ;
    AOI21_X0P5M_A12TS ix2366 (.Y (nx3468), .A0 (rd_addr_m_6), .A1 (nx21946), .B0 (
                      nx21058)) ;
    OAI21_X0P5M_A12TS ix21947 (.Y (nx21946), .A0 (rd_addr_m_5), .A1 (nx3469), .B0 (
                      nx3478)) ;
    AOI21_X0P5M_A12TS ix2877 (.Y (nx3469), .A0 (rd_addr_m_4), .A1 (nx21494), .B0 (
                      nx21278)) ;
    MXT4_X0P5M_A12TS ix21495 (.Y (nx21494), .A (nx21326), .B (nx21434), .C (
                     nx21378), .D (nx21486), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix21327 (.Y (nx21326), .A (modgen_ram_ix167_a_80__dup_1253)
                     , .B (modgen_ram_ix167_a_82__dup_1251), .C (
                     modgen_ram_ix167_a_81__dup_1252), .D (
                     modgen_ram_ix167_a_83__dup_1250), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21435 (.Y (nx21434), .A (modgen_ram_ix167_a_88__dup_1245)
                     , .B (modgen_ram_ix167_a_90__dup_1243), .C (
                     modgen_ram_ix167_a_89__dup_1244), .D (
                     modgen_ram_ix167_a_91__dup_1242), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21379 (.Y (nx21378), .A (modgen_ram_ix167_a_84__dup_1249)
                     , .B (modgen_ram_ix167_a_86__dup_1247), .C (
                     modgen_ram_ix167_a_85__dup_1248), .D (
                     modgen_ram_ix167_a_87__dup_1246), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21487 (.Y (nx21486), .A (modgen_ram_ix167_a_92__dup_1241)
                     , .B (modgen_ram_ix167_a_94__dup_1239), .C (
                     modgen_ram_ix167_a_93__dup_1240), .D (
                     modgen_ram_ix167_a_95__dup_1238), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21279 (.Y (nx21278), .A0 (rd_addr_m_3), .A1 (nx3470)
                          , .B0 (nx3474), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2380 (.Y (nx3470), .A0 (rd_addr_m_2), .A1 (nx21158), .B0 (
                      nx21110)) ;
    MXT4_X0P5M_A12TS ix21159 (.Y (nx21158), .A (modgen_ram_ix167_a_68__dup_1265)
                     , .B (modgen_ram_ix167_a_70__dup_1263), .C (
                     modgen_ram_ix167_a_69__dup_1264), .D (
                     modgen_ram_ix167_a_71__dup_1262), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21111 (.Y (nx21110), .A0 (rd_addr_m_1), .A1 (nx3471)
                          , .B0 (nx3473), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2878 (.Y (nx3471), .A (modgen_ram_ix167_a_64__dup_1269)
                      , .B (modgen_ram_ix167_a_65__dup_1268), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2879 (.Y (nx3473), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_1266), .B0 (nx21092), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix21093 (.Y (nx21092), .AN (
                      modgen_ram_ix167_a_66__dup_1267), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2880 (.Y (nx3474), .A0 (rd_addr_m_2), .A1 (nx21266)
                          , .B0 (nx21218), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix21267 (.Y (nx21266), .A (modgen_ram_ix167_a_76__dup_1257)
                     , .B (modgen_ram_ix167_a_78__dup_1255), .C (
                     modgen_ram_ix167_a_77__dup_1256), .D (
                     modgen_ram_ix167_a_79__dup_1254), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21219 (.Y (nx21218), .A0 (rd_addr_m_1), .A1 (nx3475)
                          , .B0 (nx3477), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2394 (.Y (nx3475), .A (modgen_ram_ix167_a_72__dup_1261)
                      , .B (modgen_ram_ix167_a_73__dup_1260), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2396 (.Y (nx3477), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_1258), .B0 (nx21200), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix21201 (.Y (nx21200), .AN (
                      modgen_ram_ix167_a_74__dup_1259), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2400 (.Y (nx3478), .A0 (rd_addr_m_4), .A1 (nx21938)
                          , .B0 (nx21722), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix21939 (.Y (nx21938), .A (nx21770), .B (nx21878), .C (
                     nx21822), .D (nx21930), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix21771 (.Y (nx21770), .A (modgen_ram_ix167_a_112__dup_1221
                     ), .B (modgen_ram_ix167_a_114__dup_1219), .C (
                     modgen_ram_ix167_a_113__dup_1220), .D (
                     modgen_ram_ix167_a_115__dup_1218), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21879 (.Y (nx21878), .A (modgen_ram_ix167_a_120__dup_1213
                     ), .B (modgen_ram_ix167_a_122__dup_1211), .C (
                     modgen_ram_ix167_a_121__dup_1212), .D (
                     modgen_ram_ix167_a_123__dup_1210), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21823 (.Y (nx21822), .A (modgen_ram_ix167_a_116__dup_1217
                     ), .B (modgen_ram_ix167_a_118__dup_1215), .C (
                     modgen_ram_ix167_a_117__dup_1216), .D (
                     modgen_ram_ix167_a_119__dup_1214), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21931 (.Y (nx21930), .A (modgen_ram_ix167_a_124__dup_1209
                     ), .B (modgen_ram_ix167_a_126__dup_1207), .C (
                     modgen_ram_ix167_a_125__dup_1208), .D (
                     modgen_ram_ix167_a_127__dup_1206), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21723 (.Y (nx21722), .A0 (rd_addr_m_3), .A1 (nx3479)
                          , .B0 (nx3482), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2881 (.Y (nx3479), .A0 (rd_addr_m_2), .A1 (nx21602), .B0 (
                      nx21554)) ;
    MXT4_X0P5M_A12TS ix21603 (.Y (nx21602), .A (modgen_ram_ix167_a_100__dup_1233
                     ), .B (modgen_ram_ix167_a_102__dup_1231), .C (
                     modgen_ram_ix167_a_101__dup_1232), .D (
                     modgen_ram_ix167_a_103__dup_1230), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21555 (.Y (nx21554), .A0 (rd_addr_m_1), .A1 (nx3480)
                          , .B0 (nx3481), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2414 (.Y (nx3480), .A (modgen_ram_ix167_a_96__dup_1237)
                      , .B (modgen_ram_ix167_a_97__dup_1236), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2416 (.Y (nx3481), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_1234), .B0 (nx21536), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix21537 (.Y (nx21536), .AN (
                      modgen_ram_ix167_a_98__dup_1235), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2420 (.Y (nx3482), .A0 (rd_addr_m_2), .A1 (nx21710)
                          , .B0 (nx21662), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix21711 (.Y (nx21710), .A (modgen_ram_ix167_a_108__dup_1225
                     ), .B (modgen_ram_ix167_a_110__dup_1223), .C (
                     modgen_ram_ix167_a_109__dup_1224), .D (
                     modgen_ram_ix167_a_111__dup_1222), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21663 (.Y (nx21662), .A0 (rd_addr_m_1), .A1 (nx3483)
                          , .B0 (nx3485), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2882 (.Y (nx3483), .A (modgen_ram_ix167_a_104__dup_1229)
                      , .B (modgen_ram_ix167_a_105__dup_1228), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2883 (.Y (nx3485), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_1226), .B0 (nx21644), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix21645 (.Y (nx21644), .AN (
                      modgen_ram_ix167_a_106__dup_1227), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix21059 (.Y (nx21058), .A0 (rd_addr_m_5), .A1 (nx3487)
                          , .B0 (nx2461), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2884 (.Y (nx3487), .A0 (rd_addr_m_4), .A1 (nx20602), .B0 (
                      nx20386)) ;
    MXT4_X0P5M_A12TS ix20603 (.Y (nx20602), .A (nx20434), .B (nx20542), .C (
                     nx20486), .D (nx20594), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix20435 (.Y (nx20434), .A (modgen_ram_ix167_a_16__dup_1317)
                     , .B (modgen_ram_ix167_a_18__dup_1315), .C (
                     modgen_ram_ix167_a_17__dup_1316), .D (
                     modgen_ram_ix167_a_19__dup_1314), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20543 (.Y (nx20542), .A (modgen_ram_ix167_a_24__dup_1309)
                     , .B (modgen_ram_ix167_a_26__dup_1307), .C (
                     modgen_ram_ix167_a_25__dup_1308), .D (
                     modgen_ram_ix167_a_27__dup_1306), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20487 (.Y (nx20486), .A (modgen_ram_ix167_a_20__dup_1313)
                     , .B (modgen_ram_ix167_a_22__dup_1311), .C (
                     modgen_ram_ix167_a_21__dup_1312), .D (
                     modgen_ram_ix167_a_23__dup_1310), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20595 (.Y (nx20594), .A (modgen_ram_ix167_a_28__dup_1305)
                     , .B (modgen_ram_ix167_a_30__dup_1303), .C (
                     modgen_ram_ix167_a_29__dup_1304), .D (
                     modgen_ram_ix167_a_31__dup_1302), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix20387 (.Y (nx20386), .A0 (rd_addr_m_3), .A1 (nx3488)
                          , .B0 (nx2451), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2441 (.Y (nx3488), .A0 (rd_addr_m_2), .A1 (nx20266), .B0 (
                      nx20218)) ;
    MXT4_X0P5M_A12TS ix20267 (.Y (nx20266), .A (modgen_ram_ix167_a_4__dup_1329)
                     , .B (modgen_ram_ix167_a_6__dup_1327), .C (
                     modgen_ram_ix167_a_5__dup_1328), .D (
                     modgen_ram_ix167_a_7__dup_1326), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix20219 (.Y (nx20218), .A0 (rd_addr_m_1), .A1 (nx3489)
                          , .B0 (nx3490), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2886 (.Y (nx3489), .A (modgen_ram_ix167_a_0__dup_1333), 
                      .B (modgen_ram_ix167_a_1__dup_1332), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2887 (.Y (nx3490), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_1330), .B0 (nx20200), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix20201 (.Y (nx20200), .AN (modgen_ram_ix167_a_2__dup_1331
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2888 (.Y (nx2451), .A0 (rd_addr_m_2), .A1 (nx20374)
                          , .B0 (nx20326), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix20375 (.Y (nx20374), .A (modgen_ram_ix167_a_12__dup_1321)
                     , .B (modgen_ram_ix167_a_14__dup_1319), .C (
                     modgen_ram_ix167_a_13__dup_1320), .D (
                     modgen_ram_ix167_a_15__dup_1318), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix20327 (.Y (nx20326), .A0 (rd_addr_m_1), .A1 (nx2456)
                          , .B0 (nx3491), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2889 (.Y (nx2456), .A (modgen_ram_ix167_a_8__dup_1325), 
                      .B (modgen_ram_ix167_a_9__dup_1324), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2890 (.Y (nx3491), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_1322), .B0 (nx20308), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix20309 (.Y (nx20308), .AN (
                      modgen_ram_ix167_a_10__dup_1323), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2891 (.Y (nx2461), .A0 (rd_addr_m_4), .A1 (nx21046)
                          , .B0 (nx20830), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix21047 (.Y (nx21046), .A (nx20878), .B (nx20986), .C (
                     nx20930), .D (nx21038), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix20879 (.Y (nx20878), .A (modgen_ram_ix167_a_48__dup_1285)
                     , .B (modgen_ram_ix167_a_50__dup_1283), .C (
                     modgen_ram_ix167_a_49__dup_1284), .D (
                     modgen_ram_ix167_a_51__dup_1282), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20987 (.Y (nx20986), .A (modgen_ram_ix167_a_56__dup_1277)
                     , .B (modgen_ram_ix167_a_58__dup_1275), .C (
                     modgen_ram_ix167_a_57__dup_1276), .D (
                     modgen_ram_ix167_a_59__dup_1274), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix20931 (.Y (nx20930), .A (modgen_ram_ix167_a_52__dup_1281)
                     , .B (modgen_ram_ix167_a_54__dup_1279), .C (
                     modgen_ram_ix167_a_53__dup_1280), .D (
                     modgen_ram_ix167_a_55__dup_1278), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix21039 (.Y (nx21038), .A (modgen_ram_ix167_a_60__dup_1273)
                     , .B (modgen_ram_ix167_a_62__dup_1271), .C (
                     modgen_ram_ix167_a_61__dup_1272), .D (
                     modgen_ram_ix167_a_63__dup_1270), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix20831 (.Y (nx20830), .A0 (rd_addr_m_3), .A1 (nx3492)
                          , .B0 (nx2480), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2892 (.Y (nx3492), .A0 (rd_addr_m_2), .A1 (nx20710), .B0 (
                      nx20662)) ;
    MXT4_X0P5M_A12TS ix20711 (.Y (nx20710), .A (modgen_ram_ix167_a_36__dup_1297)
                     , .B (modgen_ram_ix167_a_38__dup_1295), .C (
                     modgen_ram_ix167_a_37__dup_1296), .D (
                     modgen_ram_ix167_a_39__dup_1294), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix20663 (.Y (nx20662), .A0 (rd_addr_m_1), .A1 (nx2475)
                          , .B0 (nx2477), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2894 (.Y (nx2475), .A (modgen_ram_ix167_a_32__dup_1301)
                      , .B (modgen_ram_ix167_a_33__dup_1300), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2895 (.Y (nx2477), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_1298), .B0 (nx20644), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix20645 (.Y (nx20644), .AN (
                      modgen_ram_ix167_a_34__dup_1299), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2896 (.Y (nx2480), .A0 (rd_addr_m_2), .A1 (nx20818)
                          , .B0 (nx20770), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix20819 (.Y (nx20818), .A (modgen_ram_ix167_a_44__dup_1289)
                     , .B (modgen_ram_ix167_a_46__dup_1287), .C (
                     modgen_ram_ix167_a_45__dup_1288), .D (
                     modgen_ram_ix167_a_47__dup_1286), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix20771 (.Y (nx20770), .A0 (rd_addr_m_1), .A1 (nx2485)
                          , .B0 (nx2487), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2897 (.Y (nx2485), .A (modgen_ram_ix167_a_40__dup_1293)
                      , .B (modgen_ram_ix167_a_41__dup_1292), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2898 (.Y (nx2487), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_1290), .B0 (nx20752), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix20753 (.Y (nx20752), .AN (
                      modgen_ram_ix167_a_42__dup_1291), .B (rd_addr_m_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_6 (.Q (rd_data_m_6), .CK (wb_clk_i), .D (
                        nx27338), .R (wb_rst_i), .SE (NOT_nx50), .SI (
                        rd_data_m_6)) ;
    MXIT2_X0P5M_A12TS ix27339 (.Y (nx27338), .A (nx2493), .B (nx3493), .S0 (
                      nx1127)) ;
    INV_X0P5B_A12TS ix2900 (.Y (nx2493), .A (wr_data_m_6)) ;
    OA21A1OI2_X0P5M_A12TS ix2901 (.Y (nx3493), .A0 (nx27324), .A1 (nx26434), .B0 (
                          rd_addr_7), .C0 (nx25542)) ;
    OA21A1OI2_X0P5M_A12TS ix27325 (.Y (nx27324), .A0 (rd_addr_m_5), .A1 (nx2498)
                          , .B0 (nx2531), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2902 (.Y (nx2498), .A0 (rd_addr_m_4), .A1 (nx26870), .B0 (
                      nx26654)) ;
    MXT4_X0P5M_A12TS ix26871 (.Y (nx26870), .A (nx26702), .B (nx26810), .C (
                     nx26754), .D (nx26862), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix26703 (.Y (nx26702), .A (modgen_ram_ix167_a_208__dup_861)
                     , .B (modgen_ram_ix167_a_210__dup_859), .C (
                     modgen_ram_ix167_a_209__dup_860), .D (
                     modgen_ram_ix167_a_211__dup_858), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix26811 (.Y (nx26810), .A (modgen_ram_ix167_a_216__dup_853)
                     , .B (modgen_ram_ix167_a_218__dup_851), .C (
                     modgen_ram_ix167_a_217__dup_852), .D (
                     modgen_ram_ix167_a_219__dup_850), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix26755 (.Y (nx26754), .A (modgen_ram_ix167_a_212__dup_857)
                     , .B (modgen_ram_ix167_a_214__dup_855), .C (
                     modgen_ram_ix167_a_213__dup_856), .D (
                     modgen_ram_ix167_a_215__dup_854), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix26863 (.Y (nx26862), .A (modgen_ram_ix167_a_220__dup_849)
                     , .B (modgen_ram_ix167_a_222__dup_847), .C (
                     modgen_ram_ix167_a_221__dup_848), .D (
                     modgen_ram_ix167_a_223__dup_846), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26655 (.Y (nx26654), .A0 (rd_addr_m_3), .A1 (nx2511)
                          , .B0 (nx3495), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2903 (.Y (nx2511), .A0 (rd_addr_m_2), .A1 (nx26534), .B0 (
                      nx26486)) ;
    MXT4_X0P5M_A12TS ix26535 (.Y (nx26534), .A (modgen_ram_ix167_a_196__dup_873)
                     , .B (modgen_ram_ix167_a_198__dup_871), .C (
                     modgen_ram_ix167_a_197__dup_872), .D (
                     modgen_ram_ix167_a_199__dup_870), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26487 (.Y (nx26486), .A0 (rd_addr_m_1), .A1 (nx3494)
                          , .B0 (nx2517), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2904 (.Y (nx3494), .A (modgen_ram_ix167_a_192__dup_877)
                      , .B (modgen_ram_ix167_a_193__dup_876), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2906 (.Y (nx2517), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195__dup_874), .B0 (nx26468), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix26469 (.Y (nx26468), .AN (
                      modgen_ram_ix167_a_194__dup_875), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2907 (.Y (nx3495), .A0 (rd_addr_m_2), .A1 (nx26642)
                          , .B0 (nx26594), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix26643 (.Y (nx26642), .A (modgen_ram_ix167_a_204__dup_865)
                     , .B (modgen_ram_ix167_a_206__dup_863), .C (
                     modgen_ram_ix167_a_205__dup_864), .D (
                     modgen_ram_ix167_a_207__dup_862), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26595 (.Y (nx26594), .A0 (rd_addr_m_1), .A1 (nx2525)
                          , .B0 (nx2527), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2908 (.Y (nx2525), .A (modgen_ram_ix167_a_200__dup_869)
                      , .B (modgen_ram_ix167_a_201__dup_868), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2909 (.Y (nx2527), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203__dup_866), .B0 (nx26576), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix26577 (.Y (nx26576), .AN (
                      modgen_ram_ix167_a_202__dup_867), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2910 (.Y (nx2531), .A0 (rd_addr_m_4), .A1 (nx27314)
                          , .B0 (nx27098), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix27315 (.Y (nx27314), .A (nx27146), .B (nx27254), .C (
                     nx27198), .D (nx27306), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix27147 (.Y (nx27146), .A (modgen_ram_ix167_a_240__dup_829)
                     , .B (modgen_ram_ix167_a_242__dup_827), .C (
                     modgen_ram_ix167_a_241__dup_828), .D (
                     modgen_ram_ix167_a_243__dup_826), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix27255 (.Y (nx27254), .A (modgen_ram_ix167_a_248__dup_821)
                     , .B (modgen_ram_ix167_a_250__dup_819), .C (
                     modgen_ram_ix167_a_249__dup_820), .D (
                     modgen_ram_ix167_a_251__dup_818), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix27199 (.Y (nx27198), .A (modgen_ram_ix167_a_244__dup_825)
                     , .B (modgen_ram_ix167_a_246__dup_823), .C (
                     modgen_ram_ix167_a_245__dup_824), .D (
                     modgen_ram_ix167_a_247__dup_822), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix27307 (.Y (nx27306), .A (modgen_ram_ix167_a_252__dup_817)
                     , .B (modgen_ram_ix167_a_254__dup_815), .C (
                     modgen_ram_ix167_a_253__dup_816), .D (
                     modgen_ram_ix167_a_255__dup_814), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix27099 (.Y (nx27098), .A0 (rd_addr_m_3), .A1 (nx2541)
                          , .B0 (nx2551), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2911 (.Y (nx2541), .A0 (rd_addr_m_2), .A1 (nx26978), .B0 (
                      nx26930)) ;
    MXT4_X0P5M_A12TS ix26979 (.Y (nx26978), .A (modgen_ram_ix167_a_228__dup_841)
                     , .B (modgen_ram_ix167_a_230__dup_839), .C (
                     modgen_ram_ix167_a_229__dup_840), .D (
                     modgen_ram_ix167_a_231__dup_838), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26931 (.Y (nx26930), .A0 (rd_addr_m_1), .A1 (nx2545)
                          , .B0 (nx2547), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2912 (.Y (nx2545), .A (modgen_ram_ix167_a_224__dup_845)
                      , .B (modgen_ram_ix167_a_225__dup_844), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2913 (.Y (nx2547), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227__dup_842), .B0 (nx26912), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix26913 (.Y (nx26912), .AN (
                      modgen_ram_ix167_a_226__dup_843), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2914 (.Y (nx2551), .A0 (rd_addr_m_2), .A1 (nx27086)
                          , .B0 (nx27038), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix27087 (.Y (nx27086), .A (modgen_ram_ix167_a_236__dup_833)
                     , .B (modgen_ram_ix167_a_238__dup_831), .C (
                     modgen_ram_ix167_a_237__dup_832), .D (
                     modgen_ram_ix167_a_239__dup_830), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix27039 (.Y (nx27038), .A0 (rd_addr_m_1), .A1 (nx2555)
                          , .B0 (nx3497), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2915 (.Y (nx2555), .A (modgen_ram_ix167_a_232__dup_837)
                      , .B (modgen_ram_ix167_a_233__dup_836), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2916 (.Y (nx3497), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235__dup_834), .B0 (nx27020), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix27021 (.Y (nx27020), .AN (
                      modgen_ram_ix167_a_234__dup_835), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26435 (.Y (nx26434), .A0 (rd_addr_m_5), .A1 (nx3498)
                          , .B0 (nx2593), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2918 (.Y (nx3498), .A0 (rd_addr_m_4), .A1 (nx25978), .B0 (
                      nx25762)) ;
    MXT4_X0P5M_A12TS ix25979 (.Y (nx25978), .A (nx25810), .B (nx25918), .C (
                     nx25862), .D (nx25970), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix25811 (.Y (nx25810), .A (modgen_ram_ix167_a_144__dup_925)
                     , .B (modgen_ram_ix167_a_146__dup_923), .C (
                     modgen_ram_ix167_a_145__dup_924), .D (
                     modgen_ram_ix167_a_147__dup_922), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25919 (.Y (nx25918), .A (modgen_ram_ix167_a_152__dup_917)
                     , .B (modgen_ram_ix167_a_154__dup_915), .C (
                     modgen_ram_ix167_a_153__dup_916), .D (
                     modgen_ram_ix167_a_155__dup_914), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25863 (.Y (nx25862), .A (modgen_ram_ix167_a_148__dup_921)
                     , .B (modgen_ram_ix167_a_150__dup_919), .C (
                     modgen_ram_ix167_a_149__dup_920), .D (
                     modgen_ram_ix167_a_151__dup_918), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25971 (.Y (nx25970), .A (modgen_ram_ix167_a_156__dup_913)
                     , .B (modgen_ram_ix167_a_158__dup_911), .C (
                     modgen_ram_ix167_a_157__dup_912), .D (
                     modgen_ram_ix167_a_159__dup_910), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix25763 (.Y (nx25762), .A0 (rd_addr_m_3), .A1 (nx2571)
                          , .B0 (nx3499), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2919 (.Y (nx2571), .A0 (rd_addr_m_2), .A1 (nx25642), .B0 (
                      nx25594)) ;
    MXT4_X0P5M_A12TS ix25643 (.Y (nx25642), .A (modgen_ram_ix167_a_132__dup_937)
                     , .B (modgen_ram_ix167_a_134__dup_935), .C (
                     modgen_ram_ix167_a_133__dup_936), .D (
                     modgen_ram_ix167_a_135__dup_934), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix25595 (.Y (nx25594), .A0 (rd_addr_m_1), .A1 (nx2577)
                          , .B0 (nx2579), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2920 (.Y (nx2577), .A (modgen_ram_ix167_a_128__dup_941)
                      , .B (modgen_ram_ix167_a_129__dup_940), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2921 (.Y (nx2579), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131__dup_938), .B0 (nx25576), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix25577 (.Y (nx25576), .AN (
                      modgen_ram_ix167_a_130__dup_939), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2922 (.Y (nx3499), .A0 (rd_addr_m_2), .A1 (nx25750)
                          , .B0 (nx25702), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix25751 (.Y (nx25750), .A (modgen_ram_ix167_a_140__dup_929)
                     , .B (modgen_ram_ix167_a_142__dup_927), .C (
                     modgen_ram_ix167_a_141__dup_928), .D (
                     modgen_ram_ix167_a_143__dup_926), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix25703 (.Y (nx25702), .A0 (rd_addr_m_1), .A1 (nx3500)
                          , .B0 (nx3501), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2923 (.Y (nx3500), .A (modgen_ram_ix167_a_136__dup_933)
                      , .B (modgen_ram_ix167_a_137__dup_932), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2924 (.Y (nx3501), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139__dup_930), .B0 (nx25684), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix25685 (.Y (nx25684), .AN (
                      modgen_ram_ix167_a_138__dup_931), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2925 (.Y (nx2593), .A0 (rd_addr_m_4), .A1 (nx26422)
                          , .B0 (nx26206), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix26423 (.Y (nx26422), .A (nx26254), .B (nx26362), .C (
                     nx26306), .D (nx26414), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix26255 (.Y (nx26254), .A (modgen_ram_ix167_a_176__dup_893)
                     , .B (modgen_ram_ix167_a_178__dup_891), .C (
                     modgen_ram_ix167_a_177__dup_892), .D (
                     modgen_ram_ix167_a_179__dup_890), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix26363 (.Y (nx26362), .A (modgen_ram_ix167_a_184__dup_885)
                     , .B (modgen_ram_ix167_a_186__dup_883), .C (
                     modgen_ram_ix167_a_185__dup_884), .D (
                     modgen_ram_ix167_a_187__dup_882), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix26307 (.Y (nx26306), .A (modgen_ram_ix167_a_180__dup_889)
                     , .B (modgen_ram_ix167_a_182__dup_887), .C (
                     modgen_ram_ix167_a_181__dup_888), .D (
                     modgen_ram_ix167_a_183__dup_886), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix26415 (.Y (nx26414), .A (modgen_ram_ix167_a_188__dup_881)
                     , .B (modgen_ram_ix167_a_190__dup_879), .C (
                     modgen_ram_ix167_a_189__dup_880), .D (
                     modgen_ram_ix167_a_191__dup_878), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26207 (.Y (nx26206), .A0 (rd_addr_m_3), .A1 (nx2605)
                          , .B0 (nx2615), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2926 (.Y (nx2605), .A0 (rd_addr_m_2), .A1 (nx26086), .B0 (
                      nx26038)) ;
    MXT4_X0P5M_A12TS ix26087 (.Y (nx26086), .A (modgen_ram_ix167_a_164__dup_905)
                     , .B (modgen_ram_ix167_a_166__dup_903), .C (
                     modgen_ram_ix167_a_165__dup_904), .D (
                     modgen_ram_ix167_a_167__dup_902), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26039 (.Y (nx26038), .A0 (rd_addr_m_1), .A1 (nx2609)
                          , .B0 (nx2611), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2927 (.Y (nx2609), .A (modgen_ram_ix167_a_160__dup_909)
                      , .B (modgen_ram_ix167_a_161__dup_908), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2928 (.Y (nx2611), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163__dup_906), .B0 (nx26020), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix26021 (.Y (nx26020), .AN (
                      modgen_ram_ix167_a_162__dup_907), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2929 (.Y (nx2615), .A0 (rd_addr_m_2), .A1 (nx26194)
                          , .B0 (nx26146), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix26195 (.Y (nx26194), .A (modgen_ram_ix167_a_172__dup_897)
                     , .B (modgen_ram_ix167_a_174__dup_895), .C (
                     modgen_ram_ix167_a_173__dup_896), .D (
                     modgen_ram_ix167_a_175__dup_894), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix26147 (.Y (nx26146), .A0 (rd_addr_m_1), .A1 (nx3503)
                          , .B0 (nx3504), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2930 (.Y (nx3503), .A (modgen_ram_ix167_a_168__dup_901)
                      , .B (modgen_ram_ix167_a_169__dup_900), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2931 (.Y (nx3504), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171__dup_898), .B0 (nx26128), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix26129 (.Y (nx26128), .AN (
                      modgen_ram_ix167_a_170__dup_899), .B (rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix25543 (.Y (nx25542), .A (rd_addr_7), .B (nx2627)) ;
    AOI21_X0P5M_A12TS ix2932 (.Y (nx2627), .A0 (rd_addr_m_6), .A1 (nx25534), .B0 (
                      nx24646)) ;
    OAI21_X0P5M_A12TS ix25535 (.Y (nx25534), .A0 (rd_addr_m_5), .A1 (nx2631), .B0 (
                      nx2661)) ;
    AOI21_X0P5M_A12TS ix2934 (.Y (nx2631), .A0 (rd_addr_m_4), .A1 (nx25082), .B0 (
                      nx24866)) ;
    MXT4_X0P5M_A12TS ix25083 (.Y (nx25082), .A (nx24914), .B (nx25022), .C (
                     nx24966), .D (nx25074), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix24915 (.Y (nx24914), .A (modgen_ram_ix167_a_80__dup_989)
                     , .B (modgen_ram_ix167_a_82__dup_987), .C (
                     modgen_ram_ix167_a_81__dup_988), .D (
                     modgen_ram_ix167_a_83__dup_986), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25023 (.Y (nx25022), .A (modgen_ram_ix167_a_88__dup_981)
                     , .B (modgen_ram_ix167_a_90__dup_979), .C (
                     modgen_ram_ix167_a_89__dup_980), .D (
                     modgen_ram_ix167_a_91__dup_978), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24967 (.Y (nx24966), .A (modgen_ram_ix167_a_84__dup_985)
                     , .B (modgen_ram_ix167_a_86__dup_983), .C (
                     modgen_ram_ix167_a_85__dup_984), .D (
                     modgen_ram_ix167_a_87__dup_982), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25075 (.Y (nx25074), .A (modgen_ram_ix167_a_92__dup_977)
                     , .B (modgen_ram_ix167_a_94__dup_975), .C (
                     modgen_ram_ix167_a_93__dup_976), .D (
                     modgen_ram_ix167_a_95__dup_974), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24867 (.Y (nx24866), .A0 (rd_addr_m_3), .A1 (nx2639)
                          , .B0 (nx3506), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2935 (.Y (nx2639), .A0 (rd_addr_m_2), .A1 (nx24746), .B0 (
                      nx24698)) ;
    MXT4_X0P5M_A12TS ix24747 (.Y (nx24746), .A (modgen_ram_ix167_a_68__dup_1001)
                     , .B (modgen_ram_ix167_a_70__dup_999), .C (
                     modgen_ram_ix167_a_69__dup_1000), .D (
                     modgen_ram_ix167_a_71__dup_998), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24699 (.Y (nx24698), .A0 (rd_addr_m_1), .A1 (nx2645)
                          , .B0 (nx3505), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2936 (.Y (nx2645), .A (modgen_ram_ix167_a_64__dup_1005)
                      , .B (modgen_ram_ix167_a_65__dup_1004), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2937 (.Y (nx3505), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67__dup_1002), .B0 (nx24680), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix24681 (.Y (nx24680), .AN (
                      modgen_ram_ix167_a_66__dup_1003), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2938 (.Y (nx3506), .A0 (rd_addr_m_2), .A1 (nx24854)
                          , .B0 (nx24806), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix24855 (.Y (nx24854), .A (modgen_ram_ix167_a_76__dup_993)
                     , .B (modgen_ram_ix167_a_78__dup_991), .C (
                     modgen_ram_ix167_a_77__dup_992), .D (
                     modgen_ram_ix167_a_79__dup_990), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24807 (.Y (nx24806), .A0 (rd_addr_m_1), .A1 (nx3507)
                          , .B0 (nx3509), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2940 (.Y (nx3507), .A (modgen_ram_ix167_a_72__dup_997), 
                      .B (modgen_ram_ix167_a_73__dup_996), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2942 (.Y (nx3509), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75__dup_994), .B0 (nx24788), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix24789 (.Y (nx24788), .AN (modgen_ram_ix167_a_74__dup_995
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2943 (.Y (nx2661), .A0 (rd_addr_m_4), .A1 (nx25526)
                          , .B0 (nx25310), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix25527 (.Y (nx25526), .A (nx25358), .B (nx25466), .C (
                     nx25410), .D (nx25518), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix25359 (.Y (nx25358), .A (modgen_ram_ix167_a_112__dup_957)
                     , .B (modgen_ram_ix167_a_114__dup_955), .C (
                     modgen_ram_ix167_a_113__dup_956), .D (
                     modgen_ram_ix167_a_115__dup_954), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25467 (.Y (nx25466), .A (modgen_ram_ix167_a_120__dup_949)
                     , .B (modgen_ram_ix167_a_122__dup_947), .C (
                     modgen_ram_ix167_a_121__dup_948), .D (
                     modgen_ram_ix167_a_123__dup_946), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25411 (.Y (nx25410), .A (modgen_ram_ix167_a_116__dup_953)
                     , .B (modgen_ram_ix167_a_118__dup_951), .C (
                     modgen_ram_ix167_a_117__dup_952), .D (
                     modgen_ram_ix167_a_119__dup_950), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix25519 (.Y (nx25518), .A (modgen_ram_ix167_a_124__dup_945)
                     , .B (modgen_ram_ix167_a_126__dup_943), .C (
                     modgen_ram_ix167_a_125__dup_944), .D (
                     modgen_ram_ix167_a_127__dup_942), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix25311 (.Y (nx25310), .A0 (rd_addr_m_3), .A1 (nx2671)
                          , .B0 (nx3511), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2944 (.Y (nx2671), .A0 (rd_addr_m_2), .A1 (nx25190), .B0 (
                      nx25142)) ;
    MXT4_X0P5M_A12TS ix25191 (.Y (nx25190), .A (modgen_ram_ix167_a_100__dup_969)
                     , .B (modgen_ram_ix167_a_102__dup_967), .C (
                     modgen_ram_ix167_a_101__dup_968), .D (
                     modgen_ram_ix167_a_103__dup_966), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix25143 (.Y (nx25142), .A0 (rd_addr_m_1), .A1 (nx2675)
                          , .B0 (nx3510), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2945 (.Y (nx2675), .A (modgen_ram_ix167_a_96__dup_973), 
                      .B (modgen_ram_ix167_a_97__dup_972), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2946 (.Y (nx3510), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99__dup_970), .B0 (nx25124), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix25125 (.Y (nx25124), .AN (modgen_ram_ix167_a_98__dup_971
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2947 (.Y (nx3511), .A0 (rd_addr_m_2), .A1 (nx25298)
                          , .B0 (nx25250), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix25299 (.Y (nx25298), .A (modgen_ram_ix167_a_108__dup_961)
                     , .B (modgen_ram_ix167_a_110__dup_959), .C (
                     modgen_ram_ix167_a_109__dup_960), .D (
                     modgen_ram_ix167_a_111__dup_958), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix25251 (.Y (nx25250), .A0 (rd_addr_m_1), .A1 (nx2687)
                          , .B0 (nx2689), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2948 (.Y (nx2687), .A (modgen_ram_ix167_a_104__dup_965)
                      , .B (modgen_ram_ix167_a_105__dup_964), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2950 (.Y (nx2689), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107__dup_962), .B0 (nx25232), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix25233 (.Y (nx25232), .AN (
                      modgen_ram_ix167_a_106__dup_963), .B (rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24647 (.Y (nx24646), .A0 (rd_addr_m_5), .A1 (nx2693)
                          , .B0 (nx2723), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2951 (.Y (nx2693), .A0 (rd_addr_m_4), .A1 (nx24190), .B0 (
                      nx23974)) ;
    MXT4_X0P5M_A12TS ix24191 (.Y (nx24190), .A (nx24022), .B (nx24130), .C (
                     nx24074), .D (nx24182), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix24023 (.Y (nx24022), .A (modgen_ram_ix167_a_16__dup_1053)
                     , .B (modgen_ram_ix167_a_18__dup_1051), .C (
                     modgen_ram_ix167_a_17__dup_1052), .D (
                     modgen_ram_ix167_a_19__dup_1050), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24131 (.Y (nx24130), .A (modgen_ram_ix167_a_24__dup_1045)
                     , .B (modgen_ram_ix167_a_26__dup_1043), .C (
                     modgen_ram_ix167_a_25__dup_1044), .D (
                     modgen_ram_ix167_a_27__dup_1042), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24075 (.Y (nx24074), .A (modgen_ram_ix167_a_20__dup_1049)
                     , .B (modgen_ram_ix167_a_22__dup_1047), .C (
                     modgen_ram_ix167_a_21__dup_1048), .D (
                     modgen_ram_ix167_a_23__dup_1046), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24183 (.Y (nx24182), .A (modgen_ram_ix167_a_28__dup_1041)
                     , .B (modgen_ram_ix167_a_30__dup_1039), .C (
                     modgen_ram_ix167_a_29__dup_1040), .D (
                     modgen_ram_ix167_a_31__dup_1038), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23975 (.Y (nx23974), .A0 (rd_addr_m_3), .A1 (nx3512)
                          , .B0 (nx2713), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2952 (.Y (nx3512), .A0 (rd_addr_m_2), .A1 (nx23854), .B0 (
                      nx23806)) ;
    MXT4_X0P5M_A12TS ix23855 (.Y (nx23854), .A (modgen_ram_ix167_a_4__dup_1065)
                     , .B (modgen_ram_ix167_a_6__dup_1063), .C (
                     modgen_ram_ix167_a_5__dup_1064), .D (
                     modgen_ram_ix167_a_7__dup_1062), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23807 (.Y (nx23806), .A0 (rd_addr_m_1), .A1 (nx3513)
                          , .B0 (nx3514), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2953 (.Y (nx3513), .A (modgen_ram_ix167_a_0__dup_1069), 
                      .B (modgen_ram_ix167_a_1__dup_1068), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2954 (.Y (nx3514), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_1066), .B0 (nx23788), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix23789 (.Y (nx23788), .AN (modgen_ram_ix167_a_2__dup_1067
                      ), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2956 (.Y (nx2713), .A0 (rd_addr_m_2), .A1 (nx23962)
                          , .B0 (nx23914), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix23963 (.Y (nx23962), .A (modgen_ram_ix167_a_12__dup_1057)
                     , .B (modgen_ram_ix167_a_14__dup_1055), .C (
                     modgen_ram_ix167_a_13__dup_1056), .D (
                     modgen_ram_ix167_a_15__dup_1054), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix23915 (.Y (nx23914), .A0 (rd_addr_m_1), .A1 (nx3515)
                          , .B0 (nx2720), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2958 (.Y (nx3515), .A (modgen_ram_ix167_a_8__dup_1061), 
                      .B (modgen_ram_ix167_a_9__dup_1060), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2959 (.Y (nx2720), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11__dup_1058), .B0 (nx23896), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix23897 (.Y (nx23896), .AN (
                      modgen_ram_ix167_a_10__dup_1059), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2960 (.Y (nx2723), .A0 (rd_addr_m_4), .A1 (nx24634)
                          , .B0 (nx24418), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix24635 (.Y (nx24634), .A (nx24466), .B (nx24574), .C (
                     nx24518), .D (nx24626), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix24467 (.Y (nx24466), .A (modgen_ram_ix167_a_48__dup_1021)
                     , .B (modgen_ram_ix167_a_50__dup_1019), .C (
                     modgen_ram_ix167_a_49__dup_1020), .D (
                     modgen_ram_ix167_a_51__dup_1018), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24575 (.Y (nx24574), .A (modgen_ram_ix167_a_56__dup_1013)
                     , .B (modgen_ram_ix167_a_58__dup_1011), .C (
                     modgen_ram_ix167_a_57__dup_1012), .D (
                     modgen_ram_ix167_a_59__dup_1010), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24519 (.Y (nx24518), .A (modgen_ram_ix167_a_52__dup_1017)
                     , .B (modgen_ram_ix167_a_54__dup_1015), .C (
                     modgen_ram_ix167_a_53__dup_1016), .D (
                     modgen_ram_ix167_a_55__dup_1014), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix24627 (.Y (nx24626), .A (modgen_ram_ix167_a_60__dup_1009)
                     , .B (modgen_ram_ix167_a_62__dup_1007), .C (
                     modgen_ram_ix167_a_61__dup_1008), .D (
                     modgen_ram_ix167_a_63__dup_1006), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24419 (.Y (nx24418), .A0 (rd_addr_m_3), .A1 (nx2733)
                          , .B0 (nx2742), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2961 (.Y (nx2733), .A0 (rd_addr_m_2), .A1 (nx24298), .B0 (
                      nx24250)) ;
    MXT4_X0P5M_A12TS ix24299 (.Y (nx24298), .A (modgen_ram_ix167_a_36__dup_1033)
                     , .B (modgen_ram_ix167_a_38__dup_1031), .C (
                     modgen_ram_ix167_a_37__dup_1032), .D (
                     modgen_ram_ix167_a_39__dup_1030), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24251 (.Y (nx24250), .A0 (rd_addr_m_1), .A1 (nx3516)
                          , .B0 (nx3517), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2962 (.Y (nx3516), .A (modgen_ram_ix167_a_32__dup_1037)
                      , .B (modgen_ram_ix167_a_33__dup_1036), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2963 (.Y (nx3517), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35__dup_1034), .B0 (nx24232), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix24233 (.Y (nx24232), .AN (
                      modgen_ram_ix167_a_34__dup_1035), .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2964 (.Y (nx2742), .A0 (rd_addr_m_2), .A1 (nx24406)
                          , .B0 (nx24358), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix24407 (.Y (nx24406), .A (modgen_ram_ix167_a_44__dup_1025)
                     , .B (modgen_ram_ix167_a_46__dup_1023), .C (
                     modgen_ram_ix167_a_45__dup_1024), .D (
                     modgen_ram_ix167_a_47__dup_1022), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix24359 (.Y (nx24358), .A0 (rd_addr_m_1), .A1 (nx2747)
                          , .B0 (nx2749), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2966 (.Y (nx2747), .A (modgen_ram_ix167_a_40__dup_1029)
                      , .B (modgen_ram_ix167_a_41__dup_1028), .S0 (rd_addr_m_0)
                      ) ;
    AO21A1AI2_X0P5M_A12TS ix2967 (.Y (nx2749), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43__dup_1026), .B0 (nx24340), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix24341 (.Y (nx24340), .AN (
                      modgen_ram_ix167_a_42__dup_1027), .B (rd_addr_m_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_rd_data_7 (.Q (rd_data_m_7), .CK (wb_clk_i), .D (
                        nx30926), .R (wb_rst_i), .SE (NOT_nx50), .SI (
                        rd_data_m_7)) ;
    MXIT2_X0P5M_A12TS ix30927 (.Y (nx30926), .A (nx2755), .B (nx2757), .S0 (
                      nx1127)) ;
    INV_X0P5B_A12TS ix2968 (.Y (nx2755), .A (wr_data_m_7)) ;
    OA21A1OI2_X0P5M_A12TS ix2969 (.Y (nx2757), .A0 (nx30912), .A1 (nx30022), .B0 (
                          rd_addr_7), .C0 (nx29130)) ;
    OA21A1OI2_X0P5M_A12TS ix30913 (.Y (nx30912), .A0 (rd_addr_m_5), .A1 (nx2760)
                          , .B0 (nx2793), .C0 (nx933)) ;
    AOI21_X0P5M_A12TS ix2970 (.Y (nx2760), .A0 (rd_addr_m_4), .A1 (nx30458), .B0 (
                      nx30242)) ;
    MXT4_X0P5M_A12TS ix30459 (.Y (nx30458), .A (nx30290), .B (nx30398), .C (
                     nx30342), .D (nx30450), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix30291 (.Y (nx30290), .A (modgen_ram_ix167_a_208), .B (
                     modgen_ram_ix167_a_210), .C (modgen_ram_ix167_a_209), .D (
                     modgen_ram_ix167_a_211), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30399 (.Y (nx30398), .A (modgen_ram_ix167_a_216), .B (
                     modgen_ram_ix167_a_218), .C (modgen_ram_ix167_a_217), .D (
                     modgen_ram_ix167_a_219), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30343 (.Y (nx30342), .A (modgen_ram_ix167_a_212), .B (
                     modgen_ram_ix167_a_214), .C (modgen_ram_ix167_a_213), .D (
                     modgen_ram_ix167_a_215), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30451 (.Y (nx30450), .A (modgen_ram_ix167_a_220), .B (
                     modgen_ram_ix167_a_222), .C (modgen_ram_ix167_a_221), .D (
                     modgen_ram_ix167_a_223), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30243 (.Y (nx30242), .A0 (rd_addr_m_3), .A1 (nx2773)
                          , .B0 (nx2783), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2972 (.Y (nx2773), .A0 (rd_addr_m_2), .A1 (nx30122), .B0 (
                      nx30074)) ;
    MXT4_X0P5M_A12TS ix30123 (.Y (nx30122), .A (modgen_ram_ix167_a_196), .B (
                     modgen_ram_ix167_a_198), .C (modgen_ram_ix167_a_197), .D (
                     modgen_ram_ix167_a_199), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30075 (.Y (nx30074), .A0 (rd_addr_m_1), .A1 (nx2777)
                          , .B0 (nx2779), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2973 (.Y (nx2777), .A (modgen_ram_ix167_a_192), .B (
                      modgen_ram_ix167_a_193), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2974 (.Y (nx2779), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_195), .B0 (nx30056), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix30057 (.Y (nx30056), .AN (modgen_ram_ix167_a_194), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2975 (.Y (nx2783), .A0 (rd_addr_m_2), .A1 (nx30230)
                          , .B0 (nx30182), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix30231 (.Y (nx30230), .A (modgen_ram_ix167_a_204), .B (
                     modgen_ram_ix167_a_206), .C (modgen_ram_ix167_a_205), .D (
                     modgen_ram_ix167_a_207), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30183 (.Y (nx30182), .A0 (rd_addr_m_1), .A1 (nx2788)
                          , .B0 (nx2790), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2976 (.Y (nx2788), .A (modgen_ram_ix167_a_200), .B (
                      modgen_ram_ix167_a_201), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2977 (.Y (nx2790), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_203), .B0 (nx30164), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix30165 (.Y (nx30164), .AN (modgen_ram_ix167_a_202), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2978 (.Y (nx2793), .A0 (rd_addr_m_4), .A1 (nx30902)
                          , .B0 (nx30686), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix30903 (.Y (nx30902), .A (nx30734), .B (nx30842), .C (
                     nx30786), .D (nx30894), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix30735 (.Y (nx30734), .A (modgen_ram_ix167_a_240), .B (
                     modgen_ram_ix167_a_242), .C (modgen_ram_ix167_a_241), .D (
                     modgen_ram_ix167_a_243), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30843 (.Y (nx30842), .A (modgen_ram_ix167_a_248), .B (
                     modgen_ram_ix167_a_250), .C (modgen_ram_ix167_a_249), .D (
                     modgen_ram_ix167_a_251), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30787 (.Y (nx30786), .A (modgen_ram_ix167_a_244), .B (
                     modgen_ram_ix167_a_246), .C (modgen_ram_ix167_a_245), .D (
                     modgen_ram_ix167_a_247), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30895 (.Y (nx30894), .A (modgen_ram_ix167_a_252), .B (
                     modgen_ram_ix167_a_254), .C (modgen_ram_ix167_a_253), .D (
                     modgen_ram_ix167_a_255), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30687 (.Y (nx30686), .A0 (rd_addr_m_3), .A1 (nx2803)
                          , .B0 (nx2813), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2979 (.Y (nx2803), .A0 (rd_addr_m_2), .A1 (nx30566), .B0 (
                      nx30518)) ;
    MXT4_X0P5M_A12TS ix30567 (.Y (nx30566), .A (modgen_ram_ix167_a_228), .B (
                     modgen_ram_ix167_a_230), .C (modgen_ram_ix167_a_229), .D (
                     modgen_ram_ix167_a_231), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30519 (.Y (nx30518), .A0 (rd_addr_m_1), .A1 (nx2807)
                          , .B0 (nx2809), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2980 (.Y (nx2807), .A (modgen_ram_ix167_a_224), .B (
                      modgen_ram_ix167_a_225), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2981 (.Y (nx2809), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_227), .B0 (nx30500), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix30501 (.Y (nx30500), .AN (modgen_ram_ix167_a_226), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2982 (.Y (nx2813), .A0 (rd_addr_m_2), .A1 (nx30674)
                          , .B0 (nx30626), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix30675 (.Y (nx30674), .A (modgen_ram_ix167_a_236), .B (
                     modgen_ram_ix167_a_238), .C (modgen_ram_ix167_a_237), .D (
                     modgen_ram_ix167_a_239), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30627 (.Y (nx30626), .A0 (rd_addr_m_1), .A1 (nx2817)
                          , .B0 (nx2819), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2983 (.Y (nx2817), .A (modgen_ram_ix167_a_232), .B (
                      modgen_ram_ix167_a_233), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2984 (.Y (nx2819), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_235), .B0 (nx30608), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix30609 (.Y (nx30608), .AN (modgen_ram_ix167_a_234), .B (
                      rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix30023 (.Y (nx30022), .A0 (rd_addr_m_5), .A1 (nx2825)
                          , .B0 (nx2855), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix2985 (.Y (nx2825), .A0 (rd_addr_m_4), .A1 (nx29566), .B0 (
                      nx29350)) ;
    MXT4_X0P5M_A12TS ix29567 (.Y (nx29566), .A (nx29398), .B (nx29506), .C (
                     nx29450), .D (nx29558), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix29399 (.Y (nx29398), .A (modgen_ram_ix167_a_144), .B (
                     modgen_ram_ix167_a_146), .C (modgen_ram_ix167_a_145), .D (
                     modgen_ram_ix167_a_147), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29507 (.Y (nx29506), .A (modgen_ram_ix167_a_152), .B (
                     modgen_ram_ix167_a_154), .C (modgen_ram_ix167_a_153), .D (
                     modgen_ram_ix167_a_155), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29451 (.Y (nx29450), .A (modgen_ram_ix167_a_148), .B (
                     modgen_ram_ix167_a_150), .C (modgen_ram_ix167_a_149), .D (
                     modgen_ram_ix167_a_151), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29559 (.Y (nx29558), .A (modgen_ram_ix167_a_156), .B (
                     modgen_ram_ix167_a_158), .C (modgen_ram_ix167_a_157), .D (
                     modgen_ram_ix167_a_159), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix29351 (.Y (nx29350), .A0 (rd_addr_m_3), .A1 (nx2833)
                          , .B0 (nx2845), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2986 (.Y (nx2833), .A0 (rd_addr_m_2), .A1 (nx29230), .B0 (
                      nx29182)) ;
    MXT4_X0P5M_A12TS ix29231 (.Y (nx29230), .A (modgen_ram_ix167_a_132), .B (
                     modgen_ram_ix167_a_134), .C (modgen_ram_ix167_a_133), .D (
                     modgen_ram_ix167_a_135), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix29183 (.Y (nx29182), .A0 (rd_addr_m_1), .A1 (nx2839)
                          , .B0 (nx2841), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2987 (.Y (nx2839), .A (modgen_ram_ix167_a_128), .B (
                      modgen_ram_ix167_a_129), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2988 (.Y (nx2841), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_131), .B0 (nx29164), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix29165 (.Y (nx29164), .AN (modgen_ram_ix167_a_130), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2989 (.Y (nx2845), .A0 (rd_addr_m_2), .A1 (nx29338)
                          , .B0 (nx29290), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix29339 (.Y (nx29338), .A (modgen_ram_ix167_a_140), .B (
                     modgen_ram_ix167_a_142), .C (modgen_ram_ix167_a_141), .D (
                     modgen_ram_ix167_a_143), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix29291 (.Y (nx29290), .A0 (rd_addr_m_1), .A1 (nx2849)
                          , .B0 (nx2851), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2990 (.Y (nx2849), .A (modgen_ram_ix167_a_136), .B (
                      modgen_ram_ix167_a_137), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2991 (.Y (nx2851), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_139), .B0 (nx29272), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix29273 (.Y (nx29272), .AN (modgen_ram_ix167_a_138), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2992 (.Y (nx2855), .A0 (rd_addr_m_4), .A1 (nx30010)
                          , .B0 (nx29794), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix30011 (.Y (nx30010), .A (nx29842), .B (nx29950), .C (
                     nx29894), .D (nx30002), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix29843 (.Y (nx29842), .A (modgen_ram_ix167_a_176), .B (
                     modgen_ram_ix167_a_178), .C (modgen_ram_ix167_a_177), .D (
                     modgen_ram_ix167_a_179), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29951 (.Y (nx29950), .A (modgen_ram_ix167_a_184), .B (
                     modgen_ram_ix167_a_186), .C (modgen_ram_ix167_a_185), .D (
                     modgen_ram_ix167_a_187), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29895 (.Y (nx29894), .A (modgen_ram_ix167_a_180), .B (
                     modgen_ram_ix167_a_182), .C (modgen_ram_ix167_a_181), .D (
                     modgen_ram_ix167_a_183), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix30003 (.Y (nx30002), .A (modgen_ram_ix167_a_188), .B (
                     modgen_ram_ix167_a_190), .C (modgen_ram_ix167_a_189), .D (
                     modgen_ram_ix167_a_191), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix29795 (.Y (nx29794), .A0 (rd_addr_m_3), .A1 (nx2865)
                          , .B0 (nx3518), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix2993 (.Y (nx2865), .A0 (rd_addr_m_2), .A1 (nx29674), .B0 (
                      nx29626)) ;
    MXT4_X0P5M_A12TS ix29675 (.Y (nx29674), .A (modgen_ram_ix167_a_164), .B (
                     modgen_ram_ix167_a_166), .C (modgen_ram_ix167_a_165), .D (
                     modgen_ram_ix167_a_167), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix29627 (.Y (nx29626), .A0 (rd_addr_m_1), .A1 (nx2869)
                          , .B0 (nx2871), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2994 (.Y (nx2869), .A (modgen_ram_ix167_a_160), .B (
                      modgen_ram_ix167_a_161), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2995 (.Y (nx2871), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_163), .B0 (nx29608), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix29609 (.Y (nx29608), .AN (modgen_ram_ix167_a_162), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2996 (.Y (nx3518), .A0 (rd_addr_m_2), .A1 (nx29782)
                          , .B0 (nx29734), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix29783 (.Y (nx29782), .A (modgen_ram_ix167_a_172), .B (
                     modgen_ram_ix167_a_174), .C (modgen_ram_ix167_a_173), .D (
                     modgen_ram_ix167_a_175), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix29735 (.Y (nx29734), .A0 (rd_addr_m_1), .A1 (nx2879)
                          , .B0 (nx2881), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix2997 (.Y (nx2879), .A (modgen_ram_ix167_a_168), .B (
                      modgen_ram_ix167_a_169), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix2998 (.Y (nx2881), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_171), .B0 (nx29716), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix29717 (.Y (nx29716), .AN (modgen_ram_ix167_a_170), .B (
                      rd_addr_m_0)) ;
    NOR2_X0P5A_A12TS ix29131 (.Y (nx29130), .A (rd_addr_7), .B (nx2887)) ;
    AOI21_X0P5M_A12TS ix2999 (.Y (nx2887), .A0 (rd_addr_m_6), .A1 (nx29122), .B0 (
                      nx28234)) ;
    OAI21_X0P5M_A12TS ix29123 (.Y (nx29122), .A0 (rd_addr_m_5), .A1 (nx2890), .B0 (
                      nx2921)) ;
    AOI21_X0P5M_A12TS ix3000 (.Y (nx2890), .A0 (rd_addr_m_4), .A1 (nx28670), .B0 (
                      nx28454)) ;
    MXT4_X0P5M_A12TS ix28671 (.Y (nx28670), .A (nx28502), .B (nx28610), .C (
                     nx28554), .D (nx28662), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix28503 (.Y (nx28502), .A (modgen_ram_ix167_a_80), .B (
                     modgen_ram_ix167_a_82), .C (modgen_ram_ix167_a_81), .D (
                     modgen_ram_ix167_a_83), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix28611 (.Y (nx28610), .A (modgen_ram_ix167_a_88), .B (
                     modgen_ram_ix167_a_90), .C (modgen_ram_ix167_a_89), .D (
                     modgen_ram_ix167_a_91), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix28555 (.Y (nx28554), .A (modgen_ram_ix167_a_84), .B (
                     modgen_ram_ix167_a_86), .C (modgen_ram_ix167_a_85), .D (
                     modgen_ram_ix167_a_87), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix28663 (.Y (nx28662), .A (modgen_ram_ix167_a_92), .B (
                     modgen_ram_ix167_a_94), .C (modgen_ram_ix167_a_93), .D (
                     modgen_ram_ix167_a_95), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix28455 (.Y (nx28454), .A0 (rd_addr_m_3), .A1 (nx2901)
                          , .B0 (nx2911), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix3001 (.Y (nx2901), .A0 (rd_addr_m_2), .A1 (nx28334), .B0 (
                      nx28286)) ;
    MXT4_X0P5M_A12TS ix28335 (.Y (nx28334), .A (modgen_ram_ix167_a_68), .B (
                     modgen_ram_ix167_a_70), .C (modgen_ram_ix167_a_69), .D (
                     modgen_ram_ix167_a_71), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix28287 (.Y (nx28286), .A0 (rd_addr_m_1), .A1 (nx2905)
                          , .B0 (nx2907), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3002 (.Y (nx2905), .A (modgen_ram_ix167_a_64), .B (
                      modgen_ram_ix167_a_65), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3004 (.Y (nx2907), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_67), .B0 (nx28268), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix28269 (.Y (nx28268), .AN (modgen_ram_ix167_a_66), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3005 (.Y (nx2911), .A0 (rd_addr_m_2), .A1 (nx28442)
                          , .B0 (nx28394), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix28443 (.Y (nx28442), .A (modgen_ram_ix167_a_76), .B (
                     modgen_ram_ix167_a_78), .C (modgen_ram_ix167_a_77), .D (
                     modgen_ram_ix167_a_79), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix28395 (.Y (nx28394), .A0 (rd_addr_m_1), .A1 (nx2915)
                          , .B0 (nx2917), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3006 (.Y (nx2915), .A (modgen_ram_ix167_a_72), .B (
                      modgen_ram_ix167_a_73), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3007 (.Y (nx2917), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_75), .B0 (nx28376), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix28377 (.Y (nx28376), .AN (modgen_ram_ix167_a_74), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3008 (.Y (nx2921), .A0 (rd_addr_m_4), .A1 (nx29114)
                          , .B0 (nx28898), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix29115 (.Y (nx29114), .A (nx28946), .B (nx29054), .C (
                     nx28998), .D (nx29106), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix28947 (.Y (nx28946), .A (modgen_ram_ix167_a_112), .B (
                     modgen_ram_ix167_a_114), .C (modgen_ram_ix167_a_113), .D (
                     modgen_ram_ix167_a_115), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29055 (.Y (nx29054), .A (modgen_ram_ix167_a_120), .B (
                     modgen_ram_ix167_a_122), .C (modgen_ram_ix167_a_121), .D (
                     modgen_ram_ix167_a_123), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix28999 (.Y (nx28998), .A (modgen_ram_ix167_a_116), .B (
                     modgen_ram_ix167_a_118), .C (modgen_ram_ix167_a_117), .D (
                     modgen_ram_ix167_a_119), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    MXT4_X0P5M_A12TS ix29107 (.Y (nx29106), .A (modgen_ram_ix167_a_124), .B (
                     modgen_ram_ix167_a_126), .C (modgen_ram_ix167_a_125), .D (
                     modgen_ram_ix167_a_127), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix28899 (.Y (nx28898), .A0 (rd_addr_m_3), .A1 (nx2931)
                          , .B0 (nx2941), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix3009 (.Y (nx2931), .A0 (rd_addr_m_2), .A1 (nx28778), .B0 (
                      nx28730)) ;
    MXT4_X0P5M_A12TS ix28779 (.Y (nx28778), .A (modgen_ram_ix167_a_100), .B (
                     modgen_ram_ix167_a_102), .C (modgen_ram_ix167_a_101), .D (
                     modgen_ram_ix167_a_103), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix28731 (.Y (nx28730), .A0 (rd_addr_m_1), .A1 (nx2935)
                          , .B0 (nx2937), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3010 (.Y (nx2935), .A (modgen_ram_ix167_a_96), .B (
                      modgen_ram_ix167_a_97), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3012 (.Y (nx2937), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_99), .B0 (nx28712), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix28713 (.Y (nx28712), .AN (modgen_ram_ix167_a_98), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3013 (.Y (nx2941), .A0 (rd_addr_m_2), .A1 (nx28886)
                          , .B0 (nx28838), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix28887 (.Y (nx28886), .A (modgen_ram_ix167_a_108), .B (
                     modgen_ram_ix167_a_110), .C (modgen_ram_ix167_a_109), .D (
                     modgen_ram_ix167_a_111), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix28839 (.Y (nx28838), .A0 (rd_addr_m_1), .A1 (nx2947)
                          , .B0 (nx2949), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3014 (.Y (nx2947), .A (modgen_ram_ix167_a_104), .B (
                      modgen_ram_ix167_a_105), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3015 (.Y (nx2949), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_107), .B0 (nx28820), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix28821 (.Y (nx28820), .AN (modgen_ram_ix167_a_106), .B (
                      rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix28235 (.Y (nx28234), .A0 (rd_addr_m_5), .A1 (nx2955)
                          , .B0 (nx2991), .C0 (rd_addr_m_6)) ;
    AOI21_X0P5M_A12TS ix3016 (.Y (nx2955), .A0 (rd_addr_m_4), .A1 (nx27778), .B0 (
                      nx27562)) ;
    MXT4_X0P5M_A12TS ix27779 (.Y (nx27778), .A (nx27610), .B (nx27718), .C (
                     nx27662), .D (nx27770), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix27611 (.Y (nx27610), .A (modgen_ram_ix167_a_16), .B (
                     modgen_ram_ix167_a_18), .C (modgen_ram_ix167_a_17), .D (
                     modgen_ram_ix167_a_19), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix27719 (.Y (nx27718), .A (modgen_ram_ix167_a_24), .B (
                     modgen_ram_ix167_a_26), .C (modgen_ram_ix167_a_25), .D (
                     modgen_ram_ix167_a_27), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix27663 (.Y (nx27662), .A (modgen_ram_ix167_a_20), .B (
                     modgen_ram_ix167_a_22), .C (modgen_ram_ix167_a_21), .D (
                     modgen_ram_ix167_a_23), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix27771 (.Y (nx27770), .A (modgen_ram_ix167_a_28), .B (
                     modgen_ram_ix167_a_30), .C (modgen_ram_ix167_a_29), .D (
                     modgen_ram_ix167_a_31), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix27563 (.Y (nx27562), .A0 (rd_addr_m_3), .A1 (nx2969)
                          , .B0 (nx2981), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix3018 (.Y (nx2969), .A0 (rd_addr_m_2), .A1 (nx27442), .B0 (
                      nx27394)) ;
    MXT4_X0P5M_A12TS ix27443 (.Y (nx27442), .A (modgen_ram_ix167_a_4__dup_807), 
                     .B (modgen_ram_ix167_a_6__dup_805), .C (
                     modgen_ram_ix167_a_5__dup_806), .D (
                     modgen_ram_ix167_a_7__dup_804), .S0 (rd_addr_m_1), .S1 (
                     rd_addr_m_0)) ;
    OA21A1OI2_X0P5M_A12TS ix27395 (.Y (nx27394), .A0 (rd_addr_m_1), .A1 (nx2975)
                          , .B0 (nx2977), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3019 (.Y (nx2975), .A (modgen_ram_ix167_a_0__dup_811), .B (
                      modgen_ram_ix167_a_1__dup_810), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3020 (.Y (nx2977), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_3__dup_808), .B0 (nx27376), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix27377 (.Y (nx27376), .AN (modgen_ram_ix167_a_2__dup_809)
                      , .B (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3021 (.Y (nx2981), .A0 (rd_addr_m_2), .A1 (nx27550)
                          , .B0 (nx27502), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix27551 (.Y (nx27550), .A (modgen_ram_ix167_a_12), .B (
                     modgen_ram_ix167_a_14), .C (modgen_ram_ix167_a_13), .D (
                     modgen_ram_ix167_a_15), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix27503 (.Y (nx27502), .A0 (rd_addr_m_1), .A1 (nx2985)
                          , .B0 (nx2987), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3022 (.Y (nx2985), .A (modgen_ram_ix167_a_8), .B (
                      modgen_ram_ix167_a_9), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3024 (.Y (nx2987), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_11), .B0 (nx27484), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix27485 (.Y (nx27484), .AN (modgen_ram_ix167_a_10), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3025 (.Y (nx2991), .A0 (rd_addr_m_4), .A1 (nx28222)
                          , .B0 (nx28006), .C0 (rd_addr_m_5)) ;
    MXT4_X0P5M_A12TS ix28223 (.Y (nx28222), .A (nx28054), .B (nx28162), .C (
                     nx28106), .D (nx28214), .S0 (rd_addr_m_3), .S1 (rd_addr_m_2
                     )) ;
    MXT4_X0P5M_A12TS ix28055 (.Y (nx28054), .A (modgen_ram_ix167_a_48), .B (
                     modgen_ram_ix167_a_50), .C (modgen_ram_ix167_a_49), .D (
                     modgen_ram_ix167_a_51), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix28163 (.Y (nx28162), .A (modgen_ram_ix167_a_56), .B (
                     modgen_ram_ix167_a_58), .C (modgen_ram_ix167_a_57), .D (
                     modgen_ram_ix167_a_59), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix28107 (.Y (nx28106), .A (modgen_ram_ix167_a_52), .B (
                     modgen_ram_ix167_a_54), .C (modgen_ram_ix167_a_53), .D (
                     modgen_ram_ix167_a_55), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    MXT4_X0P5M_A12TS ix28215 (.Y (nx28214), .A (modgen_ram_ix167_a_60), .B (
                     modgen_ram_ix167_a_62), .C (modgen_ram_ix167_a_61), .D (
                     modgen_ram_ix167_a_63), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix28007 (.Y (nx28006), .A0 (rd_addr_m_3), .A1 (nx3001)
                          , .B0 (nx3011), .C0 (rd_addr_m_4)) ;
    AOI21_X0P5M_A12TS ix3026 (.Y (nx3001), .A0 (rd_addr_m_2), .A1 (nx27886), .B0 (
                      nx27838)) ;
    MXT4_X0P5M_A12TS ix27887 (.Y (nx27886), .A (modgen_ram_ix167_a_36), .B (
                     modgen_ram_ix167_a_38), .C (modgen_ram_ix167_a_37), .D (
                     modgen_ram_ix167_a_39), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix27839 (.Y (nx27838), .A0 (rd_addr_m_1), .A1 (nx3005)
                          , .B0 (nx3007), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3027 (.Y (nx3005), .A (modgen_ram_ix167_a_32), .B (
                      modgen_ram_ix167_a_33), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3028 (.Y (nx3007), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_35), .B0 (nx27820), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix27821 (.Y (nx27820), .AN (modgen_ram_ix167_a_34), .B (
                      rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3030 (.Y (nx3011), .A0 (rd_addr_m_2), .A1 (nx27994)
                          , .B0 (nx27946), .C0 (rd_addr_m_3)) ;
    MXT4_X0P5M_A12TS ix27995 (.Y (nx27994), .A (modgen_ram_ix167_a_44), .B (
                     modgen_ram_ix167_a_46), .C (modgen_ram_ix167_a_45), .D (
                     modgen_ram_ix167_a_47), .S0 (rd_addr_m_1), .S1 (rd_addr_m_0
                     )) ;
    OA21A1OI2_X0P5M_A12TS ix27947 (.Y (nx27946), .A0 (rd_addr_m_1), .A1 (nx3015)
                          , .B0 (nx3017), .C0 (rd_addr_m_2)) ;
    MXIT2_X0P5M_A12TS ix3031 (.Y (nx3015), .A (modgen_ram_ix167_a_40), .B (
                      modgen_ram_ix167_a_41), .S0 (rd_addr_m_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3032 (.Y (nx3017), .A0 (rd_addr_m_0), .A1 (
                          modgen_ram_ix167_a_43), .B0 (nx27928), .C0 (
                          rd_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix27929 (.Y (nx27928), .AN (modgen_ram_ix167_a_42), .B (
                      rd_addr_m_0)) ;
    NOR2B_X0P7M_A12TS ix3033 (.Y (nx3287), .AN (wr_addr_m_1), .B (wr_addr_m_0)
                      ) ;
    NOR2B_X0P7M_A12TS ix444 (.Y (nx443), .AN (wr_addr_m_0), .B (wr_addr_m_1)) ;
    NOR2B_X0P7M_A12TS ix3034 (.Y (nx3289), .AN (wr_addr_m_3), .B (wr_addr_m_2)
                      ) ;
    NOR2B_X0P7M_A12TS ix3036 (.Y (nx3290), .AN (wr_addr_m_2), .B (wr_addr_m_3)
                      ) ;
    NOR2B_X0P7M_A12TS ix504 (.Y (nx503), .AN (wr_addr_m_5), .B (wr_addr_m_4)) ;
    NOR2B_X0P7M_A12TS ix530 (.Y (nx529), .AN (wr_addr_m_4), .B (wr_addr_m_5)) ;
    NOR2B_X0P7M_A12TS ix3037 (.Y (nx3291), .AN (wr_addr_7), .B (wr_addr_m_6)) ;
    NOR2B_X0P7M_A12TS ix674 (.Y (nx673), .AN (wr_addr_m_6), .B (wr_addr_7)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix297 (.Q (modgen_ram_ix167_a_255), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5764)
                         , .SI (modgen_ram_ix167_a_255), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix301 (.Q (modgen_ram_ix167_a_254), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5746)
                         , .SI (modgen_ram_ix167_a_254), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix305 (.Q (modgen_ram_ix167_a_253), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5724)
                         , .SI (modgen_ram_ix167_a_253), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix309 (.Q (modgen_ram_ix167_a_252), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5706)
                         , .SI (modgen_ram_ix167_a_252), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix313 (.Q (modgen_ram_ix167_a_251), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5680)
                         , .SI (modgen_ram_ix167_a_251), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix317 (.Q (modgen_ram_ix167_a_250), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5662)
                         , .SI (modgen_ram_ix167_a_250), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix321 (.Q (modgen_ram_ix167_a_249), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5640)
                         , .SI (modgen_ram_ix167_a_249), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix325 (.Q (modgen_ram_ix167_a_248), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5622)
                         , .SI (modgen_ram_ix167_a_248), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix329 (.Q (modgen_ram_ix167_a_247), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5592)
                         , .SI (modgen_ram_ix167_a_247), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix333 (.Q (modgen_ram_ix167_a_246), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5574)
                         , .SI (modgen_ram_ix167_a_246), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix337 (.Q (modgen_ram_ix167_a_245), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5552)
                         , .SI (modgen_ram_ix167_a_245), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix341 (.Q (modgen_ram_ix167_a_244), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5534)
                         , .SI (modgen_ram_ix167_a_244), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix345 (.Q (modgen_ram_ix167_a_243), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5508)
                         , .SI (modgen_ram_ix167_a_243), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix349 (.Q (modgen_ram_ix167_a_242), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5490)
                         , .SI (modgen_ram_ix167_a_242), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix353 (.Q (modgen_ram_ix167_a_241), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5468)
                         , .SI (modgen_ram_ix167_a_241), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix357 (.Q (modgen_ram_ix167_a_240), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5450)
                         , .SI (modgen_ram_ix167_a_240), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix361 (.Q (modgen_ram_ix167_a_239), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5414)
                         , .SI (modgen_ram_ix167_a_239), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix365 (.Q (modgen_ram_ix167_a_238), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5396)
                         , .SI (modgen_ram_ix167_a_238), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix369 (.Q (modgen_ram_ix167_a_237), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5374)
                         , .SI (modgen_ram_ix167_a_237), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix373 (.Q (modgen_ram_ix167_a_236), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5356)
                         , .SI (modgen_ram_ix167_a_236), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix377 (.Q (modgen_ram_ix167_a_235), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5330)
                         , .SI (modgen_ram_ix167_a_235), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix381 (.Q (modgen_ram_ix167_a_234), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5312)
                         , .SI (modgen_ram_ix167_a_234), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix385 (.Q (modgen_ram_ix167_a_233), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5290)
                         , .SI (modgen_ram_ix167_a_233), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix389 (.Q (modgen_ram_ix167_a_232), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5272)
                         , .SI (modgen_ram_ix167_a_232), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix393 (.Q (modgen_ram_ix167_a_231), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5242)
                         , .SI (modgen_ram_ix167_a_231), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix397 (.Q (modgen_ram_ix167_a_230), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5224)
                         , .SI (modgen_ram_ix167_a_230), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix401 (.Q (modgen_ram_ix167_a_229), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5202)
                         , .SI (modgen_ram_ix167_a_229), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix405 (.Q (modgen_ram_ix167_a_228), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5184)
                         , .SI (modgen_ram_ix167_a_228), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix409 (.Q (modgen_ram_ix167_a_227), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5158)
                         , .SI (modgen_ram_ix167_a_227), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix413 (.Q (modgen_ram_ix167_a_226), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5140)
                         , .SI (modgen_ram_ix167_a_226), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix417 (.Q (modgen_ram_ix167_a_225), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5118)
                         , .SI (modgen_ram_ix167_a_225), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix421 (.Q (modgen_ram_ix167_a_224), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5100)
                         , .SI (modgen_ram_ix167_a_224), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix425 (.Q (modgen_ram_ix167_a_223), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5060)
                         , .SI (modgen_ram_ix167_a_223), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix429 (.Q (modgen_ram_ix167_a_222), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5042)
                         , .SI (modgen_ram_ix167_a_222), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix433 (.Q (modgen_ram_ix167_a_221), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5020)
                         , .SI (modgen_ram_ix167_a_221), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix437 (.Q (modgen_ram_ix167_a_220), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx5002)
                         , .SI (modgen_ram_ix167_a_220), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix441 (.Q (modgen_ram_ix167_a_219), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4976)
                         , .SI (modgen_ram_ix167_a_219), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix445 (.Q (modgen_ram_ix167_a_218), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4958)
                         , .SI (modgen_ram_ix167_a_218), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix449 (.Q (modgen_ram_ix167_a_217), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4936)
                         , .SI (modgen_ram_ix167_a_217), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix453 (.Q (modgen_ram_ix167_a_216), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4918)
                         , .SI (modgen_ram_ix167_a_216), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix457 (.Q (modgen_ram_ix167_a_215), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4888)
                         , .SI (modgen_ram_ix167_a_215), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix461 (.Q (modgen_ram_ix167_a_214), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4870)
                         , .SI (modgen_ram_ix167_a_214), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix465 (.Q (modgen_ram_ix167_a_213), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4848)
                         , .SI (modgen_ram_ix167_a_213), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix469 (.Q (modgen_ram_ix167_a_212), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4830)
                         , .SI (modgen_ram_ix167_a_212), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix473 (.Q (modgen_ram_ix167_a_211), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4804)
                         , .SI (modgen_ram_ix167_a_211), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix477 (.Q (modgen_ram_ix167_a_210), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4786)
                         , .SI (modgen_ram_ix167_a_210), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix481 (.Q (modgen_ram_ix167_a_209), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4764)
                         , .SI (modgen_ram_ix167_a_209), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix485 (.Q (modgen_ram_ix167_a_208), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4746)
                         , .SI (modgen_ram_ix167_a_208), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix489 (.Q (modgen_ram_ix167_a_207), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4710)
                         , .SI (modgen_ram_ix167_a_207), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix493 (.Q (modgen_ram_ix167_a_206), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4692)
                         , .SI (modgen_ram_ix167_a_206), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix497 (.Q (modgen_ram_ix167_a_205), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4670)
                         , .SI (modgen_ram_ix167_a_205), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix501 (.Q (modgen_ram_ix167_a_204), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4652)
                         , .SI (modgen_ram_ix167_a_204), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix505 (.Q (modgen_ram_ix167_a_203), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4626)
                         , .SI (modgen_ram_ix167_a_203), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix509 (.Q (modgen_ram_ix167_a_202), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4608)
                         , .SI (modgen_ram_ix167_a_202), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix513 (.Q (modgen_ram_ix167_a_201), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4586)
                         , .SI (modgen_ram_ix167_a_201), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix517 (.Q (modgen_ram_ix167_a_200), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4568)
                         , .SI (modgen_ram_ix167_a_200), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix521 (.Q (modgen_ram_ix167_a_199), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4538)
                         , .SI (modgen_ram_ix167_a_199), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix525 (.Q (modgen_ram_ix167_a_198), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4520)
                         , .SI (modgen_ram_ix167_a_198), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix529 (.Q (modgen_ram_ix167_a_197), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4498)
                         , .SI (modgen_ram_ix167_a_197), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix533 (.Q (modgen_ram_ix167_a_196), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4480)
                         , .SI (modgen_ram_ix167_a_196), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix537 (.Q (modgen_ram_ix167_a_195), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4454)
                         , .SI (modgen_ram_ix167_a_195), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix541 (.Q (modgen_ram_ix167_a_194), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4436)
                         , .SI (modgen_ram_ix167_a_194), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix545 (.Q (modgen_ram_ix167_a_193), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4414)
                         , .SI (modgen_ram_ix167_a_193), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix549 (.Q (modgen_ram_ix167_a_192), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4396)
                         , .SI (modgen_ram_ix167_a_192), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix553 (.Q (modgen_ram_ix167_a_191), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4346)
                         , .SI (modgen_ram_ix167_a_191), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix557 (.Q (modgen_ram_ix167_a_190), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4328)
                         , .SI (modgen_ram_ix167_a_190), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix561 (.Q (modgen_ram_ix167_a_189), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4306)
                         , .SI (modgen_ram_ix167_a_189), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix565 (.Q (modgen_ram_ix167_a_188), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4288)
                         , .SI (modgen_ram_ix167_a_188), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix569 (.Q (modgen_ram_ix167_a_187), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4262)
                         , .SI (modgen_ram_ix167_a_187), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix573 (.Q (modgen_ram_ix167_a_186), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4244)
                         , .SI (modgen_ram_ix167_a_186), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix577 (.Q (modgen_ram_ix167_a_185), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4222)
                         , .SI (modgen_ram_ix167_a_185), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix581 (.Q (modgen_ram_ix167_a_184), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4204)
                         , .SI (modgen_ram_ix167_a_184), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix585 (.Q (modgen_ram_ix167_a_183), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4174)
                         , .SI (modgen_ram_ix167_a_183), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix589 (.Q (modgen_ram_ix167_a_182), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4156)
                         , .SI (modgen_ram_ix167_a_182), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix593 (.Q (modgen_ram_ix167_a_181), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4134)
                         , .SI (modgen_ram_ix167_a_181), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix597 (.Q (modgen_ram_ix167_a_180), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4116)
                         , .SI (modgen_ram_ix167_a_180), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix601 (.Q (modgen_ram_ix167_a_179), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4090)
                         , .SI (modgen_ram_ix167_a_179), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix605 (.Q (modgen_ram_ix167_a_178), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4072)
                         , .SI (modgen_ram_ix167_a_178), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix609 (.Q (modgen_ram_ix167_a_177), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4050)
                         , .SI (modgen_ram_ix167_a_177), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix613 (.Q (modgen_ram_ix167_a_176), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx4032)
                         , .SI (modgen_ram_ix167_a_176), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix617 (.Q (modgen_ram_ix167_a_175), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3996)
                         , .SI (modgen_ram_ix167_a_175), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix621 (.Q (modgen_ram_ix167_a_174), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3978)
                         , .SI (modgen_ram_ix167_a_174), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix625 (.Q (modgen_ram_ix167_a_173), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3956)
                         , .SI (modgen_ram_ix167_a_173), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix629 (.Q (modgen_ram_ix167_a_172), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3938)
                         , .SI (modgen_ram_ix167_a_172), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix633 (.Q (modgen_ram_ix167_a_171), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3912)
                         , .SI (modgen_ram_ix167_a_171), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix637 (.Q (modgen_ram_ix167_a_170), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3894)
                         , .SI (modgen_ram_ix167_a_170), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix641 (.Q (modgen_ram_ix167_a_169), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3872)
                         , .SI (modgen_ram_ix167_a_169), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix645 (.Q (modgen_ram_ix167_a_168), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3854)
                         , .SI (modgen_ram_ix167_a_168), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix649 (.Q (modgen_ram_ix167_a_167), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3824)
                         , .SI (modgen_ram_ix167_a_167), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix653 (.Q (modgen_ram_ix167_a_166), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3806)
                         , .SI (modgen_ram_ix167_a_166), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix657 (.Q (modgen_ram_ix167_a_165), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3784)
                         , .SI (modgen_ram_ix167_a_165), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix661 (.Q (modgen_ram_ix167_a_164), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3766)
                         , .SI (modgen_ram_ix167_a_164), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix665 (.Q (modgen_ram_ix167_a_163), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3740)
                         , .SI (modgen_ram_ix167_a_163), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix669 (.Q (modgen_ram_ix167_a_162), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3722)
                         , .SI (modgen_ram_ix167_a_162), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix673 (.Q (modgen_ram_ix167_a_161), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3700)
                         , .SI (modgen_ram_ix167_a_161), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix677 (.Q (modgen_ram_ix167_a_160), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3682)
                         , .SI (modgen_ram_ix167_a_160), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix681 (.Q (modgen_ram_ix167_a_159), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3642)
                         , .SI (modgen_ram_ix167_a_159), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix685 (.Q (modgen_ram_ix167_a_158), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3624)
                         , .SI (modgen_ram_ix167_a_158), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix689 (.Q (modgen_ram_ix167_a_157), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3602)
                         , .SI (modgen_ram_ix167_a_157), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix693 (.Q (modgen_ram_ix167_a_156), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3584)
                         , .SI (modgen_ram_ix167_a_156), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix697 (.Q (modgen_ram_ix167_a_155), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3558)
                         , .SI (modgen_ram_ix167_a_155), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix701 (.Q (modgen_ram_ix167_a_154), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3540)
                         , .SI (modgen_ram_ix167_a_154), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix705 (.Q (modgen_ram_ix167_a_153), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3518)
                         , .SI (modgen_ram_ix167_a_153), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix709 (.Q (modgen_ram_ix167_a_152), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3500)
                         , .SI (modgen_ram_ix167_a_152), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix713 (.Q (modgen_ram_ix167_a_151), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3470)
                         , .SI (modgen_ram_ix167_a_151), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix717 (.Q (modgen_ram_ix167_a_150), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3452)
                         , .SI (modgen_ram_ix167_a_150), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix721 (.Q (modgen_ram_ix167_a_149), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3430)
                         , .SI (modgen_ram_ix167_a_149), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix725 (.Q (modgen_ram_ix167_a_148), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3412)
                         , .SI (modgen_ram_ix167_a_148), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix729 (.Q (modgen_ram_ix167_a_147), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3386)
                         , .SI (modgen_ram_ix167_a_147), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix733 (.Q (modgen_ram_ix167_a_146), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3368)
                         , .SI (modgen_ram_ix167_a_146), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix737 (.Q (modgen_ram_ix167_a_145), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3346)
                         , .SI (modgen_ram_ix167_a_145), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix741 (.Q (modgen_ram_ix167_a_144), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3328)
                         , .SI (modgen_ram_ix167_a_144), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix745 (.Q (modgen_ram_ix167_a_143), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3292)
                         , .SI (modgen_ram_ix167_a_143), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix749 (.Q (modgen_ram_ix167_a_142), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3274)
                         , .SI (modgen_ram_ix167_a_142), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix753 (.Q (modgen_ram_ix167_a_141), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3252)
                         , .SI (modgen_ram_ix167_a_141), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix757 (.Q (modgen_ram_ix167_a_140), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3234)
                         , .SI (modgen_ram_ix167_a_140), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix761 (.Q (modgen_ram_ix167_a_139), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3208)
                         , .SI (modgen_ram_ix167_a_139), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix765 (.Q (modgen_ram_ix167_a_138), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3190)
                         , .SI (modgen_ram_ix167_a_138), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix769 (.Q (modgen_ram_ix167_a_137), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3168)
                         , .SI (modgen_ram_ix167_a_137), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix773 (.Q (modgen_ram_ix167_a_136), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3150)
                         , .SI (modgen_ram_ix167_a_136), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix777 (.Q (modgen_ram_ix167_a_135), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3120)
                         , .SI (modgen_ram_ix167_a_135), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix781 (.Q (modgen_ram_ix167_a_134), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3102)
                         , .SI (modgen_ram_ix167_a_134), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix785 (.Q (modgen_ram_ix167_a_133), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3080)
                         , .SI (modgen_ram_ix167_a_133), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix789 (.Q (modgen_ram_ix167_a_132), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3062)
                         , .SI (modgen_ram_ix167_a_132), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix793 (.Q (modgen_ram_ix167_a_131), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3036)
                         , .SI (modgen_ram_ix167_a_131), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix797 (.Q (modgen_ram_ix167_a_130), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx3018)
                         , .SI (modgen_ram_ix167_a_130), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix801 (.Q (modgen_ram_ix167_a_129), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2996)
                         , .SI (modgen_ram_ix167_a_129), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix805 (.Q (modgen_ram_ix167_a_128), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2978)
                         , .SI (modgen_ram_ix167_a_128), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix809 (.Q (modgen_ram_ix167_a_127), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2926)
                         , .SI (modgen_ram_ix167_a_127), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix813 (.Q (modgen_ram_ix167_a_126), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2908)
                         , .SI (modgen_ram_ix167_a_126), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix817 (.Q (modgen_ram_ix167_a_125), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2886)
                         , .SI (modgen_ram_ix167_a_125), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix821 (.Q (modgen_ram_ix167_a_124), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2868)
                         , .SI (modgen_ram_ix167_a_124), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix825 (.Q (modgen_ram_ix167_a_123), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2842)
                         , .SI (modgen_ram_ix167_a_123), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix829 (.Q (modgen_ram_ix167_a_122), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2824)
                         , .SI (modgen_ram_ix167_a_122), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix833 (.Q (modgen_ram_ix167_a_121), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2802)
                         , .SI (modgen_ram_ix167_a_121), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix837 (.Q (modgen_ram_ix167_a_120), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2784)
                         , .SI (modgen_ram_ix167_a_120), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix841 (.Q (modgen_ram_ix167_a_119), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2754)
                         , .SI (modgen_ram_ix167_a_119), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix845 (.Q (modgen_ram_ix167_a_118), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2736)
                         , .SI (modgen_ram_ix167_a_118), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix849 (.Q (modgen_ram_ix167_a_117), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2714)
                         , .SI (modgen_ram_ix167_a_117), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix853 (.Q (modgen_ram_ix167_a_116), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2696)
                         , .SI (modgen_ram_ix167_a_116), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix857 (.Q (modgen_ram_ix167_a_115), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2670)
                         , .SI (modgen_ram_ix167_a_115), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix861 (.Q (modgen_ram_ix167_a_114), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2652)
                         , .SI (modgen_ram_ix167_a_114), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix865 (.Q (modgen_ram_ix167_a_113), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2630)
                         , .SI (modgen_ram_ix167_a_113), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix869 (.Q (modgen_ram_ix167_a_112), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2612)
                         , .SI (modgen_ram_ix167_a_112), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix873 (.Q (modgen_ram_ix167_a_111), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2576)
                         , .SI (modgen_ram_ix167_a_111), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix877 (.Q (modgen_ram_ix167_a_110), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2558)
                         , .SI (modgen_ram_ix167_a_110), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix881 (.Q (modgen_ram_ix167_a_109), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2536)
                         , .SI (modgen_ram_ix167_a_109), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix885 (.Q (modgen_ram_ix167_a_108), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2518)
                         , .SI (modgen_ram_ix167_a_108), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix889 (.Q (modgen_ram_ix167_a_107), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2492)
                         , .SI (modgen_ram_ix167_a_107), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix893 (.Q (modgen_ram_ix167_a_106), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2474)
                         , .SI (modgen_ram_ix167_a_106), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix897 (.Q (modgen_ram_ix167_a_105), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2452)
                         , .SI (modgen_ram_ix167_a_105), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix901 (.Q (modgen_ram_ix167_a_104), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2434)
                         , .SI (modgen_ram_ix167_a_104), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix905 (.Q (modgen_ram_ix167_a_103), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2404)
                         , .SI (modgen_ram_ix167_a_103), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix909 (.Q (modgen_ram_ix167_a_102), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2386)
                         , .SI (modgen_ram_ix167_a_102), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix913 (.Q (modgen_ram_ix167_a_101), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2364)
                         , .SI (modgen_ram_ix167_a_101), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix917 (.Q (modgen_ram_ix167_a_100), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2346)
                         , .SI (modgen_ram_ix167_a_100), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix921 (.Q (modgen_ram_ix167_a_99), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2320)
                         , .SI (modgen_ram_ix167_a_99), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix925 (.Q (modgen_ram_ix167_a_98), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2302)
                         , .SI (modgen_ram_ix167_a_98), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix929 (.Q (modgen_ram_ix167_a_97), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2280)
                         , .SI (modgen_ram_ix167_a_97), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix933 (.Q (modgen_ram_ix167_a_96), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2262)
                         , .SI (modgen_ram_ix167_a_96), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix937 (.Q (modgen_ram_ix167_a_95), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2222)
                         , .SI (modgen_ram_ix167_a_95), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix941 (.Q (modgen_ram_ix167_a_94), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2204)
                         , .SI (modgen_ram_ix167_a_94), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix945 (.Q (modgen_ram_ix167_a_93), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2182)
                         , .SI (modgen_ram_ix167_a_93), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix949 (.Q (modgen_ram_ix167_a_92), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2164)
                         , .SI (modgen_ram_ix167_a_92), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix953 (.Q (modgen_ram_ix167_a_91), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2138)
                         , .SI (modgen_ram_ix167_a_91), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix957 (.Q (modgen_ram_ix167_a_90), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2120)
                         , .SI (modgen_ram_ix167_a_90), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix961 (.Q (modgen_ram_ix167_a_89), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2098)
                         , .SI (modgen_ram_ix167_a_89), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix965 (.Q (modgen_ram_ix167_a_88), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2080)
                         , .SI (modgen_ram_ix167_a_88), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix969 (.Q (modgen_ram_ix167_a_87), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2050)
                         , .SI (modgen_ram_ix167_a_87), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix973 (.Q (modgen_ram_ix167_a_86), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2032)
                         , .SI (modgen_ram_ix167_a_86), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix977 (.Q (modgen_ram_ix167_a_85), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx2010)
                         , .SI (modgen_ram_ix167_a_85), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix981 (.Q (modgen_ram_ix167_a_84), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1992)
                         , .SI (modgen_ram_ix167_a_84), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix985 (.Q (modgen_ram_ix167_a_83), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1966)
                         , .SI (modgen_ram_ix167_a_83), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix989 (.Q (modgen_ram_ix167_a_82), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1948)
                         , .SI (modgen_ram_ix167_a_82), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix993 (.Q (modgen_ram_ix167_a_81), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1926)
                         , .SI (modgen_ram_ix167_a_81), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix997 (.Q (modgen_ram_ix167_a_80), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1908)
                         , .SI (modgen_ram_ix167_a_80), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1001 (.Q (modgen_ram_ix167_a_79), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1872)
                         , .SI (modgen_ram_ix167_a_79), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1005 (.Q (modgen_ram_ix167_a_78), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1854)
                         , .SI (modgen_ram_ix167_a_78), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1009 (.Q (modgen_ram_ix167_a_77), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1832)
                         , .SI (modgen_ram_ix167_a_77), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1013 (.Q (modgen_ram_ix167_a_76), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1814)
                         , .SI (modgen_ram_ix167_a_76), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1017 (.Q (modgen_ram_ix167_a_75), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1788)
                         , .SI (modgen_ram_ix167_a_75), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1021 (.Q (modgen_ram_ix167_a_74), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1770)
                         , .SI (modgen_ram_ix167_a_74), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1025 (.Q (modgen_ram_ix167_a_73), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1748)
                         , .SI (modgen_ram_ix167_a_73), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1029 (.Q (modgen_ram_ix167_a_72), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1730)
                         , .SI (modgen_ram_ix167_a_72), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1033 (.Q (modgen_ram_ix167_a_71), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1700)
                         , .SI (modgen_ram_ix167_a_71), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1037 (.Q (modgen_ram_ix167_a_70), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1682)
                         , .SI (modgen_ram_ix167_a_70), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1041 (.Q (modgen_ram_ix167_a_69), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1660)
                         , .SI (modgen_ram_ix167_a_69), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1045 (.Q (modgen_ram_ix167_a_68), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1642)
                         , .SI (modgen_ram_ix167_a_68), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1049 (.Q (modgen_ram_ix167_a_67), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1616)
                         , .SI (modgen_ram_ix167_a_67), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1053 (.Q (modgen_ram_ix167_a_66), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1598)
                         , .SI (modgen_ram_ix167_a_66), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1057 (.Q (modgen_ram_ix167_a_65), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1576)
                         , .SI (modgen_ram_ix167_a_65), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1061 (.Q (modgen_ram_ix167_a_64), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1558)
                         , .SI (modgen_ram_ix167_a_64), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1065 (.Q (modgen_ram_ix167_a_63), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1510)
                         , .SI (modgen_ram_ix167_a_63), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1069 (.Q (modgen_ram_ix167_a_62), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1492)
                         , .SI (modgen_ram_ix167_a_62), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1073 (.Q (modgen_ram_ix167_a_61), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1470)
                         , .SI (modgen_ram_ix167_a_61), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1077 (.Q (modgen_ram_ix167_a_60), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1452)
                         , .SI (modgen_ram_ix167_a_60), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1081 (.Q (modgen_ram_ix167_a_59), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1426)
                         , .SI (modgen_ram_ix167_a_59), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1085 (.Q (modgen_ram_ix167_a_58), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1408)
                         , .SI (modgen_ram_ix167_a_58), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1089 (.Q (modgen_ram_ix167_a_57), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1386)
                         , .SI (modgen_ram_ix167_a_57), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1093 (.Q (modgen_ram_ix167_a_56), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1368)
                         , .SI (modgen_ram_ix167_a_56), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1097 (.Q (modgen_ram_ix167_a_55), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1338)
                         , .SI (modgen_ram_ix167_a_55), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1101 (.Q (modgen_ram_ix167_a_54), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1320)
                         , .SI (modgen_ram_ix167_a_54), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1105 (.Q (modgen_ram_ix167_a_53), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1298)
                         , .SI (modgen_ram_ix167_a_53), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1109 (.Q (modgen_ram_ix167_a_52), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1280)
                         , .SI (modgen_ram_ix167_a_52), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1113 (.Q (modgen_ram_ix167_a_51), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1254)
                         , .SI (modgen_ram_ix167_a_51), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1117 (.Q (modgen_ram_ix167_a_50), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1236)
                         , .SI (modgen_ram_ix167_a_50), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1121 (.Q (modgen_ram_ix167_a_49), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1214)
                         , .SI (modgen_ram_ix167_a_49), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1125 (.Q (modgen_ram_ix167_a_48), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1196)
                         , .SI (modgen_ram_ix167_a_48), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1129 (.Q (modgen_ram_ix167_a_47), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1154)
                         , .SI (modgen_ram_ix167_a_47), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1133 (.Q (modgen_ram_ix167_a_46), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1136)
                         , .SI (modgen_ram_ix167_a_46), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1137 (.Q (modgen_ram_ix167_a_45), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1114)
                         , .SI (modgen_ram_ix167_a_45), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1141 (.Q (modgen_ram_ix167_a_44), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1096)
                         , .SI (modgen_ram_ix167_a_44), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1145 (.Q (modgen_ram_ix167_a_43), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1070)
                         , .SI (modgen_ram_ix167_a_43), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1149 (.Q (modgen_ram_ix167_a_42), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1052)
                         , .SI (modgen_ram_ix167_a_42), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1153 (.Q (modgen_ram_ix167_a_41), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1030)
                         , .SI (modgen_ram_ix167_a_41), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1157 (.Q (modgen_ram_ix167_a_40), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx1012)
                         , .SI (modgen_ram_ix167_a_40), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1161 (.Q (modgen_ram_ix167_a_39), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx982), 
                         .SI (modgen_ram_ix167_a_39), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1165 (.Q (modgen_ram_ix167_a_38), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx964), 
                         .SI (modgen_ram_ix167_a_38), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1169 (.Q (modgen_ram_ix167_a_37), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx942), 
                         .SI (modgen_ram_ix167_a_37), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1173 (.Q (modgen_ram_ix167_a_36), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx924), 
                         .SI (modgen_ram_ix167_a_36), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1177 (.Q (modgen_ram_ix167_a_35), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx898), 
                         .SI (modgen_ram_ix167_a_35), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1181 (.Q (modgen_ram_ix167_a_34), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx880), 
                         .SI (modgen_ram_ix167_a_34), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1185 (.Q (modgen_ram_ix167_a_33), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx858), 
                         .SI (modgen_ram_ix167_a_33), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1189 (.Q (modgen_ram_ix167_a_32), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx840), 
                         .SI (modgen_ram_ix167_a_32), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1193 (.Q (modgen_ram_ix167_a_31), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx796), 
                         .SI (modgen_ram_ix167_a_31), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1197 (.Q (modgen_ram_ix167_a_30), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx778), 
                         .SI (modgen_ram_ix167_a_30), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1201 (.Q (modgen_ram_ix167_a_29), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx756), 
                         .SI (modgen_ram_ix167_a_29), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1205 (.Q (modgen_ram_ix167_a_28), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx738), 
                         .SI (modgen_ram_ix167_a_28), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1209 (.Q (modgen_ram_ix167_a_27), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx712), 
                         .SI (modgen_ram_ix167_a_27), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1213 (.Q (modgen_ram_ix167_a_26), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx694), 
                         .SI (modgen_ram_ix167_a_26), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1217 (.Q (modgen_ram_ix167_a_25), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx672), 
                         .SI (modgen_ram_ix167_a_25), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1221 (.Q (modgen_ram_ix167_a_24), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx654), 
                         .SI (modgen_ram_ix167_a_24), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1225 (.Q (modgen_ram_ix167_a_23), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx624), 
                         .SI (modgen_ram_ix167_a_23), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1229 (.Q (modgen_ram_ix167_a_22), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx606), 
                         .SI (modgen_ram_ix167_a_22), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1233 (.Q (modgen_ram_ix167_a_21), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx584), 
                         .SI (modgen_ram_ix167_a_21), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1237 (.Q (modgen_ram_ix167_a_20), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx566), 
                         .SI (modgen_ram_ix167_a_20), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1241 (.Q (modgen_ram_ix167_a_19), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx540), 
                         .SI (modgen_ram_ix167_a_19), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1245 (.Q (modgen_ram_ix167_a_18), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx522), 
                         .SI (modgen_ram_ix167_a_18), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1249 (.Q (modgen_ram_ix167_a_17), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx500), 
                         .SI (modgen_ram_ix167_a_17), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1253 (.Q (modgen_ram_ix167_a_16), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx482), 
                         .SI (modgen_ram_ix167_a_16), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1257 (.Q (modgen_ram_ix167_a_15), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx442), 
                         .SI (modgen_ram_ix167_a_15), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1261 (.Q (modgen_ram_ix167_a_14), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx422), 
                         .SI (modgen_ram_ix167_a_14), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1265 (.Q (modgen_ram_ix167_a_13), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx398), 
                         .SI (modgen_ram_ix167_a_13), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1269 (.Q (modgen_ram_ix167_a_12), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx378), 
                         .SI (modgen_ram_ix167_a_12), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1273 (.Q (modgen_ram_ix167_a_11), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx344), 
                         .SI (modgen_ram_ix167_a_11), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1277 (.Q (modgen_ram_ix167_a_10), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx324), 
                         .SI (modgen_ram_ix167_a_10), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1281 (.Q (modgen_ram_ix167_a_9), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx340), 
                         .SI (modgen_ram_ix167_a_9), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1285 (.Q (modgen_ram_ix167_a_8), .CK (
                         wb_clk_i), .D (nx28509), .R (nx3204), .SE (NOT_nx280), 
                         .SI (modgen_ram_ix167_a_8), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1289 (.Q (
                         modgen_ram_ix167_a_7__dup_804), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_804), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1293 (.Q (
                         modgen_ram_ix167_a_6__dup_805), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_805), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1297 (.Q (
                         modgen_ram_ix167_a_5__dup_806), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_806), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1301 (.Q (
                         modgen_ram_ix167_a_4__dup_807), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_807), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1305 (.Q (
                         modgen_ram_ix167_a_3__dup_808), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_808), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1309 (.Q (
                         modgen_ram_ix167_a_2__dup_809), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_809), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1313 (.Q (
                         modgen_ram_ix167_a_1__dup_810), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_810), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1317 (.Q (
                         modgen_ram_ix167_a_0__dup_811), .CK (wb_clk_i), .D (
                         nx28509), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_811), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1324 (.Q (
                         modgen_ram_ix167_a_255__dup_814), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_814), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1328 (.Q (
                         modgen_ram_ix167_a_254__dup_815), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_815), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1332 (.Q (
                         modgen_ram_ix167_a_253__dup_816), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_816), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1336 (.Q (
                         modgen_ram_ix167_a_252__dup_817), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_817), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1340 (.Q (
                         modgen_ram_ix167_a_251__dup_818), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_818), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1344 (.Q (
                         modgen_ram_ix167_a_250__dup_819), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_819), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1348 (.Q (
                         modgen_ram_ix167_a_249__dup_820), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_820), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1352 (.Q (
                         modgen_ram_ix167_a_248__dup_821), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_821), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1356 (.Q (
                         modgen_ram_ix167_a_247__dup_822), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_822), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1360 (.Q (
                         modgen_ram_ix167_a_246__dup_823), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_823), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1364 (.Q (
                         modgen_ram_ix167_a_245__dup_824), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_824), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1368 (.Q (
                         modgen_ram_ix167_a_244__dup_825), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_825), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1372 (.Q (
                         modgen_ram_ix167_a_243__dup_826), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_826), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1376 (.Q (
                         modgen_ram_ix167_a_242__dup_827), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_827), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1380 (.Q (
                         modgen_ram_ix167_a_241__dup_828), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_828), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1384 (.Q (
                         modgen_ram_ix167_a_240__dup_829), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_829), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1388 (.Q (
                         modgen_ram_ix167_a_239__dup_830), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_830), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1392 (.Q (
                         modgen_ram_ix167_a_238__dup_831), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_831), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1396 (.Q (
                         modgen_ram_ix167_a_237__dup_832), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_832), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1400 (.Q (
                         modgen_ram_ix167_a_236__dup_833), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_833), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1404 (.Q (
                         modgen_ram_ix167_a_235__dup_834), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_834), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1408 (.Q (
                         modgen_ram_ix167_a_234__dup_835), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_835), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1412 (.Q (
                         modgen_ram_ix167_a_233__dup_836), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_836), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1416 (.Q (
                         modgen_ram_ix167_a_232__dup_837), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_837), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1420 (.Q (
                         modgen_ram_ix167_a_231__dup_838), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_838), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1424 (.Q (
                         modgen_ram_ix167_a_230__dup_839), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_839), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1428 (.Q (
                         modgen_ram_ix167_a_229__dup_840), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_840), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1432 (.Q (
                         modgen_ram_ix167_a_228__dup_841), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_841), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1436 (.Q (
                         modgen_ram_ix167_a_227__dup_842), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_842), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1440 (.Q (
                         modgen_ram_ix167_a_226__dup_843), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_843), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1444 (.Q (
                         modgen_ram_ix167_a_225__dup_844), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_844), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1448 (.Q (
                         modgen_ram_ix167_a_224__dup_845), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_845), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1452 (.Q (
                         modgen_ram_ix167_a_223__dup_846), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_846), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1456 (.Q (
                         modgen_ram_ix167_a_222__dup_847), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_847), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1460 (.Q (
                         modgen_ram_ix167_a_221__dup_848), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_848), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1464 (.Q (
                         modgen_ram_ix167_a_220__dup_849), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_849), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1468 (.Q (
                         modgen_ram_ix167_a_219__dup_850), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_850), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1472 (.Q (
                         modgen_ram_ix167_a_218__dup_851), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_851), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1476 (.Q (
                         modgen_ram_ix167_a_217__dup_852), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_852), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1480 (.Q (
                         modgen_ram_ix167_a_216__dup_853), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_853), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1484 (.Q (
                         modgen_ram_ix167_a_215__dup_854), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_854), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1488 (.Q (
                         modgen_ram_ix167_a_214__dup_855), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_855), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1492 (.Q (
                         modgen_ram_ix167_a_213__dup_856), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_856), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1496 (.Q (
                         modgen_ram_ix167_a_212__dup_857), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_857), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1500 (.Q (
                         modgen_ram_ix167_a_211__dup_858), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_858), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1504 (.Q (
                         modgen_ram_ix167_a_210__dup_859), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_859), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1508 (.Q (
                         modgen_ram_ix167_a_209__dup_860), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_860), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1512 (.Q (
                         modgen_ram_ix167_a_208__dup_861), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_861), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1516 (.Q (
                         modgen_ram_ix167_a_207__dup_862), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_862), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1520 (.Q (
                         modgen_ram_ix167_a_206__dup_863), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_863), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1524 (.Q (
                         modgen_ram_ix167_a_205__dup_864), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_864), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1528 (.Q (
                         modgen_ram_ix167_a_204__dup_865), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_865), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1532 (.Q (
                         modgen_ram_ix167_a_203__dup_866), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_866), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1536 (.Q (
                         modgen_ram_ix167_a_202__dup_867), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_867), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1540 (.Q (
                         modgen_ram_ix167_a_201__dup_868), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_868), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1544 (.Q (
                         modgen_ram_ix167_a_200__dup_869), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_869), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1548 (.Q (
                         modgen_ram_ix167_a_199__dup_870), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_870), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1552 (.Q (
                         modgen_ram_ix167_a_198__dup_871), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_871), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1556 (.Q (
                         modgen_ram_ix167_a_197__dup_872), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_872), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1560 (.Q (
                         modgen_ram_ix167_a_196__dup_873), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_873), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1564 (.Q (
                         modgen_ram_ix167_a_195__dup_874), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_874), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1568 (.Q (
                         modgen_ram_ix167_a_194__dup_875), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_875), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1572 (.Q (
                         modgen_ram_ix167_a_193__dup_876), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_876), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1576 (.Q (
                         modgen_ram_ix167_a_192__dup_877), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_877), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1580 (.Q (
                         modgen_ram_ix167_a_191__dup_878), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_878), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1584 (.Q (
                         modgen_ram_ix167_a_190__dup_879), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_879), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1588 (.Q (
                         modgen_ram_ix167_a_189__dup_880), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_880), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1592 (.Q (
                         modgen_ram_ix167_a_188__dup_881), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_881), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1596 (.Q (
                         modgen_ram_ix167_a_187__dup_882), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_882), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1600 (.Q (
                         modgen_ram_ix167_a_186__dup_883), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_883), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1604 (.Q (
                         modgen_ram_ix167_a_185__dup_884), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_884), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1608 (.Q (
                         modgen_ram_ix167_a_184__dup_885), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_885), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1612 (.Q (
                         modgen_ram_ix167_a_183__dup_886), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_886), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1616 (.Q (
                         modgen_ram_ix167_a_182__dup_887), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_887), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1620 (.Q (
                         modgen_ram_ix167_a_181__dup_888), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_888), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1624 (.Q (
                         modgen_ram_ix167_a_180__dup_889), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_889), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1628 (.Q (
                         modgen_ram_ix167_a_179__dup_890), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_890), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1632 (.Q (
                         modgen_ram_ix167_a_178__dup_891), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_891), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1636 (.Q (
                         modgen_ram_ix167_a_177__dup_892), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_892), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1640 (.Q (
                         modgen_ram_ix167_a_176__dup_893), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_893), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1644 (.Q (
                         modgen_ram_ix167_a_175__dup_894), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_894), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1648 (.Q (
                         modgen_ram_ix167_a_174__dup_895), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_895), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1652 (.Q (
                         modgen_ram_ix167_a_173__dup_896), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_896), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1656 (.Q (
                         modgen_ram_ix167_a_172__dup_897), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_897), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1660 (.Q (
                         modgen_ram_ix167_a_171__dup_898), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_898), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1664 (.Q (
                         modgen_ram_ix167_a_170__dup_899), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_899), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1668 (.Q (
                         modgen_ram_ix167_a_169__dup_900), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_900), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1672 (.Q (
                         modgen_ram_ix167_a_168__dup_901), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_901), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1676 (.Q (
                         modgen_ram_ix167_a_167__dup_902), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_902), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1680 (.Q (
                         modgen_ram_ix167_a_166__dup_903), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_903), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1684 (.Q (
                         modgen_ram_ix167_a_165__dup_904), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_904), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1688 (.Q (
                         modgen_ram_ix167_a_164__dup_905), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_905), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1692 (.Q (
                         modgen_ram_ix167_a_163__dup_906), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_906), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1696 (.Q (
                         modgen_ram_ix167_a_162__dup_907), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_907), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1700 (.Q (
                         modgen_ram_ix167_a_161__dup_908), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_908), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1704 (.Q (
                         modgen_ram_ix167_a_160__dup_909), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_909), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1708 (.Q (
                         modgen_ram_ix167_a_159__dup_910), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_910), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1712 (.Q (
                         modgen_ram_ix167_a_158__dup_911), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_911), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1716 (.Q (
                         modgen_ram_ix167_a_157__dup_912), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_912), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1720 (.Q (
                         modgen_ram_ix167_a_156__dup_913), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_913), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1724 (.Q (
                         modgen_ram_ix167_a_155__dup_914), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_914), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1728 (.Q (
                         modgen_ram_ix167_a_154__dup_915), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_915), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1732 (.Q (
                         modgen_ram_ix167_a_153__dup_916), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_916), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1736 (.Q (
                         modgen_ram_ix167_a_152__dup_917), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_917), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1740 (.Q (
                         modgen_ram_ix167_a_151__dup_918), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_918), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1744 (.Q (
                         modgen_ram_ix167_a_150__dup_919), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_919), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1748 (.Q (
                         modgen_ram_ix167_a_149__dup_920), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_920), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1752 (.Q (
                         modgen_ram_ix167_a_148__dup_921), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_921), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1756 (.Q (
                         modgen_ram_ix167_a_147__dup_922), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_922), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1760 (.Q (
                         modgen_ram_ix167_a_146__dup_923), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_923), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1764 (.Q (
                         modgen_ram_ix167_a_145__dup_924), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_924), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1768 (.Q (
                         modgen_ram_ix167_a_144__dup_925), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_925), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1772 (.Q (
                         modgen_ram_ix167_a_143__dup_926), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_926), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1776 (.Q (
                         modgen_ram_ix167_a_142__dup_927), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_927), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1780 (.Q (
                         modgen_ram_ix167_a_141__dup_928), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_928), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1784 (.Q (
                         modgen_ram_ix167_a_140__dup_929), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_929), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1788 (.Q (
                         modgen_ram_ix167_a_139__dup_930), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_930), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1792 (.Q (
                         modgen_ram_ix167_a_138__dup_931), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_931), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1796 (.Q (
                         modgen_ram_ix167_a_137__dup_932), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_932), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1800 (.Q (
                         modgen_ram_ix167_a_136__dup_933), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_933), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1804 (.Q (
                         modgen_ram_ix167_a_135__dup_934), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_934), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1808 (.Q (
                         modgen_ram_ix167_a_134__dup_935), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_935), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1812 (.Q (
                         modgen_ram_ix167_a_133__dup_936), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_936), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1816 (.Q (
                         modgen_ram_ix167_a_132__dup_937), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_937), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1820 (.Q (
                         modgen_ram_ix167_a_131__dup_938), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_938), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1824 (.Q (
                         modgen_ram_ix167_a_130__dup_939), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_939), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1828 (.Q (
                         modgen_ram_ix167_a_129__dup_940), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_940), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1832 (.Q (
                         modgen_ram_ix167_a_128__dup_941), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_941), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1836 (.Q (
                         modgen_ram_ix167_a_127__dup_942), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_942), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1840 (.Q (
                         modgen_ram_ix167_a_126__dup_943), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_943), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1844 (.Q (
                         modgen_ram_ix167_a_125__dup_944), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_944), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1848 (.Q (
                         modgen_ram_ix167_a_124__dup_945), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_945), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1852 (.Q (
                         modgen_ram_ix167_a_123__dup_946), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_946), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1856 (.Q (
                         modgen_ram_ix167_a_122__dup_947), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_947), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1860 (.Q (
                         modgen_ram_ix167_a_121__dup_948), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_948), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1864 (.Q (
                         modgen_ram_ix167_a_120__dup_949), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_949), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1868 (.Q (
                         modgen_ram_ix167_a_119__dup_950), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_950), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1872 (.Q (
                         modgen_ram_ix167_a_118__dup_951), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_951), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1876 (.Q (
                         modgen_ram_ix167_a_117__dup_952), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_952), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1880 (.Q (
                         modgen_ram_ix167_a_116__dup_953), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_953), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1884 (.Q (
                         modgen_ram_ix167_a_115__dup_954), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_954), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1888 (.Q (
                         modgen_ram_ix167_a_114__dup_955), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_955), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1892 (.Q (
                         modgen_ram_ix167_a_113__dup_956), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_956), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1896 (.Q (
                         modgen_ram_ix167_a_112__dup_957), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_957), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1900 (.Q (
                         modgen_ram_ix167_a_111__dup_958), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_958), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1904 (.Q (
                         modgen_ram_ix167_a_110__dup_959), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_959), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1908 (.Q (
                         modgen_ram_ix167_a_109__dup_960), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_960), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1912 (.Q (
                         modgen_ram_ix167_a_108__dup_961), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_961), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1916 (.Q (
                         modgen_ram_ix167_a_107__dup_962), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_962), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1920 (.Q (
                         modgen_ram_ix167_a_106__dup_963), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_963), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1924 (.Q (
                         modgen_ram_ix167_a_105__dup_964), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_964), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1928 (.Q (
                         modgen_ram_ix167_a_104__dup_965), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_965), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1932 (.Q (
                         modgen_ram_ix167_a_103__dup_966), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_966), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1936 (.Q (
                         modgen_ram_ix167_a_102__dup_967), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_967), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1940 (.Q (
                         modgen_ram_ix167_a_101__dup_968), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_968), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1944 (.Q (
                         modgen_ram_ix167_a_100__dup_969), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_969), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1948 (.Q (
                         modgen_ram_ix167_a_99__dup_970), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_970), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1952 (.Q (
                         modgen_ram_ix167_a_98__dup_971), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_971), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1956 (.Q (
                         modgen_ram_ix167_a_97__dup_972), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_972), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1960 (.Q (
                         modgen_ram_ix167_a_96__dup_973), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_973), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1964 (.Q (
                         modgen_ram_ix167_a_95__dup_974), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_974), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1968 (.Q (
                         modgen_ram_ix167_a_94__dup_975), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_975), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1972 (.Q (
                         modgen_ram_ix167_a_93__dup_976), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_976), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1976 (.Q (
                         modgen_ram_ix167_a_92__dup_977), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_977), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1980 (.Q (
                         modgen_ram_ix167_a_91__dup_978), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_978), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1984 (.Q (
                         modgen_ram_ix167_a_90__dup_979), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_979), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1988 (.Q (
                         modgen_ram_ix167_a_89__dup_980), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_980), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1992 (.Q (
                         modgen_ram_ix167_a_88__dup_981), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_981), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix1996 (.Q (
                         modgen_ram_ix167_a_87__dup_982), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_982), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2000 (.Q (
                         modgen_ram_ix167_a_86__dup_983), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_983), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2004 (.Q (
                         modgen_ram_ix167_a_85__dup_984), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_984), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2008 (.Q (
                         modgen_ram_ix167_a_84__dup_985), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_985), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2012 (.Q (
                         modgen_ram_ix167_a_83__dup_986), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_986), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2016 (.Q (
                         modgen_ram_ix167_a_82__dup_987), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_987), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2020 (.Q (
                         modgen_ram_ix167_a_81__dup_988), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_988), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2024 (.Q (
                         modgen_ram_ix167_a_80__dup_989), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_989), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2028 (.Q (
                         modgen_ram_ix167_a_79__dup_990), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_990), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2032 (.Q (
                         modgen_ram_ix167_a_78__dup_991), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_991), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2036 (.Q (
                         modgen_ram_ix167_a_77__dup_992), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_992), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2040 (.Q (
                         modgen_ram_ix167_a_76__dup_993), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_993), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2044 (.Q (
                         modgen_ram_ix167_a_75__dup_994), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_994), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2048 (.Q (
                         modgen_ram_ix167_a_74__dup_995), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_995), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2052 (.Q (
                         modgen_ram_ix167_a_73__dup_996), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_996), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2056 (.Q (
                         modgen_ram_ix167_a_72__dup_997), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_997), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2060 (.Q (
                         modgen_ram_ix167_a_71__dup_998), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_998), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2064 (.Q (
                         modgen_ram_ix167_a_70__dup_999), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_999), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2068 (.Q (
                         modgen_ram_ix167_a_69__dup_1000), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_1000), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2072 (.Q (
                         modgen_ram_ix167_a_68__dup_1001), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_1001), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2076 (.Q (
                         modgen_ram_ix167_a_67__dup_1002), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_1002), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2080 (.Q (
                         modgen_ram_ix167_a_66__dup_1003), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_1003), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2084 (.Q (
                         modgen_ram_ix167_a_65__dup_1004), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_1004), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2088 (.Q (
                         modgen_ram_ix167_a_64__dup_1005), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_1005), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2092 (.Q (
                         modgen_ram_ix167_a_63__dup_1006), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_1006), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2096 (.Q (
                         modgen_ram_ix167_a_62__dup_1007), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_1007), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2100 (.Q (
                         modgen_ram_ix167_a_61__dup_1008), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_1008), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2104 (.Q (
                         modgen_ram_ix167_a_60__dup_1009), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_1009), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2108 (.Q (
                         modgen_ram_ix167_a_59__dup_1010), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_1010), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2112 (.Q (
                         modgen_ram_ix167_a_58__dup_1011), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_1011), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2116 (.Q (
                         modgen_ram_ix167_a_57__dup_1012), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_1012), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2120 (.Q (
                         modgen_ram_ix167_a_56__dup_1013), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_1013), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2124 (.Q (
                         modgen_ram_ix167_a_55__dup_1014), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_1014), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2128 (.Q (
                         modgen_ram_ix167_a_54__dup_1015), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_1015), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2132 (.Q (
                         modgen_ram_ix167_a_53__dup_1016), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_1016), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2136 (.Q (
                         modgen_ram_ix167_a_52__dup_1017), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_1017), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2140 (.Q (
                         modgen_ram_ix167_a_51__dup_1018), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_1018), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2144 (.Q (
                         modgen_ram_ix167_a_50__dup_1019), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_1019), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2148 (.Q (
                         modgen_ram_ix167_a_49__dup_1020), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_1020), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2152 (.Q (
                         modgen_ram_ix167_a_48__dup_1021), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_1021), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2156 (.Q (
                         modgen_ram_ix167_a_47__dup_1022), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_1022), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2160 (.Q (
                         modgen_ram_ix167_a_46__dup_1023), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_1023), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2164 (.Q (
                         modgen_ram_ix167_a_45__dup_1024), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_1024), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2168 (.Q (
                         modgen_ram_ix167_a_44__dup_1025), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_1025), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2172 (.Q (
                         modgen_ram_ix167_a_43__dup_1026), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_1026), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2176 (.Q (
                         modgen_ram_ix167_a_42__dup_1027), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_1027), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2180 (.Q (
                         modgen_ram_ix167_a_41__dup_1028), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_1028), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2184 (.Q (
                         modgen_ram_ix167_a_40__dup_1029), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_1029), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2188 (.Q (
                         modgen_ram_ix167_a_39__dup_1030), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_1030), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2192 (.Q (
                         modgen_ram_ix167_a_38__dup_1031), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_1031), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2196 (.Q (
                         modgen_ram_ix167_a_37__dup_1032), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_1032), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2200 (.Q (
                         modgen_ram_ix167_a_36__dup_1033), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_1033), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2204 (.Q (
                         modgen_ram_ix167_a_35__dup_1034), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_1034), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2208 (.Q (
                         modgen_ram_ix167_a_34__dup_1035), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_1035), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2212 (.Q (
                         modgen_ram_ix167_a_33__dup_1036), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_1036), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2216 (.Q (
                         modgen_ram_ix167_a_32__dup_1037), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_1037), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2220 (.Q (
                         modgen_ram_ix167_a_31__dup_1038), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_1038), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2224 (.Q (
                         modgen_ram_ix167_a_30__dup_1039), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_1039), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2228 (.Q (
                         modgen_ram_ix167_a_29__dup_1040), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_1040), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2232 (.Q (
                         modgen_ram_ix167_a_28__dup_1041), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_1041), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2236 (.Q (
                         modgen_ram_ix167_a_27__dup_1042), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_1042), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2240 (.Q (
                         modgen_ram_ix167_a_26__dup_1043), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_1043), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2244 (.Q (
                         modgen_ram_ix167_a_25__dup_1044), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_1044), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2248 (.Q (
                         modgen_ram_ix167_a_24__dup_1045), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_1045), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2252 (.Q (
                         modgen_ram_ix167_a_23__dup_1046), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_1046), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2256 (.Q (
                         modgen_ram_ix167_a_22__dup_1047), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_1047), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2260 (.Q (
                         modgen_ram_ix167_a_21__dup_1048), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_1048), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2264 (.Q (
                         modgen_ram_ix167_a_20__dup_1049), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_1049), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2268 (.Q (
                         modgen_ram_ix167_a_19__dup_1050), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_1050), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2272 (.Q (
                         modgen_ram_ix167_a_18__dup_1051), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_1051), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2276 (.Q (
                         modgen_ram_ix167_a_17__dup_1052), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_1052), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2280 (.Q (
                         modgen_ram_ix167_a_16__dup_1053), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_1053), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2284 (.Q (
                         modgen_ram_ix167_a_15__dup_1054), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_1054), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2288 (.Q (
                         modgen_ram_ix167_a_14__dup_1055), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_1055), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2292 (.Q (
                         modgen_ram_ix167_a_13__dup_1056), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_1056), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2296 (.Q (
                         modgen_ram_ix167_a_12__dup_1057), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_1057), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2300 (.Q (
                         modgen_ram_ix167_a_11__dup_1058), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_1058), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2304 (.Q (
                         modgen_ram_ix167_a_10__dup_1059), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_1059), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2308 (.Q (
                         modgen_ram_ix167_a_9__dup_1060), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_1060), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2312 (.Q (
                         modgen_ram_ix167_a_8__dup_1061), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_1061), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2316 (.Q (
                         modgen_ram_ix167_a_7__dup_1062), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_1062), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2320 (.Q (
                         modgen_ram_ix167_a_6__dup_1063), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_1063), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2324 (.Q (
                         modgen_ram_ix167_a_5__dup_1064), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_1064), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2328 (.Q (
                         modgen_ram_ix167_a_4__dup_1065), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_1065), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2332 (.Q (
                         modgen_ram_ix167_a_3__dup_1066), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_1066), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2336 (.Q (
                         modgen_ram_ix167_a_2__dup_1067), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_1067), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2340 (.Q (
                         modgen_ram_ix167_a_1__dup_1068), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_1068), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2344 (.Q (
                         modgen_ram_ix167_a_0__dup_1069), .CK (wb_clk_i), .D (
                         nx28511), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_1069), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2349 (.Q (
                         modgen_ram_ix167_a_255__dup_1078), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_1078), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2353 (.Q (
                         modgen_ram_ix167_a_254__dup_1079), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_1079), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2357 (.Q (
                         modgen_ram_ix167_a_253__dup_1080), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_1080), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2361 (.Q (
                         modgen_ram_ix167_a_252__dup_1081), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_1081), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2365 (.Q (
                         modgen_ram_ix167_a_251__dup_1082), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_1082), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2369 (.Q (
                         modgen_ram_ix167_a_250__dup_1083), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_1083), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2373 (.Q (
                         modgen_ram_ix167_a_249__dup_1084), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_1084), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2377 (.Q (
                         modgen_ram_ix167_a_248__dup_1085), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_1085), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2381 (.Q (
                         modgen_ram_ix167_a_247__dup_1086), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_1086), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2385 (.Q (
                         modgen_ram_ix167_a_246__dup_1087), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_1087), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2389 (.Q (
                         modgen_ram_ix167_a_245__dup_1088), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_1088), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2393 (.Q (
                         modgen_ram_ix167_a_244__dup_1089), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_1089), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2397 (.Q (
                         modgen_ram_ix167_a_243__dup_1090), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_1090), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2401 (.Q (
                         modgen_ram_ix167_a_242__dup_1091), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_1091), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2405 (.Q (
                         modgen_ram_ix167_a_241__dup_1092), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_1092), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2409 (.Q (
                         modgen_ram_ix167_a_240__dup_1093), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_1093), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2413 (.Q (
                         modgen_ram_ix167_a_239__dup_1094), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_1094), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2417 (.Q (
                         modgen_ram_ix167_a_238__dup_1095), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_1095), .SN (nx28497)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2421 (.Q (
                         modgen_ram_ix167_a_237__dup_1096), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_1096), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2425 (.Q (
                         modgen_ram_ix167_a_236__dup_1097), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_1097), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2429 (.Q (
                         modgen_ram_ix167_a_235__dup_1098), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_1098), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2433 (.Q (
                         modgen_ram_ix167_a_234__dup_1099), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_1099), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2437 (.Q (
                         modgen_ram_ix167_a_233__dup_1100), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_1100), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2441 (.Q (
                         modgen_ram_ix167_a_232__dup_1101), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_1101), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2445 (.Q (
                         modgen_ram_ix167_a_231__dup_1102), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_1102), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2449 (.Q (
                         modgen_ram_ix167_a_230__dup_1103), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_1103), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2453 (.Q (
                         modgen_ram_ix167_a_229__dup_1104), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_1104), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2457 (.Q (
                         modgen_ram_ix167_a_228__dup_1105), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_1105), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2461 (.Q (
                         modgen_ram_ix167_a_227__dup_1106), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_1106), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2465 (.Q (
                         modgen_ram_ix167_a_226__dup_1107), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_1107), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2469 (.Q (
                         modgen_ram_ix167_a_225__dup_1108), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_1108), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2473 (.Q (
                         modgen_ram_ix167_a_224__dup_1109), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_1109), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2477 (.Q (
                         modgen_ram_ix167_a_223__dup_1110), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_1110), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2481 (.Q (
                         modgen_ram_ix167_a_222__dup_1111), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_1111), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2485 (.Q (
                         modgen_ram_ix167_a_221__dup_1112), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_1112), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2489 (.Q (
                         modgen_ram_ix167_a_220__dup_1113), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_1113), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2493 (.Q (
                         modgen_ram_ix167_a_219__dup_1114), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_1114), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2497 (.Q (
                         modgen_ram_ix167_a_218__dup_1115), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_1115), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2501 (.Q (
                         modgen_ram_ix167_a_217__dup_1116), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_1116), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2505 (.Q (
                         modgen_ram_ix167_a_216__dup_1117), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_1117), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2509 (.Q (
                         modgen_ram_ix167_a_215__dup_1118), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_1118), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2513 (.Q (
                         modgen_ram_ix167_a_214__dup_1119), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_1119), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2517 (.Q (
                         modgen_ram_ix167_a_213__dup_1120), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_1120), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2521 (.Q (
                         modgen_ram_ix167_a_212__dup_1121), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_1121), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2525 (.Q (
                         modgen_ram_ix167_a_211__dup_1122), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_1122), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2529 (.Q (
                         modgen_ram_ix167_a_210__dup_1123), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_1123), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2533 (.Q (
                         modgen_ram_ix167_a_209__dup_1124), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_1124), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2537 (.Q (
                         modgen_ram_ix167_a_208__dup_1125), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_1125), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2541 (.Q (
                         modgen_ram_ix167_a_207__dup_1126), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_1126), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2545 (.Q (
                         modgen_ram_ix167_a_206__dup_1127), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_1127), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2549 (.Q (
                         modgen_ram_ix167_a_205__dup_1128), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_1128), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2553 (.Q (
                         modgen_ram_ix167_a_204__dup_1129), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_1129), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2557 (.Q (
                         modgen_ram_ix167_a_203__dup_1130), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_1130), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2561 (.Q (
                         modgen_ram_ix167_a_202__dup_1131), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_1131), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2565 (.Q (
                         modgen_ram_ix167_a_201__dup_1132), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_1132), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2569 (.Q (
                         modgen_ram_ix167_a_200__dup_1133), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_1133), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2573 (.Q (
                         modgen_ram_ix167_a_199__dup_1134), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_1134), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2577 (.Q (
                         modgen_ram_ix167_a_198__dup_1135), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_1135), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2581 (.Q (
                         modgen_ram_ix167_a_197__dup_1136), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_1136), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2585 (.Q (
                         modgen_ram_ix167_a_196__dup_1137), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_1137), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2589 (.Q (
                         modgen_ram_ix167_a_195__dup_1138), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_1138), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2593 (.Q (
                         modgen_ram_ix167_a_194__dup_1139), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_1139), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2597 (.Q (
                         modgen_ram_ix167_a_193__dup_1140), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_1140), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2601 (.Q (
                         modgen_ram_ix167_a_192__dup_1141), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_1141), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2605 (.Q (
                         modgen_ram_ix167_a_191__dup_1142), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_1142), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2609 (.Q (
                         modgen_ram_ix167_a_190__dup_1143), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_1143), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2613 (.Q (
                         modgen_ram_ix167_a_189__dup_1144), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_1144), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2617 (.Q (
                         modgen_ram_ix167_a_188__dup_1145), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_1145), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2621 (.Q (
                         modgen_ram_ix167_a_187__dup_1146), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_1146), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2625 (.Q (
                         modgen_ram_ix167_a_186__dup_1147), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_1147), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2629 (.Q (
                         modgen_ram_ix167_a_185__dup_1148), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_1148), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2633 (.Q (
                         modgen_ram_ix167_a_184__dup_1149), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_1149), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2637 (.Q (
                         modgen_ram_ix167_a_183__dup_1150), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_1150), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2641 (.Q (
                         modgen_ram_ix167_a_182__dup_1151), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_1151), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2645 (.Q (
                         modgen_ram_ix167_a_181__dup_1152), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_1152), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2649 (.Q (
                         modgen_ram_ix167_a_180__dup_1153), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_1153), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2653 (.Q (
                         modgen_ram_ix167_a_179__dup_1154), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_1154), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2657 (.Q (
                         modgen_ram_ix167_a_178__dup_1155), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_1155), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2661 (.Q (
                         modgen_ram_ix167_a_177__dup_1156), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_1156), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2665 (.Q (
                         modgen_ram_ix167_a_176__dup_1157), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_1157), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2669 (.Q (
                         modgen_ram_ix167_a_175__dup_1158), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_1158), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2673 (.Q (
                         modgen_ram_ix167_a_174__dup_1159), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_1159), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2677 (.Q (
                         modgen_ram_ix167_a_173__dup_1160), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_1160), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2681 (.Q (
                         modgen_ram_ix167_a_172__dup_1161), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_1161), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2685 (.Q (
                         modgen_ram_ix167_a_171__dup_1162), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_1162), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2689 (.Q (
                         modgen_ram_ix167_a_170__dup_1163), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_1163), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2693 (.Q (
                         modgen_ram_ix167_a_169__dup_1164), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_1164), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2697 (.Q (
                         modgen_ram_ix167_a_168__dup_1165), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_1165), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2701 (.Q (
                         modgen_ram_ix167_a_167__dup_1166), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_1166), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2705 (.Q (
                         modgen_ram_ix167_a_166__dup_1167), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_1167), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2709 (.Q (
                         modgen_ram_ix167_a_165__dup_1168), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_1168), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2713 (.Q (
                         modgen_ram_ix167_a_164__dup_1169), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_1169), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2717 (.Q (
                         modgen_ram_ix167_a_163__dup_1170), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_1170), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2721 (.Q (
                         modgen_ram_ix167_a_162__dup_1171), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_1171), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2725 (.Q (
                         modgen_ram_ix167_a_161__dup_1172), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_1172), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2729 (.Q (
                         modgen_ram_ix167_a_160__dup_1173), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_1173), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2733 (.Q (
                         modgen_ram_ix167_a_159__dup_1174), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_1174), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2737 (.Q (
                         modgen_ram_ix167_a_158__dup_1175), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_1175), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2741 (.Q (
                         modgen_ram_ix167_a_157__dup_1176), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_1176), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2745 (.Q (
                         modgen_ram_ix167_a_156__dup_1177), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_1177), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2749 (.Q (
                         modgen_ram_ix167_a_155__dup_1178), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_1178), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2753 (.Q (
                         modgen_ram_ix167_a_154__dup_1179), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_1179), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2757 (.Q (
                         modgen_ram_ix167_a_153__dup_1180), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_1180), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2761 (.Q (
                         modgen_ram_ix167_a_152__dup_1181), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_1181), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2765 (.Q (
                         modgen_ram_ix167_a_151__dup_1182), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_1182), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2769 (.Q (
                         modgen_ram_ix167_a_150__dup_1183), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_1183), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2773 (.Q (
                         modgen_ram_ix167_a_149__dup_1184), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_1184), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2777 (.Q (
                         modgen_ram_ix167_a_148__dup_1185), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_1185), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2781 (.Q (
                         modgen_ram_ix167_a_147__dup_1186), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_1186), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2785 (.Q (
                         modgen_ram_ix167_a_146__dup_1187), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_1187), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2789 (.Q (
                         modgen_ram_ix167_a_145__dup_1188), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_1188), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2793 (.Q (
                         modgen_ram_ix167_a_144__dup_1189), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_1189), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2797 (.Q (
                         modgen_ram_ix167_a_143__dup_1190), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_1190), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2801 (.Q (
                         modgen_ram_ix167_a_142__dup_1191), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_1191), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2805 (.Q (
                         modgen_ram_ix167_a_141__dup_1192), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_1192), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2809 (.Q (
                         modgen_ram_ix167_a_140__dup_1193), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_1193), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2813 (.Q (
                         modgen_ram_ix167_a_139__dup_1194), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_1194), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2817 (.Q (
                         modgen_ram_ix167_a_138__dup_1195), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_1195), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2821 (.Q (
                         modgen_ram_ix167_a_137__dup_1196), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_1196), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2825 (.Q (
                         modgen_ram_ix167_a_136__dup_1197), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_1197), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2829 (.Q (
                         modgen_ram_ix167_a_135__dup_1198), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_1198), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2833 (.Q (
                         modgen_ram_ix167_a_134__dup_1199), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_1199), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2837 (.Q (
                         modgen_ram_ix167_a_133__dup_1200), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_1200), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2841 (.Q (
                         modgen_ram_ix167_a_132__dup_1201), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_1201), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2845 (.Q (
                         modgen_ram_ix167_a_131__dup_1202), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_1202), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2849 (.Q (
                         modgen_ram_ix167_a_130__dup_1203), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_1203), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2853 (.Q (
                         modgen_ram_ix167_a_129__dup_1204), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_1204), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2857 (.Q (
                         modgen_ram_ix167_a_128__dup_1205), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_1205), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2861 (.Q (
                         modgen_ram_ix167_a_127__dup_1206), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_1206), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2865 (.Q (
                         modgen_ram_ix167_a_126__dup_1207), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_1207), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2869 (.Q (
                         modgen_ram_ix167_a_125__dup_1208), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_1208), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2873 (.Q (
                         modgen_ram_ix167_a_124__dup_1209), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_1209), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2877 (.Q (
                         modgen_ram_ix167_a_123__dup_1210), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_1210), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2881 (.Q (
                         modgen_ram_ix167_a_122__dup_1211), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_1211), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2885 (.Q (
                         modgen_ram_ix167_a_121__dup_1212), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_1212), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2889 (.Q (
                         modgen_ram_ix167_a_120__dup_1213), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_1213), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2893 (.Q (
                         modgen_ram_ix167_a_119__dup_1214), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_1214), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2897 (.Q (
                         modgen_ram_ix167_a_118__dup_1215), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_1215), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2901 (.Q (
                         modgen_ram_ix167_a_117__dup_1216), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_1216), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2905 (.Q (
                         modgen_ram_ix167_a_116__dup_1217), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_1217), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2909 (.Q (
                         modgen_ram_ix167_a_115__dup_1218), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_1218), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2913 (.Q (
                         modgen_ram_ix167_a_114__dup_1219), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_1219), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2917 (.Q (
                         modgen_ram_ix167_a_113__dup_1220), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_1220), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2921 (.Q (
                         modgen_ram_ix167_a_112__dup_1221), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_1221), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2925 (.Q (
                         modgen_ram_ix167_a_111__dup_1222), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_1222), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2929 (.Q (
                         modgen_ram_ix167_a_110__dup_1223), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_1223), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2933 (.Q (
                         modgen_ram_ix167_a_109__dup_1224), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_1224), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2937 (.Q (
                         modgen_ram_ix167_a_108__dup_1225), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_1225), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2941 (.Q (
                         modgen_ram_ix167_a_107__dup_1226), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_1226), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2945 (.Q (
                         modgen_ram_ix167_a_106__dup_1227), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_1227), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2949 (.Q (
                         modgen_ram_ix167_a_105__dup_1228), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_1228), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2953 (.Q (
                         modgen_ram_ix167_a_104__dup_1229), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_1229), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2957 (.Q (
                         modgen_ram_ix167_a_103__dup_1230), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_1230), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2961 (.Q (
                         modgen_ram_ix167_a_102__dup_1231), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_1231), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2965 (.Q (
                         modgen_ram_ix167_a_101__dup_1232), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_1232), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2969 (.Q (
                         modgen_ram_ix167_a_100__dup_1233), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_1233), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2973 (.Q (
                         modgen_ram_ix167_a_99__dup_1234), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_1234), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2977 (.Q (
                         modgen_ram_ix167_a_98__dup_1235), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_1235), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2981 (.Q (
                         modgen_ram_ix167_a_97__dup_1236), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_1236), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2985 (.Q (
                         modgen_ram_ix167_a_96__dup_1237), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_1237), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2989 (.Q (
                         modgen_ram_ix167_a_95__dup_1238), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_1238), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2993 (.Q (
                         modgen_ram_ix167_a_94__dup_1239), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_1239), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix2997 (.Q (
                         modgen_ram_ix167_a_93__dup_1240), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_1240), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3001 (.Q (
                         modgen_ram_ix167_a_92__dup_1241), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_1241), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3005 (.Q (
                         modgen_ram_ix167_a_91__dup_1242), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_1242), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3009 (.Q (
                         modgen_ram_ix167_a_90__dup_1243), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_1243), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3013 (.Q (
                         modgen_ram_ix167_a_89__dup_1244), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_1244), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3017 (.Q (
                         modgen_ram_ix167_a_88__dup_1245), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_1245), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3021 (.Q (
                         modgen_ram_ix167_a_87__dup_1246), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_1246), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3025 (.Q (
                         modgen_ram_ix167_a_86__dup_1247), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_1247), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3029 (.Q (
                         modgen_ram_ix167_a_85__dup_1248), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_1248), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3033 (.Q (
                         modgen_ram_ix167_a_84__dup_1249), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_1249), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3037 (.Q (
                         modgen_ram_ix167_a_83__dup_1250), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_1250), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3041 (.Q (
                         modgen_ram_ix167_a_82__dup_1251), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_1251), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3045 (.Q (
                         modgen_ram_ix167_a_81__dup_1252), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_1252), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3049 (.Q (
                         modgen_ram_ix167_a_80__dup_1253), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_1253), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3053 (.Q (
                         modgen_ram_ix167_a_79__dup_1254), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_1254), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3057 (.Q (
                         modgen_ram_ix167_a_78__dup_1255), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_1255), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3061 (.Q (
                         modgen_ram_ix167_a_77__dup_1256), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_1256), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3065 (.Q (
                         modgen_ram_ix167_a_76__dup_1257), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_1257), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3069 (.Q (
                         modgen_ram_ix167_a_75__dup_1258), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_1258), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3073 (.Q (
                         modgen_ram_ix167_a_74__dup_1259), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_1259), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3077 (.Q (
                         modgen_ram_ix167_a_73__dup_1260), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_1260), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3081 (.Q (
                         modgen_ram_ix167_a_72__dup_1261), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_1261), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3085 (.Q (
                         modgen_ram_ix167_a_71__dup_1262), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_1262), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3089 (.Q (
                         modgen_ram_ix167_a_70__dup_1263), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_1263), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3093 (.Q (
                         modgen_ram_ix167_a_69__dup_1264), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_1264), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3097 (.Q (
                         modgen_ram_ix167_a_68__dup_1265), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_1265), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3101 (.Q (
                         modgen_ram_ix167_a_67__dup_1266), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_1266), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3105 (.Q (
                         modgen_ram_ix167_a_66__dup_1267), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_1267), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3109 (.Q (
                         modgen_ram_ix167_a_65__dup_1268), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_1268), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3113 (.Q (
                         modgen_ram_ix167_a_64__dup_1269), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_1269), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3117 (.Q (
                         modgen_ram_ix167_a_63__dup_1270), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_1270), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3121 (.Q (
                         modgen_ram_ix167_a_62__dup_1271), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_1271), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3125 (.Q (
                         modgen_ram_ix167_a_61__dup_1272), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_1272), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3129 (.Q (
                         modgen_ram_ix167_a_60__dup_1273), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_1273), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3133 (.Q (
                         modgen_ram_ix167_a_59__dup_1274), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_1274), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3137 (.Q (
                         modgen_ram_ix167_a_58__dup_1275), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_1275), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3141 (.Q (
                         modgen_ram_ix167_a_57__dup_1276), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_1276), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3145 (.Q (
                         modgen_ram_ix167_a_56__dup_1277), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_1277), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3149 (.Q (
                         modgen_ram_ix167_a_55__dup_1278), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_1278), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3153 (.Q (
                         modgen_ram_ix167_a_54__dup_1279), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_1279), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3157 (.Q (
                         modgen_ram_ix167_a_53__dup_1280), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_1280), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3161 (.Q (
                         modgen_ram_ix167_a_52__dup_1281), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_1281), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3165 (.Q (
                         modgen_ram_ix167_a_51__dup_1282), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_1282), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3169 (.Q (
                         modgen_ram_ix167_a_50__dup_1283), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_1283), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3173 (.Q (
                         modgen_ram_ix167_a_49__dup_1284), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_1284), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3177 (.Q (
                         modgen_ram_ix167_a_48__dup_1285), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_1285), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3181 (.Q (
                         modgen_ram_ix167_a_47__dup_1286), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_1286), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3185 (.Q (
                         modgen_ram_ix167_a_46__dup_1287), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_1287), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3189 (.Q (
                         modgen_ram_ix167_a_45__dup_1288), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_1288), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3193 (.Q (
                         modgen_ram_ix167_a_44__dup_1289), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_1289), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3197 (.Q (
                         modgen_ram_ix167_a_43__dup_1290), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_1290), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3201 (.Q (
                         modgen_ram_ix167_a_42__dup_1291), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_1291), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3205 (.Q (
                         modgen_ram_ix167_a_41__dup_1292), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_1292), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3209 (.Q (
                         modgen_ram_ix167_a_40__dup_1293), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_1293), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3213 (.Q (
                         modgen_ram_ix167_a_39__dup_1294), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_1294), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3217 (.Q (
                         modgen_ram_ix167_a_38__dup_1295), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_1295), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3221 (.Q (
                         modgen_ram_ix167_a_37__dup_1296), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_1296), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3225 (.Q (
                         modgen_ram_ix167_a_36__dup_1297), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_1297), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3229 (.Q (
                         modgen_ram_ix167_a_35__dup_1298), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_1298), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3233 (.Q (
                         modgen_ram_ix167_a_34__dup_1299), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_1299), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3237 (.Q (
                         modgen_ram_ix167_a_33__dup_1300), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_1300), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3241 (.Q (
                         modgen_ram_ix167_a_32__dup_1301), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_1301), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3245 (.Q (
                         modgen_ram_ix167_a_31__dup_1302), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_1302), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3249 (.Q (
                         modgen_ram_ix167_a_30__dup_1303), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_1303), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3253 (.Q (
                         modgen_ram_ix167_a_29__dup_1304), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_1304), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3257 (.Q (
                         modgen_ram_ix167_a_28__dup_1305), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_1305), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3261 (.Q (
                         modgen_ram_ix167_a_27__dup_1306), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_1306), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3265 (.Q (
                         modgen_ram_ix167_a_26__dup_1307), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_1307), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3269 (.Q (
                         modgen_ram_ix167_a_25__dup_1308), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_1308), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3273 (.Q (
                         modgen_ram_ix167_a_24__dup_1309), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_1309), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3277 (.Q (
                         modgen_ram_ix167_a_23__dup_1310), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_1310), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3281 (.Q (
                         modgen_ram_ix167_a_22__dup_1311), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_1311), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3285 (.Q (
                         modgen_ram_ix167_a_21__dup_1312), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_1312), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3289 (.Q (
                         modgen_ram_ix167_a_20__dup_1313), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_1313), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3293 (.Q (
                         modgen_ram_ix167_a_19__dup_1314), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_1314), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3297 (.Q (
                         modgen_ram_ix167_a_18__dup_1315), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_1315), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3301 (.Q (
                         modgen_ram_ix167_a_17__dup_1316), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_1316), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3305 (.Q (
                         modgen_ram_ix167_a_16__dup_1317), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_1317), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3309 (.Q (
                         modgen_ram_ix167_a_15__dup_1318), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_1318), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3313 (.Q (
                         modgen_ram_ix167_a_14__dup_1319), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_1319), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3317 (.Q (
                         modgen_ram_ix167_a_13__dup_1320), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_1320), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3321 (.Q (
                         modgen_ram_ix167_a_12__dup_1321), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_1321), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3325 (.Q (
                         modgen_ram_ix167_a_11__dup_1322), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_1322), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3329 (.Q (
                         modgen_ram_ix167_a_10__dup_1323), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_1323), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3333 (.Q (
                         modgen_ram_ix167_a_9__dup_1324), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_1324), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3337 (.Q (
                         modgen_ram_ix167_a_8__dup_1325), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_1325), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3341 (.Q (
                         modgen_ram_ix167_a_7__dup_1326), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_1326), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3345 (.Q (
                         modgen_ram_ix167_a_6__dup_1327), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_1327), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3349 (.Q (
                         modgen_ram_ix167_a_5__dup_1328), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_1328), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3353 (.Q (
                         modgen_ram_ix167_a_4__dup_1329), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_1329), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3357 (.Q (
                         modgen_ram_ix167_a_3__dup_1330), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_1330), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3361 (.Q (
                         modgen_ram_ix167_a_2__dup_1331), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_1331), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3365 (.Q (
                         modgen_ram_ix167_a_1__dup_1332), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_1332), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3369 (.Q (
                         modgen_ram_ix167_a_0__dup_1333), .CK (wb_clk_i), .D (
                         nx28513), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_1333), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3374 (.Q (
                         modgen_ram_ix167_a_255__dup_1342), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_1342), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3378 (.Q (
                         modgen_ram_ix167_a_254__dup_1343), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_1343), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3382 (.Q (
                         modgen_ram_ix167_a_253__dup_1344), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_1344), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3386 (.Q (
                         modgen_ram_ix167_a_252__dup_1345), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_1345), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3390 (.Q (
                         modgen_ram_ix167_a_251__dup_1346), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_1346), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3394 (.Q (
                         modgen_ram_ix167_a_250__dup_1347), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_1347), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3398 (.Q (
                         modgen_ram_ix167_a_249__dup_1348), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_1348), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3402 (.Q (
                         modgen_ram_ix167_a_248__dup_1349), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_1349), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3406 (.Q (
                         modgen_ram_ix167_a_247__dup_1350), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_1350), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3410 (.Q (
                         modgen_ram_ix167_a_246__dup_1351), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_1351), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3414 (.Q (
                         modgen_ram_ix167_a_245__dup_1352), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_1352), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3418 (.Q (
                         modgen_ram_ix167_a_244__dup_1353), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_1353), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3422 (.Q (
                         modgen_ram_ix167_a_243__dup_1354), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_1354), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3426 (.Q (
                         modgen_ram_ix167_a_242__dup_1355), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_1355), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3430 (.Q (
                         modgen_ram_ix167_a_241__dup_1356), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_1356), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3434 (.Q (
                         modgen_ram_ix167_a_240__dup_1357), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_1357), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3438 (.Q (
                         modgen_ram_ix167_a_239__dup_1358), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_1358), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3442 (.Q (
                         modgen_ram_ix167_a_238__dup_1359), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_1359), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3446 (.Q (
                         modgen_ram_ix167_a_237__dup_1360), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_1360), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3450 (.Q (
                         modgen_ram_ix167_a_236__dup_1361), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_1361), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3454 (.Q (
                         modgen_ram_ix167_a_235__dup_1362), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_1362), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3458 (.Q (
                         modgen_ram_ix167_a_234__dup_1363), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_1363), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3462 (.Q (
                         modgen_ram_ix167_a_233__dup_1364), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_1364), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3466 (.Q (
                         modgen_ram_ix167_a_232__dup_1365), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_1365), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3470 (.Q (
                         modgen_ram_ix167_a_231__dup_1366), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_1366), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3474 (.Q (
                         modgen_ram_ix167_a_230__dup_1367), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_1367), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3478 (.Q (
                         modgen_ram_ix167_a_229__dup_1368), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_1368), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3482 (.Q (
                         modgen_ram_ix167_a_228__dup_1369), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_1369), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3486 (.Q (
                         modgen_ram_ix167_a_227__dup_1370), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_1370), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3490 (.Q (
                         modgen_ram_ix167_a_226__dup_1371), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_1371), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3494 (.Q (
                         modgen_ram_ix167_a_225__dup_1372), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_1372), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3498 (.Q (
                         modgen_ram_ix167_a_224__dup_1373), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_1373), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3502 (.Q (
                         modgen_ram_ix167_a_223__dup_1374), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_1374), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3506 (.Q (
                         modgen_ram_ix167_a_222__dup_1375), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_1375), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3510 (.Q (
                         modgen_ram_ix167_a_221__dup_1376), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_1376), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3514 (.Q (
                         modgen_ram_ix167_a_220__dup_1377), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_1377), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3518 (.Q (
                         modgen_ram_ix167_a_219__dup_1378), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_1378), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3522 (.Q (
                         modgen_ram_ix167_a_218__dup_1379), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_1379), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3526 (.Q (
                         modgen_ram_ix167_a_217__dup_1380), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_1380), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3530 (.Q (
                         modgen_ram_ix167_a_216__dup_1381), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_1381), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3534 (.Q (
                         modgen_ram_ix167_a_215__dup_1382), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_1382), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3538 (.Q (
                         modgen_ram_ix167_a_214__dup_1383), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_1383), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3542 (.Q (
                         modgen_ram_ix167_a_213__dup_1384), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_1384), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3546 (.Q (
                         modgen_ram_ix167_a_212__dup_1385), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_1385), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3550 (.Q (
                         modgen_ram_ix167_a_211__dup_1386), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_1386), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3554 (.Q (
                         modgen_ram_ix167_a_210__dup_1387), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_1387), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3558 (.Q (
                         modgen_ram_ix167_a_209__dup_1388), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_1388), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3562 (.Q (
                         modgen_ram_ix167_a_208__dup_1389), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_1389), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3566 (.Q (
                         modgen_ram_ix167_a_207__dup_1390), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_1390), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3570 (.Q (
                         modgen_ram_ix167_a_206__dup_1391), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_1391), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3574 (.Q (
                         modgen_ram_ix167_a_205__dup_1392), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_1392), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3578 (.Q (
                         modgen_ram_ix167_a_204__dup_1393), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_1393), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3582 (.Q (
                         modgen_ram_ix167_a_203__dup_1394), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_1394), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3586 (.Q (
                         modgen_ram_ix167_a_202__dup_1395), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_1395), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3590 (.Q (
                         modgen_ram_ix167_a_201__dup_1396), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_1396), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3594 (.Q (
                         modgen_ram_ix167_a_200__dup_1397), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_1397), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3598 (.Q (
                         modgen_ram_ix167_a_199__dup_1398), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_1398), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3602 (.Q (
                         modgen_ram_ix167_a_198__dup_1399), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_1399), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3606 (.Q (
                         modgen_ram_ix167_a_197__dup_1400), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_1400), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3610 (.Q (
                         modgen_ram_ix167_a_196__dup_1401), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_1401), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3614 (.Q (
                         modgen_ram_ix167_a_195__dup_1402), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_1402), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3618 (.Q (
                         modgen_ram_ix167_a_194__dup_1403), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_1403), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3622 (.Q (
                         modgen_ram_ix167_a_193__dup_1404), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_1404), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3626 (.Q (
                         modgen_ram_ix167_a_192__dup_1405), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_1405), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3630 (.Q (
                         modgen_ram_ix167_a_191__dup_1406), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_1406), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3634 (.Q (
                         modgen_ram_ix167_a_190__dup_1407), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_1407), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3638 (.Q (
                         modgen_ram_ix167_a_189__dup_1408), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_1408), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3642 (.Q (
                         modgen_ram_ix167_a_188__dup_1409), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_1409), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3646 (.Q (
                         modgen_ram_ix167_a_187__dup_1410), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_1410), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3650 (.Q (
                         modgen_ram_ix167_a_186__dup_1411), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_1411), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3654 (.Q (
                         modgen_ram_ix167_a_185__dup_1412), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_1412), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3658 (.Q (
                         modgen_ram_ix167_a_184__dup_1413), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_1413), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3662 (.Q (
                         modgen_ram_ix167_a_183__dup_1414), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_1414), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3666 (.Q (
                         modgen_ram_ix167_a_182__dup_1415), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_1415), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3670 (.Q (
                         modgen_ram_ix167_a_181__dup_1416), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_1416), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3674 (.Q (
                         modgen_ram_ix167_a_180__dup_1417), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_1417), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3678 (.Q (
                         modgen_ram_ix167_a_179__dup_1418), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_1418), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3682 (.Q (
                         modgen_ram_ix167_a_178__dup_1419), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_1419), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3686 (.Q (
                         modgen_ram_ix167_a_177__dup_1420), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_1420), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3690 (.Q (
                         modgen_ram_ix167_a_176__dup_1421), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_1421), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3694 (.Q (
                         modgen_ram_ix167_a_175__dup_1422), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_1422), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3698 (.Q (
                         modgen_ram_ix167_a_174__dup_1423), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_1423), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3702 (.Q (
                         modgen_ram_ix167_a_173__dup_1424), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_1424), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3706 (.Q (
                         modgen_ram_ix167_a_172__dup_1425), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_1425), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3710 (.Q (
                         modgen_ram_ix167_a_171__dup_1426), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_1426), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3714 (.Q (
                         modgen_ram_ix167_a_170__dup_1427), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_1427), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3718 (.Q (
                         modgen_ram_ix167_a_169__dup_1428), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_1428), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3722 (.Q (
                         modgen_ram_ix167_a_168__dup_1429), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_1429), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3726 (.Q (
                         modgen_ram_ix167_a_167__dup_1430), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_1430), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3730 (.Q (
                         modgen_ram_ix167_a_166__dup_1431), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_1431), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3734 (.Q (
                         modgen_ram_ix167_a_165__dup_1432), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_1432), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3738 (.Q (
                         modgen_ram_ix167_a_164__dup_1433), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_1433), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3742 (.Q (
                         modgen_ram_ix167_a_163__dup_1434), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_1434), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3746 (.Q (
                         modgen_ram_ix167_a_162__dup_1435), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_1435), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3750 (.Q (
                         modgen_ram_ix167_a_161__dup_1436), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_1436), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3754 (.Q (
                         modgen_ram_ix167_a_160__dup_1437), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_1437), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3758 (.Q (
                         modgen_ram_ix167_a_159__dup_1438), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_1438), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3762 (.Q (
                         modgen_ram_ix167_a_158__dup_1439), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_1439), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3766 (.Q (
                         modgen_ram_ix167_a_157__dup_1440), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_1440), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3770 (.Q (
                         modgen_ram_ix167_a_156__dup_1441), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_1441), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3774 (.Q (
                         modgen_ram_ix167_a_155__dup_1442), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_1442), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3778 (.Q (
                         modgen_ram_ix167_a_154__dup_1443), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_1443), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3782 (.Q (
                         modgen_ram_ix167_a_153__dup_1444), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_1444), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3786 (.Q (
                         modgen_ram_ix167_a_152__dup_1445), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_1445), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3790 (.Q (
                         modgen_ram_ix167_a_151__dup_1446), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_1446), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3794 (.Q (
                         modgen_ram_ix167_a_150__dup_1447), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_1447), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3798 (.Q (
                         modgen_ram_ix167_a_149__dup_1448), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_1448), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3802 (.Q (
                         modgen_ram_ix167_a_148__dup_1449), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_1449), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3806 (.Q (
                         modgen_ram_ix167_a_147__dup_1450), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_1450), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3810 (.Q (
                         modgen_ram_ix167_a_146__dup_1451), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_1451), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3814 (.Q (
                         modgen_ram_ix167_a_145__dup_1452), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_1452), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3818 (.Q (
                         modgen_ram_ix167_a_144__dup_1453), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_1453), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3822 (.Q (
                         modgen_ram_ix167_a_143__dup_1454), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_1454), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3826 (.Q (
                         modgen_ram_ix167_a_142__dup_1455), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_1455), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3830 (.Q (
                         modgen_ram_ix167_a_141__dup_1456), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_1456), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3834 (.Q (
                         modgen_ram_ix167_a_140__dup_1457), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_1457), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3838 (.Q (
                         modgen_ram_ix167_a_139__dup_1458), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_1458), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3842 (.Q (
                         modgen_ram_ix167_a_138__dup_1459), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_1459), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3846 (.Q (
                         modgen_ram_ix167_a_137__dup_1460), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_1460), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3850 (.Q (
                         modgen_ram_ix167_a_136__dup_1461), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_1461), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3854 (.Q (
                         modgen_ram_ix167_a_135__dup_1462), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_1462), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3858 (.Q (
                         modgen_ram_ix167_a_134__dup_1463), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_1463), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3862 (.Q (
                         modgen_ram_ix167_a_133__dup_1464), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_1464), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3866 (.Q (
                         modgen_ram_ix167_a_132__dup_1465), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_1465), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3870 (.Q (
                         modgen_ram_ix167_a_131__dup_1466), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_1466), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3874 (.Q (
                         modgen_ram_ix167_a_130__dup_1467), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_1467), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3878 (.Q (
                         modgen_ram_ix167_a_129__dup_1468), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_1468), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3882 (.Q (
                         modgen_ram_ix167_a_128__dup_1469), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_1469), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3886 (.Q (
                         modgen_ram_ix167_a_127__dup_1470), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_1470), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3890 (.Q (
                         modgen_ram_ix167_a_126__dup_1471), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_1471), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3894 (.Q (
                         modgen_ram_ix167_a_125__dup_1472), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_1472), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3898 (.Q (
                         modgen_ram_ix167_a_124__dup_1473), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_1473), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3902 (.Q (
                         modgen_ram_ix167_a_123__dup_1474), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_1474), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3906 (.Q (
                         modgen_ram_ix167_a_122__dup_1475), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_1475), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3910 (.Q (
                         modgen_ram_ix167_a_121__dup_1476), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_1476), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3914 (.Q (
                         modgen_ram_ix167_a_120__dup_1477), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_1477), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3918 (.Q (
                         modgen_ram_ix167_a_119__dup_1478), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_1478), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3922 (.Q (
                         modgen_ram_ix167_a_118__dup_1479), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_1479), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3926 (.Q (
                         modgen_ram_ix167_a_117__dup_1480), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_1480), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3930 (.Q (
                         modgen_ram_ix167_a_116__dup_1481), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_1481), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3934 (.Q (
                         modgen_ram_ix167_a_115__dup_1482), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_1482), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3938 (.Q (
                         modgen_ram_ix167_a_114__dup_1483), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_1483), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3942 (.Q (
                         modgen_ram_ix167_a_113__dup_1484), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_1484), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3946 (.Q (
                         modgen_ram_ix167_a_112__dup_1485), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_1485), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3950 (.Q (
                         modgen_ram_ix167_a_111__dup_1486), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_1486), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3954 (.Q (
                         modgen_ram_ix167_a_110__dup_1487), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_1487), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3958 (.Q (
                         modgen_ram_ix167_a_109__dup_1488), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_1488), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3962 (.Q (
                         modgen_ram_ix167_a_108__dup_1489), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_1489), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3966 (.Q (
                         modgen_ram_ix167_a_107__dup_1490), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_1490), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3970 (.Q (
                         modgen_ram_ix167_a_106__dup_1491), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_1491), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3974 (.Q (
                         modgen_ram_ix167_a_105__dup_1492), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_1492), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3978 (.Q (
                         modgen_ram_ix167_a_104__dup_1493), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_1493), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3982 (.Q (
                         modgen_ram_ix167_a_103__dup_1494), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_1494), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3986 (.Q (
                         modgen_ram_ix167_a_102__dup_1495), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_1495), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3990 (.Q (
                         modgen_ram_ix167_a_101__dup_1496), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_1496), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3994 (.Q (
                         modgen_ram_ix167_a_100__dup_1497), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_1497), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix3998 (.Q (
                         modgen_ram_ix167_a_99__dup_1498), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_1498), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4002 (.Q (
                         modgen_ram_ix167_a_98__dup_1499), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_1499), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4006 (.Q (
                         modgen_ram_ix167_a_97__dup_1500), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_1500), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4010 (.Q (
                         modgen_ram_ix167_a_96__dup_1501), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_1501), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4014 (.Q (
                         modgen_ram_ix167_a_95__dup_1502), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_1502), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4018 (.Q (
                         modgen_ram_ix167_a_94__dup_1503), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_1503), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4022 (.Q (
                         modgen_ram_ix167_a_93__dup_1504), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_1504), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4026 (.Q (
                         modgen_ram_ix167_a_92__dup_1505), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_1505), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4030 (.Q (
                         modgen_ram_ix167_a_91__dup_1506), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_1506), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4034 (.Q (
                         modgen_ram_ix167_a_90__dup_1507), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_1507), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4038 (.Q (
                         modgen_ram_ix167_a_89__dup_1508), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_1508), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4042 (.Q (
                         modgen_ram_ix167_a_88__dup_1509), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_1509), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4046 (.Q (
                         modgen_ram_ix167_a_87__dup_1510), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_1510), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4050 (.Q (
                         modgen_ram_ix167_a_86__dup_1511), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_1511), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4054 (.Q (
                         modgen_ram_ix167_a_85__dup_1512), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_1512), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4058 (.Q (
                         modgen_ram_ix167_a_84__dup_1513), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_1513), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4062 (.Q (
                         modgen_ram_ix167_a_83__dup_1514), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_1514), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4066 (.Q (
                         modgen_ram_ix167_a_82__dup_1515), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_1515), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4070 (.Q (
                         modgen_ram_ix167_a_81__dup_1516), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_1516), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4074 (.Q (
                         modgen_ram_ix167_a_80__dup_1517), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_1517), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4078 (.Q (
                         modgen_ram_ix167_a_79__dup_1518), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_1518), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4082 (.Q (
                         modgen_ram_ix167_a_78__dup_1519), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_1519), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4086 (.Q (
                         modgen_ram_ix167_a_77__dup_1520), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_1520), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4090 (.Q (
                         modgen_ram_ix167_a_76__dup_1521), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_1521), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4094 (.Q (
                         modgen_ram_ix167_a_75__dup_1522), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_1522), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4098 (.Q (
                         modgen_ram_ix167_a_74__dup_1523), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_1523), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4102 (.Q (
                         modgen_ram_ix167_a_73__dup_1524), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_1524), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4106 (.Q (
                         modgen_ram_ix167_a_72__dup_1525), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_1525), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4110 (.Q (
                         modgen_ram_ix167_a_71__dup_1526), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_1526), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4114 (.Q (
                         modgen_ram_ix167_a_70__dup_1527), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_1527), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4118 (.Q (
                         modgen_ram_ix167_a_69__dup_1528), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_1528), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4122 (.Q (
                         modgen_ram_ix167_a_68__dup_1529), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_1529), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4126 (.Q (
                         modgen_ram_ix167_a_67__dup_1530), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_1530), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4130 (.Q (
                         modgen_ram_ix167_a_66__dup_1531), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_1531), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4134 (.Q (
                         modgen_ram_ix167_a_65__dup_1532), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_1532), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4138 (.Q (
                         modgen_ram_ix167_a_64__dup_1533), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_1533), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4142 (.Q (
                         modgen_ram_ix167_a_63__dup_1534), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_1534), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4146 (.Q (
                         modgen_ram_ix167_a_62__dup_1535), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_1535), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4150 (.Q (
                         modgen_ram_ix167_a_61__dup_1536), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_1536), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4154 (.Q (
                         modgen_ram_ix167_a_60__dup_1537), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_1537), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4158 (.Q (
                         modgen_ram_ix167_a_59__dup_1538), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_1538), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4162 (.Q (
                         modgen_ram_ix167_a_58__dup_1539), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_1539), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4166 (.Q (
                         modgen_ram_ix167_a_57__dup_1540), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_1540), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4170 (.Q (
                         modgen_ram_ix167_a_56__dup_1541), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_1541), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4174 (.Q (
                         modgen_ram_ix167_a_55__dup_1542), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_1542), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4178 (.Q (
                         modgen_ram_ix167_a_54__dup_1543), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_1543), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4182 (.Q (
                         modgen_ram_ix167_a_53__dup_1544), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_1544), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4186 (.Q (
                         modgen_ram_ix167_a_52__dup_1545), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_1545), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4190 (.Q (
                         modgen_ram_ix167_a_51__dup_1546), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_1546), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4194 (.Q (
                         modgen_ram_ix167_a_50__dup_1547), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_1547), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4198 (.Q (
                         modgen_ram_ix167_a_49__dup_1548), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_1548), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4202 (.Q (
                         modgen_ram_ix167_a_48__dup_1549), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_1549), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4206 (.Q (
                         modgen_ram_ix167_a_47__dup_1550), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_1550), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4210 (.Q (
                         modgen_ram_ix167_a_46__dup_1551), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_1551), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4214 (.Q (
                         modgen_ram_ix167_a_45__dup_1552), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_1552), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4218 (.Q (
                         modgen_ram_ix167_a_44__dup_1553), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_1553), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4222 (.Q (
                         modgen_ram_ix167_a_43__dup_1554), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_1554), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4226 (.Q (
                         modgen_ram_ix167_a_42__dup_1555), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_1555), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4230 (.Q (
                         modgen_ram_ix167_a_41__dup_1556), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_1556), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4234 (.Q (
                         modgen_ram_ix167_a_40__dup_1557), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_1557), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4238 (.Q (
                         modgen_ram_ix167_a_39__dup_1558), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_1558), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4242 (.Q (
                         modgen_ram_ix167_a_38__dup_1559), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_1559), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4246 (.Q (
                         modgen_ram_ix167_a_37__dup_1560), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_1560), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4250 (.Q (
                         modgen_ram_ix167_a_36__dup_1561), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_1561), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4254 (.Q (
                         modgen_ram_ix167_a_35__dup_1562), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_1562), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4258 (.Q (
                         modgen_ram_ix167_a_34__dup_1563), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_1563), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4262 (.Q (
                         modgen_ram_ix167_a_33__dup_1564), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_1564), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4266 (.Q (
                         modgen_ram_ix167_a_32__dup_1565), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_1565), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4270 (.Q (
                         modgen_ram_ix167_a_31__dup_1566), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_1566), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4274 (.Q (
                         modgen_ram_ix167_a_30__dup_1567), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_1567), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4278 (.Q (
                         modgen_ram_ix167_a_29__dup_1568), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_1568), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4282 (.Q (
                         modgen_ram_ix167_a_28__dup_1569), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_1569), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4286 (.Q (
                         modgen_ram_ix167_a_27__dup_1570), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_1570), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4290 (.Q (
                         modgen_ram_ix167_a_26__dup_1571), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_1571), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4294 (.Q (
                         modgen_ram_ix167_a_25__dup_1572), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_1572), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4298 (.Q (
                         modgen_ram_ix167_a_24__dup_1573), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_1573), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4302 (.Q (
                         modgen_ram_ix167_a_23__dup_1574), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_1574), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4306 (.Q (
                         modgen_ram_ix167_a_22__dup_1575), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_1575), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4310 (.Q (
                         modgen_ram_ix167_a_21__dup_1576), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_1576), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4314 (.Q (
                         modgen_ram_ix167_a_20__dup_1577), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_1577), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4318 (.Q (
                         modgen_ram_ix167_a_19__dup_1578), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_1578), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4322 (.Q (
                         modgen_ram_ix167_a_18__dup_1579), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_1579), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4326 (.Q (
                         modgen_ram_ix167_a_17__dup_1580), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_1580), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4330 (.Q (
                         modgen_ram_ix167_a_16__dup_1581), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_1581), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4334 (.Q (
                         modgen_ram_ix167_a_15__dup_1582), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_1582), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4338 (.Q (
                         modgen_ram_ix167_a_14__dup_1583), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_1583), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4342 (.Q (
                         modgen_ram_ix167_a_13__dup_1584), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_1584), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4346 (.Q (
                         modgen_ram_ix167_a_12__dup_1585), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_1585), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4350 (.Q (
                         modgen_ram_ix167_a_11__dup_1586), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_1586), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4354 (.Q (
                         modgen_ram_ix167_a_10__dup_1587), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_1587), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4358 (.Q (
                         modgen_ram_ix167_a_9__dup_1588), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_1588), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4362 (.Q (
                         modgen_ram_ix167_a_8__dup_1589), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_1589), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4366 (.Q (
                         modgen_ram_ix167_a_7__dup_1590), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_1590), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4370 (.Q (
                         modgen_ram_ix167_a_6__dup_1591), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_1591), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4374 (.Q (
                         modgen_ram_ix167_a_5__dup_1592), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_1592), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4378 (.Q (
                         modgen_ram_ix167_a_4__dup_1593), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_1593), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4382 (.Q (
                         modgen_ram_ix167_a_3__dup_1594), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_1594), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4386 (.Q (
                         modgen_ram_ix167_a_2__dup_1595), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_1595), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4390 (.Q (
                         modgen_ram_ix167_a_1__dup_1596), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_1596), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4394 (.Q (
                         modgen_ram_ix167_a_0__dup_1597), .CK (wb_clk_i), .D (
                         nx28515), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_1597), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4399 (.Q (
                         modgen_ram_ix167_a_255__dup_1606), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_1606), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4403 (.Q (
                         modgen_ram_ix167_a_254__dup_1607), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_1607), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4407 (.Q (
                         modgen_ram_ix167_a_253__dup_1608), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_1608), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4411 (.Q (
                         modgen_ram_ix167_a_252__dup_1609), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_1609), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4415 (.Q (
                         modgen_ram_ix167_a_251__dup_1610), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_1610), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4419 (.Q (
                         modgen_ram_ix167_a_250__dup_1611), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_1611), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4423 (.Q (
                         modgen_ram_ix167_a_249__dup_1612), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_1612), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4427 (.Q (
                         modgen_ram_ix167_a_248__dup_1613), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_1613), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4431 (.Q (
                         modgen_ram_ix167_a_247__dup_1614), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_1614), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4435 (.Q (
                         modgen_ram_ix167_a_246__dup_1615), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_1615), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4439 (.Q (
                         modgen_ram_ix167_a_245__dup_1616), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_1616), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4443 (.Q (
                         modgen_ram_ix167_a_244__dup_1617), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_1617), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4447 (.Q (
                         modgen_ram_ix167_a_243__dup_1618), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_1618), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4451 (.Q (
                         modgen_ram_ix167_a_242__dup_1619), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_1619), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4455 (.Q (
                         modgen_ram_ix167_a_241__dup_1620), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_1620), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4459 (.Q (
                         modgen_ram_ix167_a_240__dup_1621), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_1621), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4463 (.Q (
                         modgen_ram_ix167_a_239__dup_1622), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_1622), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4467 (.Q (
                         modgen_ram_ix167_a_238__dup_1623), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_1623), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4471 (.Q (
                         modgen_ram_ix167_a_237__dup_1624), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_1624), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4475 (.Q (
                         modgen_ram_ix167_a_236__dup_1625), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_1625), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4479 (.Q (
                         modgen_ram_ix167_a_235__dup_1626), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_1626), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4483 (.Q (
                         modgen_ram_ix167_a_234__dup_1627), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_1627), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4487 (.Q (
                         modgen_ram_ix167_a_233__dup_1628), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_1628), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4491 (.Q (
                         modgen_ram_ix167_a_232__dup_1629), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_1629), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4495 (.Q (
                         modgen_ram_ix167_a_231__dup_1630), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_1630), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4499 (.Q (
                         modgen_ram_ix167_a_230__dup_1631), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_1631), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4503 (.Q (
                         modgen_ram_ix167_a_229__dup_1632), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_1632), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4507 (.Q (
                         modgen_ram_ix167_a_228__dup_1633), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_1633), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4511 (.Q (
                         modgen_ram_ix167_a_227__dup_1634), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_1634), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4515 (.Q (
                         modgen_ram_ix167_a_226__dup_1635), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_1635), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4519 (.Q (
                         modgen_ram_ix167_a_225__dup_1636), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_1636), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4523 (.Q (
                         modgen_ram_ix167_a_224__dup_1637), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_1637), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4527 (.Q (
                         modgen_ram_ix167_a_223__dup_1638), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_1638), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4531 (.Q (
                         modgen_ram_ix167_a_222__dup_1639), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_1639), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4535 (.Q (
                         modgen_ram_ix167_a_221__dup_1640), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_1640), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4539 (.Q (
                         modgen_ram_ix167_a_220__dup_1641), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_1641), .SN (nx28499)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4543 (.Q (
                         modgen_ram_ix167_a_219__dup_1642), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_1642), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4547 (.Q (
                         modgen_ram_ix167_a_218__dup_1643), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_1643), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4551 (.Q (
                         modgen_ram_ix167_a_217__dup_1644), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_1644), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4555 (.Q (
                         modgen_ram_ix167_a_216__dup_1645), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_1645), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4559 (.Q (
                         modgen_ram_ix167_a_215__dup_1646), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_1646), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4563 (.Q (
                         modgen_ram_ix167_a_214__dup_1647), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_1647), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4567 (.Q (
                         modgen_ram_ix167_a_213__dup_1648), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_1648), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4571 (.Q (
                         modgen_ram_ix167_a_212__dup_1649), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_1649), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4575 (.Q (
                         modgen_ram_ix167_a_211__dup_1650), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_1650), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4579 (.Q (
                         modgen_ram_ix167_a_210__dup_1651), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_1651), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4583 (.Q (
                         modgen_ram_ix167_a_209__dup_1652), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_1652), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4587 (.Q (
                         modgen_ram_ix167_a_208__dup_1653), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_1653), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4591 (.Q (
                         modgen_ram_ix167_a_207__dup_1654), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_1654), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4595 (.Q (
                         modgen_ram_ix167_a_206__dup_1655), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_1655), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4599 (.Q (
                         modgen_ram_ix167_a_205__dup_1656), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_1656), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4603 (.Q (
                         modgen_ram_ix167_a_204__dup_1657), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_1657), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4607 (.Q (
                         modgen_ram_ix167_a_203__dup_1658), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_1658), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4611 (.Q (
                         modgen_ram_ix167_a_202__dup_1659), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_1659), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4615 (.Q (
                         modgen_ram_ix167_a_201__dup_1660), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_1660), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4619 (.Q (
                         modgen_ram_ix167_a_200__dup_1661), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_1661), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4623 (.Q (
                         modgen_ram_ix167_a_199__dup_1662), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_1662), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4627 (.Q (
                         modgen_ram_ix167_a_198__dup_1663), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_1663), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4631 (.Q (
                         modgen_ram_ix167_a_197__dup_1664), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_1664), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4635 (.Q (
                         modgen_ram_ix167_a_196__dup_1665), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_1665), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4639 (.Q (
                         modgen_ram_ix167_a_195__dup_1666), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_1666), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4643 (.Q (
                         modgen_ram_ix167_a_194__dup_1667), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_1667), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4647 (.Q (
                         modgen_ram_ix167_a_193__dup_1668), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_1668), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4651 (.Q (
                         modgen_ram_ix167_a_192__dup_1669), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_1669), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4655 (.Q (
                         modgen_ram_ix167_a_191__dup_1670), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_1670), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4659 (.Q (
                         modgen_ram_ix167_a_190__dup_1671), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_1671), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4663 (.Q (
                         modgen_ram_ix167_a_189__dup_1672), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_1672), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4667 (.Q (
                         modgen_ram_ix167_a_188__dup_1673), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_1673), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4671 (.Q (
                         modgen_ram_ix167_a_187__dup_1674), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_1674), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4675 (.Q (
                         modgen_ram_ix167_a_186__dup_1675), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_1675), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4679 (.Q (
                         modgen_ram_ix167_a_185__dup_1676), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_1676), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4683 (.Q (
                         modgen_ram_ix167_a_184__dup_1677), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_1677), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4687 (.Q (
                         modgen_ram_ix167_a_183__dup_1678), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_1678), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4691 (.Q (
                         modgen_ram_ix167_a_182__dup_1679), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_1679), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4695 (.Q (
                         modgen_ram_ix167_a_181__dup_1680), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_1680), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4699 (.Q (
                         modgen_ram_ix167_a_180__dup_1681), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_1681), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4703 (.Q (
                         modgen_ram_ix167_a_179__dup_1682), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_1682), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4707 (.Q (
                         modgen_ram_ix167_a_178__dup_1683), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_1683), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4711 (.Q (
                         modgen_ram_ix167_a_177__dup_1684), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_1684), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4715 (.Q (
                         modgen_ram_ix167_a_176__dup_1685), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_1685), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4719 (.Q (
                         modgen_ram_ix167_a_175__dup_1686), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_1686), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4723 (.Q (
                         modgen_ram_ix167_a_174__dup_1687), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_1687), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4727 (.Q (
                         modgen_ram_ix167_a_173__dup_1688), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_1688), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4731 (.Q (
                         modgen_ram_ix167_a_172__dup_1689), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_1689), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4735 (.Q (
                         modgen_ram_ix167_a_171__dup_1690), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_1690), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4739 (.Q (
                         modgen_ram_ix167_a_170__dup_1691), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_1691), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4743 (.Q (
                         modgen_ram_ix167_a_169__dup_1692), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_1692), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4747 (.Q (
                         modgen_ram_ix167_a_168__dup_1693), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_1693), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4751 (.Q (
                         modgen_ram_ix167_a_167__dup_1694), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_1694), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4755 (.Q (
                         modgen_ram_ix167_a_166__dup_1695), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_1695), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4759 (.Q (
                         modgen_ram_ix167_a_165__dup_1696), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_1696), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4763 (.Q (
                         modgen_ram_ix167_a_164__dup_1697), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_1697), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4767 (.Q (
                         modgen_ram_ix167_a_163__dup_1698), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_1698), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4771 (.Q (
                         modgen_ram_ix167_a_162__dup_1699), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_1699), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4775 (.Q (
                         modgen_ram_ix167_a_161__dup_1700), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_1700), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4779 (.Q (
                         modgen_ram_ix167_a_160__dup_1701), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_1701), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4783 (.Q (
                         modgen_ram_ix167_a_159__dup_1702), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_1702), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4787 (.Q (
                         modgen_ram_ix167_a_158__dup_1703), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_1703), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4791 (.Q (
                         modgen_ram_ix167_a_157__dup_1704), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_1704), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4795 (.Q (
                         modgen_ram_ix167_a_156__dup_1705), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_1705), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4799 (.Q (
                         modgen_ram_ix167_a_155__dup_1706), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_1706), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4803 (.Q (
                         modgen_ram_ix167_a_154__dup_1707), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_1707), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4807 (.Q (
                         modgen_ram_ix167_a_153__dup_1708), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_1708), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4811 (.Q (
                         modgen_ram_ix167_a_152__dup_1709), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_1709), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4815 (.Q (
                         modgen_ram_ix167_a_151__dup_1710), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_1710), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4819 (.Q (
                         modgen_ram_ix167_a_150__dup_1711), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_1711), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4823 (.Q (
                         modgen_ram_ix167_a_149__dup_1712), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_1712), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4827 (.Q (
                         modgen_ram_ix167_a_148__dup_1713), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_1713), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4831 (.Q (
                         modgen_ram_ix167_a_147__dup_1714), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_1714), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4835 (.Q (
                         modgen_ram_ix167_a_146__dup_1715), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_1715), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4839 (.Q (
                         modgen_ram_ix167_a_145__dup_1716), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_1716), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4843 (.Q (
                         modgen_ram_ix167_a_144__dup_1717), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_1717), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4847 (.Q (
                         modgen_ram_ix167_a_143__dup_1718), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_1718), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4851 (.Q (
                         modgen_ram_ix167_a_142__dup_1719), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_1719), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4855 (.Q (
                         modgen_ram_ix167_a_141__dup_1720), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_1720), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4859 (.Q (
                         modgen_ram_ix167_a_140__dup_1721), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_1721), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4863 (.Q (
                         modgen_ram_ix167_a_139__dup_1722), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_1722), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4867 (.Q (
                         modgen_ram_ix167_a_138__dup_1723), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_1723), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4871 (.Q (
                         modgen_ram_ix167_a_137__dup_1724), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_1724), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4875 (.Q (
                         modgen_ram_ix167_a_136__dup_1725), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_1725), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4879 (.Q (
                         modgen_ram_ix167_a_135__dup_1726), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_1726), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4883 (.Q (
                         modgen_ram_ix167_a_134__dup_1727), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_1727), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4887 (.Q (
                         modgen_ram_ix167_a_133__dup_1728), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_1728), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4891 (.Q (
                         modgen_ram_ix167_a_132__dup_1729), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_1729), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4895 (.Q (
                         modgen_ram_ix167_a_131__dup_1730), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_1730), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4899 (.Q (
                         modgen_ram_ix167_a_130__dup_1731), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_1731), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4903 (.Q (
                         modgen_ram_ix167_a_129__dup_1732), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_1732), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4907 (.Q (
                         modgen_ram_ix167_a_128__dup_1733), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_1733), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4911 (.Q (
                         modgen_ram_ix167_a_127__dup_1734), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_1734), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4915 (.Q (
                         modgen_ram_ix167_a_126__dup_1735), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_1735), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4919 (.Q (
                         modgen_ram_ix167_a_125__dup_1736), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_1736), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4923 (.Q (
                         modgen_ram_ix167_a_124__dup_1737), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_1737), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4927 (.Q (
                         modgen_ram_ix167_a_123__dup_1738), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_1738), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4931 (.Q (
                         modgen_ram_ix167_a_122__dup_1739), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_1739), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4935 (.Q (
                         modgen_ram_ix167_a_121__dup_1740), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_1740), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4939 (.Q (
                         modgen_ram_ix167_a_120__dup_1741), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_1741), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4943 (.Q (
                         modgen_ram_ix167_a_119__dup_1742), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_1742), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4947 (.Q (
                         modgen_ram_ix167_a_118__dup_1743), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_1743), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4951 (.Q (
                         modgen_ram_ix167_a_117__dup_1744), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_1744), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4955 (.Q (
                         modgen_ram_ix167_a_116__dup_1745), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_1745), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4959 (.Q (
                         modgen_ram_ix167_a_115__dup_1746), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_1746), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4963 (.Q (
                         modgen_ram_ix167_a_114__dup_1747), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_1747), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4967 (.Q (
                         modgen_ram_ix167_a_113__dup_1748), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_1748), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4971 (.Q (
                         modgen_ram_ix167_a_112__dup_1749), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_1749), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4975 (.Q (
                         modgen_ram_ix167_a_111__dup_1750), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_1750), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4979 (.Q (
                         modgen_ram_ix167_a_110__dup_1751), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_1751), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4983 (.Q (
                         modgen_ram_ix167_a_109__dup_1752), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_1752), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4987 (.Q (
                         modgen_ram_ix167_a_108__dup_1753), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_1753), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4991 (.Q (
                         modgen_ram_ix167_a_107__dup_1754), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_1754), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4995 (.Q (
                         modgen_ram_ix167_a_106__dup_1755), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_1755), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix4999 (.Q (
                         modgen_ram_ix167_a_105__dup_1756), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_1756), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5003 (.Q (
                         modgen_ram_ix167_a_104__dup_1757), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_1757), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5007 (.Q (
                         modgen_ram_ix167_a_103__dup_1758), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_1758), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5011 (.Q (
                         modgen_ram_ix167_a_102__dup_1759), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_1759), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5015 (.Q (
                         modgen_ram_ix167_a_101__dup_1760), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_1760), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5019 (.Q (
                         modgen_ram_ix167_a_100__dup_1761), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_1761), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5023 (.Q (
                         modgen_ram_ix167_a_99__dup_1762), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_1762), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5027 (.Q (
                         modgen_ram_ix167_a_98__dup_1763), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_1763), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5031 (.Q (
                         modgen_ram_ix167_a_97__dup_1764), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_1764), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5035 (.Q (
                         modgen_ram_ix167_a_96__dup_1765), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_1765), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5039 (.Q (
                         modgen_ram_ix167_a_95__dup_1766), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_1766), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5043 (.Q (
                         modgen_ram_ix167_a_94__dup_1767), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_1767), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5047 (.Q (
                         modgen_ram_ix167_a_93__dup_1768), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_1768), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5051 (.Q (
                         modgen_ram_ix167_a_92__dup_1769), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_1769), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5055 (.Q (
                         modgen_ram_ix167_a_91__dup_1770), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_1770), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5059 (.Q (
                         modgen_ram_ix167_a_90__dup_1771), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_1771), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5063 (.Q (
                         modgen_ram_ix167_a_89__dup_1772), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_1772), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5067 (.Q (
                         modgen_ram_ix167_a_88__dup_1773), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_1773), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5071 (.Q (
                         modgen_ram_ix167_a_87__dup_1774), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_1774), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5075 (.Q (
                         modgen_ram_ix167_a_86__dup_1775), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_1775), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5079 (.Q (
                         modgen_ram_ix167_a_85__dup_1776), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_1776), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5083 (.Q (
                         modgen_ram_ix167_a_84__dup_1777), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_1777), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5087 (.Q (
                         modgen_ram_ix167_a_83__dup_1778), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_1778), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5091 (.Q (
                         modgen_ram_ix167_a_82__dup_1779), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_1779), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5095 (.Q (
                         modgen_ram_ix167_a_81__dup_1780), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_1780), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5099 (.Q (
                         modgen_ram_ix167_a_80__dup_1781), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_1781), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5103 (.Q (
                         modgen_ram_ix167_a_79__dup_1782), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_1782), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5107 (.Q (
                         modgen_ram_ix167_a_78__dup_1783), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_1783), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5111 (.Q (
                         modgen_ram_ix167_a_77__dup_1784), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_1784), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5115 (.Q (
                         modgen_ram_ix167_a_76__dup_1785), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_1785), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5119 (.Q (
                         modgen_ram_ix167_a_75__dup_1786), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_1786), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5123 (.Q (
                         modgen_ram_ix167_a_74__dup_1787), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_1787), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5127 (.Q (
                         modgen_ram_ix167_a_73__dup_1788), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_1788), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5131 (.Q (
                         modgen_ram_ix167_a_72__dup_1789), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_1789), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5135 (.Q (
                         modgen_ram_ix167_a_71__dup_1790), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_1790), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5139 (.Q (
                         modgen_ram_ix167_a_70__dup_1791), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_1791), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5143 (.Q (
                         modgen_ram_ix167_a_69__dup_1792), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_1792), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5147 (.Q (
                         modgen_ram_ix167_a_68__dup_1793), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_1793), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5151 (.Q (
                         modgen_ram_ix167_a_67__dup_1794), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_1794), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5155 (.Q (
                         modgen_ram_ix167_a_66__dup_1795), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_1795), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5159 (.Q (
                         modgen_ram_ix167_a_65__dup_1796), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_1796), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5163 (.Q (
                         modgen_ram_ix167_a_64__dup_1797), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_1797), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5167 (.Q (
                         modgen_ram_ix167_a_63__dup_1798), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_1798), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5171 (.Q (
                         modgen_ram_ix167_a_62__dup_1799), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_1799), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5175 (.Q (
                         modgen_ram_ix167_a_61__dup_1800), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_1800), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5179 (.Q (
                         modgen_ram_ix167_a_60__dup_1801), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_1801), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5183 (.Q (
                         modgen_ram_ix167_a_59__dup_1802), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_1802), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5187 (.Q (
                         modgen_ram_ix167_a_58__dup_1803), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_1803), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5191 (.Q (
                         modgen_ram_ix167_a_57__dup_1804), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_1804), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5195 (.Q (
                         modgen_ram_ix167_a_56__dup_1805), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_1805), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5199 (.Q (
                         modgen_ram_ix167_a_55__dup_1806), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_1806), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5203 (.Q (
                         modgen_ram_ix167_a_54__dup_1807), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_1807), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5207 (.Q (
                         modgen_ram_ix167_a_53__dup_1808), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_1808), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5211 (.Q (
                         modgen_ram_ix167_a_52__dup_1809), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_1809), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5215 (.Q (
                         modgen_ram_ix167_a_51__dup_1810), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_1810), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5219 (.Q (
                         modgen_ram_ix167_a_50__dup_1811), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_1811), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5223 (.Q (
                         modgen_ram_ix167_a_49__dup_1812), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_1812), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5227 (.Q (
                         modgen_ram_ix167_a_48__dup_1813), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_1813), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5231 (.Q (
                         modgen_ram_ix167_a_47__dup_1814), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_1814), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5235 (.Q (
                         modgen_ram_ix167_a_46__dup_1815), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_1815), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5239 (.Q (
                         modgen_ram_ix167_a_45__dup_1816), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_1816), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5243 (.Q (
                         modgen_ram_ix167_a_44__dup_1817), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_1817), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5247 (.Q (
                         modgen_ram_ix167_a_43__dup_1818), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_1818), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5251 (.Q (
                         modgen_ram_ix167_a_42__dup_1819), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_1819), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5255 (.Q (
                         modgen_ram_ix167_a_41__dup_1820), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_1820), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5259 (.Q (
                         modgen_ram_ix167_a_40__dup_1821), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_1821), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5263 (.Q (
                         modgen_ram_ix167_a_39__dup_1822), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_1822), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5267 (.Q (
                         modgen_ram_ix167_a_38__dup_1823), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_1823), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5271 (.Q (
                         modgen_ram_ix167_a_37__dup_1824), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_1824), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5275 (.Q (
                         modgen_ram_ix167_a_36__dup_1825), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_1825), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5279 (.Q (
                         modgen_ram_ix167_a_35__dup_1826), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_1826), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5283 (.Q (
                         modgen_ram_ix167_a_34__dup_1827), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_1827), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5287 (.Q (
                         modgen_ram_ix167_a_33__dup_1828), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_1828), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5291 (.Q (
                         modgen_ram_ix167_a_32__dup_1829), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_1829), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5295 (.Q (
                         modgen_ram_ix167_a_31__dup_1830), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_1830), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5299 (.Q (
                         modgen_ram_ix167_a_30__dup_1831), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_1831), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5303 (.Q (
                         modgen_ram_ix167_a_29__dup_1832), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_1832), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5307 (.Q (
                         modgen_ram_ix167_a_28__dup_1833), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_1833), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5311 (.Q (
                         modgen_ram_ix167_a_27__dup_1834), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_1834), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5315 (.Q (
                         modgen_ram_ix167_a_26__dup_1835), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_1835), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5319 (.Q (
                         modgen_ram_ix167_a_25__dup_1836), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_1836), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5323 (.Q (
                         modgen_ram_ix167_a_24__dup_1837), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_1837), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5327 (.Q (
                         modgen_ram_ix167_a_23__dup_1838), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_1838), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5331 (.Q (
                         modgen_ram_ix167_a_22__dup_1839), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_1839), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5335 (.Q (
                         modgen_ram_ix167_a_21__dup_1840), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_1840), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5339 (.Q (
                         modgen_ram_ix167_a_20__dup_1841), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_1841), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5343 (.Q (
                         modgen_ram_ix167_a_19__dup_1842), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_1842), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5347 (.Q (
                         modgen_ram_ix167_a_18__dup_1843), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_1843), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5351 (.Q (
                         modgen_ram_ix167_a_17__dup_1844), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_1844), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5355 (.Q (
                         modgen_ram_ix167_a_16__dup_1845), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_1845), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5359 (.Q (
                         modgen_ram_ix167_a_15__dup_1846), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_1846), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5363 (.Q (
                         modgen_ram_ix167_a_14__dup_1847), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_1847), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5367 (.Q (
                         modgen_ram_ix167_a_13__dup_1848), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_1848), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5371 (.Q (
                         modgen_ram_ix167_a_12__dup_1849), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_1849), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5375 (.Q (
                         modgen_ram_ix167_a_11__dup_1850), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_1850), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5379 (.Q (
                         modgen_ram_ix167_a_10__dup_1851), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_1851), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5383 (.Q (
                         modgen_ram_ix167_a_9__dup_1852), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_1852), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5387 (.Q (
                         modgen_ram_ix167_a_8__dup_1853), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_1853), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5391 (.Q (
                         modgen_ram_ix167_a_7__dup_1854), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_1854), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5395 (.Q (
                         modgen_ram_ix167_a_6__dup_1855), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_1855), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5399 (.Q (
                         modgen_ram_ix167_a_5__dup_1856), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_1856), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5403 (.Q (
                         modgen_ram_ix167_a_4__dup_1857), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_1857), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5407 (.Q (
                         modgen_ram_ix167_a_3__dup_1858), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_1858), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5411 (.Q (
                         modgen_ram_ix167_a_2__dup_1859), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_1859), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5415 (.Q (
                         modgen_ram_ix167_a_1__dup_1860), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_1860), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5419 (.Q (
                         modgen_ram_ix167_a_0__dup_1861), .CK (wb_clk_i), .D (
                         nx28517), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_1861), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5424 (.Q (
                         modgen_ram_ix167_a_255__dup_1870), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_1870), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5428 (.Q (
                         modgen_ram_ix167_a_254__dup_1871), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_1871), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5432 (.Q (
                         modgen_ram_ix167_a_253__dup_1872), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_1872), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5436 (.Q (
                         modgen_ram_ix167_a_252__dup_1873), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_1873), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5440 (.Q (
                         modgen_ram_ix167_a_251__dup_1874), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_1874), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5444 (.Q (
                         modgen_ram_ix167_a_250__dup_1875), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_1875), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5448 (.Q (
                         modgen_ram_ix167_a_249__dup_1876), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_1876), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5452 (.Q (
                         modgen_ram_ix167_a_248__dup_1877), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_1877), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5456 (.Q (
                         modgen_ram_ix167_a_247__dup_1878), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_1878), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5460 (.Q (
                         modgen_ram_ix167_a_246__dup_1879), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_1879), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5464 (.Q (
                         modgen_ram_ix167_a_245__dup_1880), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_1880), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5468 (.Q (
                         modgen_ram_ix167_a_244__dup_1881), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_1881), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5472 (.Q (
                         modgen_ram_ix167_a_243__dup_1882), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_1882), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5476 (.Q (
                         modgen_ram_ix167_a_242__dup_1883), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_1883), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5480 (.Q (
                         modgen_ram_ix167_a_241__dup_1884), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_1884), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5484 (.Q (
                         modgen_ram_ix167_a_240__dup_1885), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_1885), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5488 (.Q (
                         modgen_ram_ix167_a_239__dup_1886), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_1886), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5492 (.Q (
                         modgen_ram_ix167_a_238__dup_1887), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_1887), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5496 (.Q (
                         modgen_ram_ix167_a_237__dup_1888), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_1888), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5500 (.Q (
                         modgen_ram_ix167_a_236__dup_1889), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_1889), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5504 (.Q (
                         modgen_ram_ix167_a_235__dup_1890), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_1890), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5508 (.Q (
                         modgen_ram_ix167_a_234__dup_1891), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_1891), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5512 (.Q (
                         modgen_ram_ix167_a_233__dup_1892), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_1892), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5516 (.Q (
                         modgen_ram_ix167_a_232__dup_1893), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_1893), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5520 (.Q (
                         modgen_ram_ix167_a_231__dup_1894), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_1894), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5524 (.Q (
                         modgen_ram_ix167_a_230__dup_1895), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_1895), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5528 (.Q (
                         modgen_ram_ix167_a_229__dup_1896), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_1896), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5532 (.Q (
                         modgen_ram_ix167_a_228__dup_1897), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_1897), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5536 (.Q (
                         modgen_ram_ix167_a_227__dup_1898), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_1898), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5540 (.Q (
                         modgen_ram_ix167_a_226__dup_1899), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_1899), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5544 (.Q (
                         modgen_ram_ix167_a_225__dup_1900), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_1900), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5548 (.Q (
                         modgen_ram_ix167_a_224__dup_1901), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_1901), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5552 (.Q (
                         modgen_ram_ix167_a_223__dup_1902), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_1902), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5556 (.Q (
                         modgen_ram_ix167_a_222__dup_1903), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_1903), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5560 (.Q (
                         modgen_ram_ix167_a_221__dup_1904), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_1904), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5564 (.Q (
                         modgen_ram_ix167_a_220__dup_1905), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_1905), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5568 (.Q (
                         modgen_ram_ix167_a_219__dup_1906), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_1906), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5572 (.Q (
                         modgen_ram_ix167_a_218__dup_1907), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_1907), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5576 (.Q (
                         modgen_ram_ix167_a_217__dup_1908), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_1908), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5580 (.Q (
                         modgen_ram_ix167_a_216__dup_1909), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_1909), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5584 (.Q (
                         modgen_ram_ix167_a_215__dup_1910), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_1910), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5588 (.Q (
                         modgen_ram_ix167_a_214__dup_1911), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_1911), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5592 (.Q (
                         modgen_ram_ix167_a_213__dup_1912), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_1912), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5596 (.Q (
                         modgen_ram_ix167_a_212__dup_1913), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_1913), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5600 (.Q (
                         modgen_ram_ix167_a_211__dup_1914), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_1914), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5604 (.Q (
                         modgen_ram_ix167_a_210__dup_1915), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_1915), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5608 (.Q (
                         modgen_ram_ix167_a_209__dup_1916), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_1916), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5612 (.Q (
                         modgen_ram_ix167_a_208__dup_1917), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_1917), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5616 (.Q (
                         modgen_ram_ix167_a_207__dup_1918), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_1918), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5620 (.Q (
                         modgen_ram_ix167_a_206__dup_1919), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_1919), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5624 (.Q (
                         modgen_ram_ix167_a_205__dup_1920), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_1920), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5628 (.Q (
                         modgen_ram_ix167_a_204__dup_1921), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_1921), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5632 (.Q (
                         modgen_ram_ix167_a_203__dup_1922), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_1922), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5636 (.Q (
                         modgen_ram_ix167_a_202__dup_1923), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_1923), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5640 (.Q (
                         modgen_ram_ix167_a_201__dup_1924), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_1924), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5644 (.Q (
                         modgen_ram_ix167_a_200__dup_1925), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_1925), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5648 (.Q (
                         modgen_ram_ix167_a_199__dup_1926), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_1926), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5652 (.Q (
                         modgen_ram_ix167_a_198__dup_1927), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_1927), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5656 (.Q (
                         modgen_ram_ix167_a_197__dup_1928), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_1928), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5660 (.Q (
                         modgen_ram_ix167_a_196__dup_1929), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_1929), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5664 (.Q (
                         modgen_ram_ix167_a_195__dup_1930), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_1930), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5668 (.Q (
                         modgen_ram_ix167_a_194__dup_1931), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_1931), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5672 (.Q (
                         modgen_ram_ix167_a_193__dup_1932), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_1932), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5676 (.Q (
                         modgen_ram_ix167_a_192__dup_1933), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_1933), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5680 (.Q (
                         modgen_ram_ix167_a_191__dup_1934), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_1934), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5684 (.Q (
                         modgen_ram_ix167_a_190__dup_1935), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_1935), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5688 (.Q (
                         modgen_ram_ix167_a_189__dup_1936), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_1936), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5692 (.Q (
                         modgen_ram_ix167_a_188__dup_1937), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_1937), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5696 (.Q (
                         modgen_ram_ix167_a_187__dup_1938), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_1938), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5700 (.Q (
                         modgen_ram_ix167_a_186__dup_1939), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_1939), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5704 (.Q (
                         modgen_ram_ix167_a_185__dup_1940), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_1940), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5708 (.Q (
                         modgen_ram_ix167_a_184__dup_1941), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_1941), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5712 (.Q (
                         modgen_ram_ix167_a_183__dup_1942), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_1942), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5716 (.Q (
                         modgen_ram_ix167_a_182__dup_1943), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_1943), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5720 (.Q (
                         modgen_ram_ix167_a_181__dup_1944), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_1944), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5724 (.Q (
                         modgen_ram_ix167_a_180__dup_1945), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_1945), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5728 (.Q (
                         modgen_ram_ix167_a_179__dup_1946), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_1946), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5732 (.Q (
                         modgen_ram_ix167_a_178__dup_1947), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_1947), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5736 (.Q (
                         modgen_ram_ix167_a_177__dup_1948), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_1948), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5740 (.Q (
                         modgen_ram_ix167_a_176__dup_1949), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_1949), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5744 (.Q (
                         modgen_ram_ix167_a_175__dup_1950), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_1950), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5748 (.Q (
                         modgen_ram_ix167_a_174__dup_1951), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_1951), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5752 (.Q (
                         modgen_ram_ix167_a_173__dup_1952), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_1952), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5756 (.Q (
                         modgen_ram_ix167_a_172__dup_1953), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_1953), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5760 (.Q (
                         modgen_ram_ix167_a_171__dup_1954), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_1954), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5764 (.Q (
                         modgen_ram_ix167_a_170__dup_1955), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_1955), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5768 (.Q (
                         modgen_ram_ix167_a_169__dup_1956), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_1956), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5772 (.Q (
                         modgen_ram_ix167_a_168__dup_1957), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_1957), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5776 (.Q (
                         modgen_ram_ix167_a_167__dup_1958), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_1958), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5780 (.Q (
                         modgen_ram_ix167_a_166__dup_1959), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_1959), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5784 (.Q (
                         modgen_ram_ix167_a_165__dup_1960), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_1960), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5788 (.Q (
                         modgen_ram_ix167_a_164__dup_1961), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_1961), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5792 (.Q (
                         modgen_ram_ix167_a_163__dup_1962), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_1962), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5796 (.Q (
                         modgen_ram_ix167_a_162__dup_1963), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_1963), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5800 (.Q (
                         modgen_ram_ix167_a_161__dup_1964), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_1964), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5804 (.Q (
                         modgen_ram_ix167_a_160__dup_1965), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_1965), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5808 (.Q (
                         modgen_ram_ix167_a_159__dup_1966), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_1966), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5812 (.Q (
                         modgen_ram_ix167_a_158__dup_1967), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_1967), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5816 (.Q (
                         modgen_ram_ix167_a_157__dup_1968), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_1968), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5820 (.Q (
                         modgen_ram_ix167_a_156__dup_1969), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_1969), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5824 (.Q (
                         modgen_ram_ix167_a_155__dup_1970), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_1970), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5828 (.Q (
                         modgen_ram_ix167_a_154__dup_1971), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_1971), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5832 (.Q (
                         modgen_ram_ix167_a_153__dup_1972), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_1972), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5836 (.Q (
                         modgen_ram_ix167_a_152__dup_1973), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_1973), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5840 (.Q (
                         modgen_ram_ix167_a_151__dup_1974), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_1974), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5844 (.Q (
                         modgen_ram_ix167_a_150__dup_1975), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_1975), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5848 (.Q (
                         modgen_ram_ix167_a_149__dup_1976), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_1976), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5852 (.Q (
                         modgen_ram_ix167_a_148__dup_1977), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_1977), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5856 (.Q (
                         modgen_ram_ix167_a_147__dup_1978), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_1978), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5860 (.Q (
                         modgen_ram_ix167_a_146__dup_1979), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_1979), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5864 (.Q (
                         modgen_ram_ix167_a_145__dup_1980), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_1980), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5868 (.Q (
                         modgen_ram_ix167_a_144__dup_1981), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_1981), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5872 (.Q (
                         modgen_ram_ix167_a_143__dup_1982), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_1982), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5876 (.Q (
                         modgen_ram_ix167_a_142__dup_1983), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_1983), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5880 (.Q (
                         modgen_ram_ix167_a_141__dup_1984), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_1984), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5884 (.Q (
                         modgen_ram_ix167_a_140__dup_1985), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_1985), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5888 (.Q (
                         modgen_ram_ix167_a_139__dup_1986), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_1986), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5892 (.Q (
                         modgen_ram_ix167_a_138__dup_1987), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_1987), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5896 (.Q (
                         modgen_ram_ix167_a_137__dup_1988), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_1988), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5900 (.Q (
                         modgen_ram_ix167_a_136__dup_1989), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_1989), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5904 (.Q (
                         modgen_ram_ix167_a_135__dup_1990), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_1990), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5908 (.Q (
                         modgen_ram_ix167_a_134__dup_1991), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_1991), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5912 (.Q (
                         modgen_ram_ix167_a_133__dup_1992), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_1992), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5916 (.Q (
                         modgen_ram_ix167_a_132__dup_1993), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_1993), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5920 (.Q (
                         modgen_ram_ix167_a_131__dup_1994), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_1994), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5924 (.Q (
                         modgen_ram_ix167_a_130__dup_1995), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_1995), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5928 (.Q (
                         modgen_ram_ix167_a_129__dup_1996), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_1996), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5932 (.Q (
                         modgen_ram_ix167_a_128__dup_1997), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_1997), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5936 (.Q (
                         modgen_ram_ix167_a_127__dup_1998), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_1998), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5940 (.Q (
                         modgen_ram_ix167_a_126__dup_1999), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_1999), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5944 (.Q (
                         modgen_ram_ix167_a_125__dup_2000), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_2000), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5948 (.Q (
                         modgen_ram_ix167_a_124__dup_2001), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_2001), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5952 (.Q (
                         modgen_ram_ix167_a_123__dup_2002), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_2002), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5956 (.Q (
                         modgen_ram_ix167_a_122__dup_2003), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_2003), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5960 (.Q (
                         modgen_ram_ix167_a_121__dup_2004), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_2004), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5964 (.Q (
                         modgen_ram_ix167_a_120__dup_2005), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_2005), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5968 (.Q (
                         modgen_ram_ix167_a_119__dup_2006), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_2006), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5972 (.Q (
                         modgen_ram_ix167_a_118__dup_2007), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_2007), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5976 (.Q (
                         modgen_ram_ix167_a_117__dup_2008), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_2008), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5980 (.Q (
                         modgen_ram_ix167_a_116__dup_2009), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_2009), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5984 (.Q (
                         modgen_ram_ix167_a_115__dup_2010), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_2010), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5988 (.Q (
                         modgen_ram_ix167_a_114__dup_2011), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_2011), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5992 (.Q (
                         modgen_ram_ix167_a_113__dup_2012), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_2012), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix5996 (.Q (
                         modgen_ram_ix167_a_112__dup_2013), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_2013), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6000 (.Q (
                         modgen_ram_ix167_a_111__dup_2014), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_2014), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6004 (.Q (
                         modgen_ram_ix167_a_110__dup_2015), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_2015), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6008 (.Q (
                         modgen_ram_ix167_a_109__dup_2016), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_2016), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6012 (.Q (
                         modgen_ram_ix167_a_108__dup_2017), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_2017), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6016 (.Q (
                         modgen_ram_ix167_a_107__dup_2018), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_2018), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6020 (.Q (
                         modgen_ram_ix167_a_106__dup_2019), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_2019), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6024 (.Q (
                         modgen_ram_ix167_a_105__dup_2020), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_2020), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6028 (.Q (
                         modgen_ram_ix167_a_104__dup_2021), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_2021), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6032 (.Q (
                         modgen_ram_ix167_a_103__dup_2022), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_2022), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6036 (.Q (
                         modgen_ram_ix167_a_102__dup_2023), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_2023), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6040 (.Q (
                         modgen_ram_ix167_a_101__dup_2024), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_2024), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6044 (.Q (
                         modgen_ram_ix167_a_100__dup_2025), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_2025), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6048 (.Q (
                         modgen_ram_ix167_a_99__dup_2026), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_2026), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6052 (.Q (
                         modgen_ram_ix167_a_98__dup_2027), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_2027), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6056 (.Q (
                         modgen_ram_ix167_a_97__dup_2028), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_2028), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6060 (.Q (
                         modgen_ram_ix167_a_96__dup_2029), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_2029), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6064 (.Q (
                         modgen_ram_ix167_a_95__dup_2030), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_2030), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6068 (.Q (
                         modgen_ram_ix167_a_94__dup_2031), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_2031), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6072 (.Q (
                         modgen_ram_ix167_a_93__dup_2032), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_2032), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6076 (.Q (
                         modgen_ram_ix167_a_92__dup_2033), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_2033), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6080 (.Q (
                         modgen_ram_ix167_a_91__dup_2034), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_2034), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6084 (.Q (
                         modgen_ram_ix167_a_90__dup_2035), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_2035), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6088 (.Q (
                         modgen_ram_ix167_a_89__dup_2036), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_2036), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6092 (.Q (
                         modgen_ram_ix167_a_88__dup_2037), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_2037), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6096 (.Q (
                         modgen_ram_ix167_a_87__dup_2038), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_2038), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6100 (.Q (
                         modgen_ram_ix167_a_86__dup_2039), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_2039), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6104 (.Q (
                         modgen_ram_ix167_a_85__dup_2040), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_2040), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6108 (.Q (
                         modgen_ram_ix167_a_84__dup_2041), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_2041), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6112 (.Q (
                         modgen_ram_ix167_a_83__dup_2042), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_2042), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6116 (.Q (
                         modgen_ram_ix167_a_82__dup_2043), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_2043), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6120 (.Q (
                         modgen_ram_ix167_a_81__dup_2044), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_2044), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6124 (.Q (
                         modgen_ram_ix167_a_80__dup_2045), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_2045), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6128 (.Q (
                         modgen_ram_ix167_a_79__dup_2046), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_2046), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6132 (.Q (
                         modgen_ram_ix167_a_78__dup_2047), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_2047), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6136 (.Q (
                         modgen_ram_ix167_a_77__dup_2048), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_2048), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6140 (.Q (
                         modgen_ram_ix167_a_76__dup_2049), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_2049), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6144 (.Q (
                         modgen_ram_ix167_a_75__dup_2050), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_2050), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6148 (.Q (
                         modgen_ram_ix167_a_74__dup_2051), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_2051), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6152 (.Q (
                         modgen_ram_ix167_a_73__dup_2052), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_2052), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6156 (.Q (
                         modgen_ram_ix167_a_72__dup_2053), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_2053), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6160 (.Q (
                         modgen_ram_ix167_a_71__dup_2054), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_2054), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6164 (.Q (
                         modgen_ram_ix167_a_70__dup_2055), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_2055), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6168 (.Q (
                         modgen_ram_ix167_a_69__dup_2056), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_2056), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6172 (.Q (
                         modgen_ram_ix167_a_68__dup_2057), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_2057), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6176 (.Q (
                         modgen_ram_ix167_a_67__dup_2058), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_2058), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6180 (.Q (
                         modgen_ram_ix167_a_66__dup_2059), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_2059), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6184 (.Q (
                         modgen_ram_ix167_a_65__dup_2060), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_2060), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6188 (.Q (
                         modgen_ram_ix167_a_64__dup_2061), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_2061), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6192 (.Q (
                         modgen_ram_ix167_a_63__dup_2062), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_2062), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6196 (.Q (
                         modgen_ram_ix167_a_62__dup_2063), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_2063), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6200 (.Q (
                         modgen_ram_ix167_a_61__dup_2064), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_2064), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6204 (.Q (
                         modgen_ram_ix167_a_60__dup_2065), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_2065), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6208 (.Q (
                         modgen_ram_ix167_a_59__dup_2066), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_2066), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6212 (.Q (
                         modgen_ram_ix167_a_58__dup_2067), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_2067), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6216 (.Q (
                         modgen_ram_ix167_a_57__dup_2068), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_2068), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6220 (.Q (
                         modgen_ram_ix167_a_56__dup_2069), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_2069), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6224 (.Q (
                         modgen_ram_ix167_a_55__dup_2070), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_2070), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6228 (.Q (
                         modgen_ram_ix167_a_54__dup_2071), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_2071), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6232 (.Q (
                         modgen_ram_ix167_a_53__dup_2072), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_2072), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6236 (.Q (
                         modgen_ram_ix167_a_52__dup_2073), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_2073), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6240 (.Q (
                         modgen_ram_ix167_a_51__dup_2074), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_2074), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6244 (.Q (
                         modgen_ram_ix167_a_50__dup_2075), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_2075), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6248 (.Q (
                         modgen_ram_ix167_a_49__dup_2076), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_2076), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6252 (.Q (
                         modgen_ram_ix167_a_48__dup_2077), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_2077), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6256 (.Q (
                         modgen_ram_ix167_a_47__dup_2078), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_2078), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6260 (.Q (
                         modgen_ram_ix167_a_46__dup_2079), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_2079), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6264 (.Q (
                         modgen_ram_ix167_a_45__dup_2080), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_2080), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6268 (.Q (
                         modgen_ram_ix167_a_44__dup_2081), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_2081), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6272 (.Q (
                         modgen_ram_ix167_a_43__dup_2082), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_2082), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6276 (.Q (
                         modgen_ram_ix167_a_42__dup_2083), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_2083), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6280 (.Q (
                         modgen_ram_ix167_a_41__dup_2084), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_2084), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6284 (.Q (
                         modgen_ram_ix167_a_40__dup_2085), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_2085), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6288 (.Q (
                         modgen_ram_ix167_a_39__dup_2086), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_2086), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6292 (.Q (
                         modgen_ram_ix167_a_38__dup_2087), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_2087), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6296 (.Q (
                         modgen_ram_ix167_a_37__dup_2088), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_2088), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6300 (.Q (
                         modgen_ram_ix167_a_36__dup_2089), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_2089), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6304 (.Q (
                         modgen_ram_ix167_a_35__dup_2090), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_2090), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6308 (.Q (
                         modgen_ram_ix167_a_34__dup_2091), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_2091), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6312 (.Q (
                         modgen_ram_ix167_a_33__dup_2092), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_2092), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6316 (.Q (
                         modgen_ram_ix167_a_32__dup_2093), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_2093), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6320 (.Q (
                         modgen_ram_ix167_a_31__dup_2094), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_2094), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6324 (.Q (
                         modgen_ram_ix167_a_30__dup_2095), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_2095), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6328 (.Q (
                         modgen_ram_ix167_a_29__dup_2096), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_2096), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6332 (.Q (
                         modgen_ram_ix167_a_28__dup_2097), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_2097), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6336 (.Q (
                         modgen_ram_ix167_a_27__dup_2098), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_2098), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6340 (.Q (
                         modgen_ram_ix167_a_26__dup_2099), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_2099), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6344 (.Q (
                         modgen_ram_ix167_a_25__dup_2100), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_2100), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6348 (.Q (
                         modgen_ram_ix167_a_24__dup_2101), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_2101), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6352 (.Q (
                         modgen_ram_ix167_a_23__dup_2102), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_2102), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6356 (.Q (
                         modgen_ram_ix167_a_22__dup_2103), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_2103), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6360 (.Q (
                         modgen_ram_ix167_a_21__dup_2104), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_2104), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6364 (.Q (
                         modgen_ram_ix167_a_20__dup_2105), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_2105), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6368 (.Q (
                         modgen_ram_ix167_a_19__dup_2106), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_2106), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6372 (.Q (
                         modgen_ram_ix167_a_18__dup_2107), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_2107), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6376 (.Q (
                         modgen_ram_ix167_a_17__dup_2108), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_2108), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6380 (.Q (
                         modgen_ram_ix167_a_16__dup_2109), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_2109), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6384 (.Q (
                         modgen_ram_ix167_a_15__dup_2110), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_2110), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6388 (.Q (
                         modgen_ram_ix167_a_14__dup_2111), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_2111), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6392 (.Q (
                         modgen_ram_ix167_a_13__dup_2112), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_2112), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6396 (.Q (
                         modgen_ram_ix167_a_12__dup_2113), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_2113), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6400 (.Q (
                         modgen_ram_ix167_a_11__dup_2114), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_2114), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6404 (.Q (
                         modgen_ram_ix167_a_10__dup_2115), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_2115), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6408 (.Q (
                         modgen_ram_ix167_a_9__dup_2116), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_2116), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6412 (.Q (
                         modgen_ram_ix167_a_8__dup_2117), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_2117), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6416 (.Q (
                         modgen_ram_ix167_a_7__dup_2118), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_2118), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6420 (.Q (
                         modgen_ram_ix167_a_6__dup_2119), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_2119), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6424 (.Q (
                         modgen_ram_ix167_a_5__dup_2120), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_2120), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6428 (.Q (
                         modgen_ram_ix167_a_4__dup_2121), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_2121), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6432 (.Q (
                         modgen_ram_ix167_a_3__dup_2122), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_2122), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6436 (.Q (
                         modgen_ram_ix167_a_2__dup_2123), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_2123), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6440 (.Q (
                         modgen_ram_ix167_a_1__dup_2124), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_2124), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6444 (.Q (
                         modgen_ram_ix167_a_0__dup_2125), .CK (wb_clk_i), .D (
                         nx28519), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_2125), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6449 (.Q (
                         modgen_ram_ix167_a_255__dup_2134), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_2134), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6453 (.Q (
                         modgen_ram_ix167_a_254__dup_2135), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_2135), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6457 (.Q (
                         modgen_ram_ix167_a_253__dup_2136), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_2136), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6461 (.Q (
                         modgen_ram_ix167_a_252__dup_2137), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_2137), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6465 (.Q (
                         modgen_ram_ix167_a_251__dup_2138), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_2138), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6469 (.Q (
                         modgen_ram_ix167_a_250__dup_2139), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_2139), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6473 (.Q (
                         modgen_ram_ix167_a_249__dup_2140), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_2140), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6477 (.Q (
                         modgen_ram_ix167_a_248__dup_2141), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_2141), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6481 (.Q (
                         modgen_ram_ix167_a_247__dup_2142), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_2142), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6485 (.Q (
                         modgen_ram_ix167_a_246__dup_2143), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_2143), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6489 (.Q (
                         modgen_ram_ix167_a_245__dup_2144), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_2144), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6493 (.Q (
                         modgen_ram_ix167_a_244__dup_2145), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_2145), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6497 (.Q (
                         modgen_ram_ix167_a_243__dup_2146), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_2146), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6501 (.Q (
                         modgen_ram_ix167_a_242__dup_2147), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_2147), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6505 (.Q (
                         modgen_ram_ix167_a_241__dup_2148), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_2148), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6509 (.Q (
                         modgen_ram_ix167_a_240__dup_2149), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_2149), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6513 (.Q (
                         modgen_ram_ix167_a_239__dup_2150), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_2150), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6517 (.Q (
                         modgen_ram_ix167_a_238__dup_2151), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_2151), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6521 (.Q (
                         modgen_ram_ix167_a_237__dup_2152), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_2152), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6525 (.Q (
                         modgen_ram_ix167_a_236__dup_2153), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_2153), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6529 (.Q (
                         modgen_ram_ix167_a_235__dup_2154), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_2154), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6533 (.Q (
                         modgen_ram_ix167_a_234__dup_2155), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_2155), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6537 (.Q (
                         modgen_ram_ix167_a_233__dup_2156), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_2156), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6541 (.Q (
                         modgen_ram_ix167_a_232__dup_2157), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_2157), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6545 (.Q (
                         modgen_ram_ix167_a_231__dup_2158), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_2158), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6549 (.Q (
                         modgen_ram_ix167_a_230__dup_2159), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_2159), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6553 (.Q (
                         modgen_ram_ix167_a_229__dup_2160), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_2160), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6557 (.Q (
                         modgen_ram_ix167_a_228__dup_2161), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_2161), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6561 (.Q (
                         modgen_ram_ix167_a_227__dup_2162), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_2162), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6565 (.Q (
                         modgen_ram_ix167_a_226__dup_2163), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_2163), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6569 (.Q (
                         modgen_ram_ix167_a_225__dup_2164), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_2164), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6573 (.Q (
                         modgen_ram_ix167_a_224__dup_2165), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_2165), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6577 (.Q (
                         modgen_ram_ix167_a_223__dup_2166), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_2166), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6581 (.Q (
                         modgen_ram_ix167_a_222__dup_2167), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_2167), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6585 (.Q (
                         modgen_ram_ix167_a_221__dup_2168), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_2168), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6589 (.Q (
                         modgen_ram_ix167_a_220__dup_2169), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_2169), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6593 (.Q (
                         modgen_ram_ix167_a_219__dup_2170), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_2170), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6597 (.Q (
                         modgen_ram_ix167_a_218__dup_2171), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_2171), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6601 (.Q (
                         modgen_ram_ix167_a_217__dup_2172), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_2172), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6605 (.Q (
                         modgen_ram_ix167_a_216__dup_2173), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_2173), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6609 (.Q (
                         modgen_ram_ix167_a_215__dup_2174), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_2174), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6613 (.Q (
                         modgen_ram_ix167_a_214__dup_2175), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_2175), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6617 (.Q (
                         modgen_ram_ix167_a_213__dup_2176), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_2176), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6621 (.Q (
                         modgen_ram_ix167_a_212__dup_2177), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_2177), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6625 (.Q (
                         modgen_ram_ix167_a_211__dup_2178), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_2178), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6629 (.Q (
                         modgen_ram_ix167_a_210__dup_2179), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_2179), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6633 (.Q (
                         modgen_ram_ix167_a_209__dup_2180), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_2180), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6637 (.Q (
                         modgen_ram_ix167_a_208__dup_2181), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_2181), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6641 (.Q (
                         modgen_ram_ix167_a_207__dup_2182), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_2182), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6645 (.Q (
                         modgen_ram_ix167_a_206__dup_2183), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_2183), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6649 (.Q (
                         modgen_ram_ix167_a_205__dup_2184), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_2184), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6653 (.Q (
                         modgen_ram_ix167_a_204__dup_2185), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_2185), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6657 (.Q (
                         modgen_ram_ix167_a_203__dup_2186), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_2186), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6661 (.Q (
                         modgen_ram_ix167_a_202__dup_2187), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_2187), .SN (nx28501)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6665 (.Q (
                         modgen_ram_ix167_a_201__dup_2188), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_2188), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6669 (.Q (
                         modgen_ram_ix167_a_200__dup_2189), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_2189), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6673 (.Q (
                         modgen_ram_ix167_a_199__dup_2190), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_2190), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6677 (.Q (
                         modgen_ram_ix167_a_198__dup_2191), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_2191), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6681 (.Q (
                         modgen_ram_ix167_a_197__dup_2192), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_2192), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6685 (.Q (
                         modgen_ram_ix167_a_196__dup_2193), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_2193), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6689 (.Q (
                         modgen_ram_ix167_a_195__dup_2194), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_2194), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6693 (.Q (
                         modgen_ram_ix167_a_194__dup_2195), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_2195), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6697 (.Q (
                         modgen_ram_ix167_a_193__dup_2196), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_2196), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6701 (.Q (
                         modgen_ram_ix167_a_192__dup_2197), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_2197), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6705 (.Q (
                         modgen_ram_ix167_a_191__dup_2198), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_2198), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6709 (.Q (
                         modgen_ram_ix167_a_190__dup_2199), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_2199), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6713 (.Q (
                         modgen_ram_ix167_a_189__dup_2200), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_2200), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6717 (.Q (
                         modgen_ram_ix167_a_188__dup_2201), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_2201), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6721 (.Q (
                         modgen_ram_ix167_a_187__dup_2202), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_2202), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6725 (.Q (
                         modgen_ram_ix167_a_186__dup_2203), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_2203), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6729 (.Q (
                         modgen_ram_ix167_a_185__dup_2204), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_2204), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6733 (.Q (
                         modgen_ram_ix167_a_184__dup_2205), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_2205), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6737 (.Q (
                         modgen_ram_ix167_a_183__dup_2206), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_2206), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6741 (.Q (
                         modgen_ram_ix167_a_182__dup_2207), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_2207), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6745 (.Q (
                         modgen_ram_ix167_a_181__dup_2208), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_2208), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6749 (.Q (
                         modgen_ram_ix167_a_180__dup_2209), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_2209), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6753 (.Q (
                         modgen_ram_ix167_a_179__dup_2210), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_2210), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6757 (.Q (
                         modgen_ram_ix167_a_178__dup_2211), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_2211), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6761 (.Q (
                         modgen_ram_ix167_a_177__dup_2212), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_2212), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6765 (.Q (
                         modgen_ram_ix167_a_176__dup_2213), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_2213), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6769 (.Q (
                         modgen_ram_ix167_a_175__dup_2214), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_2214), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6773 (.Q (
                         modgen_ram_ix167_a_174__dup_2215), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_2215), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6777 (.Q (
                         modgen_ram_ix167_a_173__dup_2216), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_2216), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6781 (.Q (
                         modgen_ram_ix167_a_172__dup_2217), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_2217), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6785 (.Q (
                         modgen_ram_ix167_a_171__dup_2218), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_2218), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6789 (.Q (
                         modgen_ram_ix167_a_170__dup_2219), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_2219), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6793 (.Q (
                         modgen_ram_ix167_a_169__dup_2220), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_2220), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6797 (.Q (
                         modgen_ram_ix167_a_168__dup_2221), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_2221), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6801 (.Q (
                         modgen_ram_ix167_a_167__dup_2222), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_2222), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6805 (.Q (
                         modgen_ram_ix167_a_166__dup_2223), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_2223), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6809 (.Q (
                         modgen_ram_ix167_a_165__dup_2224), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_2224), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6813 (.Q (
                         modgen_ram_ix167_a_164__dup_2225), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_2225), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6817 (.Q (
                         modgen_ram_ix167_a_163__dup_2226), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_2226), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6821 (.Q (
                         modgen_ram_ix167_a_162__dup_2227), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_2227), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6825 (.Q (
                         modgen_ram_ix167_a_161__dup_2228), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_2228), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6829 (.Q (
                         modgen_ram_ix167_a_160__dup_2229), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_2229), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6833 (.Q (
                         modgen_ram_ix167_a_159__dup_2230), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_2230), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6837 (.Q (
                         modgen_ram_ix167_a_158__dup_2231), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_2231), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6841 (.Q (
                         modgen_ram_ix167_a_157__dup_2232), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_2232), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6845 (.Q (
                         modgen_ram_ix167_a_156__dup_2233), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_2233), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6849 (.Q (
                         modgen_ram_ix167_a_155__dup_2234), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_2234), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6853 (.Q (
                         modgen_ram_ix167_a_154__dup_2235), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_2235), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6857 (.Q (
                         modgen_ram_ix167_a_153__dup_2236), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_2236), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6861 (.Q (
                         modgen_ram_ix167_a_152__dup_2237), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_2237), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6865 (.Q (
                         modgen_ram_ix167_a_151__dup_2238), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_2238), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6869 (.Q (
                         modgen_ram_ix167_a_150__dup_2239), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_2239), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6873 (.Q (
                         modgen_ram_ix167_a_149__dup_2240), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_2240), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6877 (.Q (
                         modgen_ram_ix167_a_148__dup_2241), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_2241), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6881 (.Q (
                         modgen_ram_ix167_a_147__dup_2242), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_2242), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6885 (.Q (
                         modgen_ram_ix167_a_146__dup_2243), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_2243), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6889 (.Q (
                         modgen_ram_ix167_a_145__dup_2244), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_2244), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6893 (.Q (
                         modgen_ram_ix167_a_144__dup_2245), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_2245), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6897 (.Q (
                         modgen_ram_ix167_a_143__dup_2246), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_2246), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6901 (.Q (
                         modgen_ram_ix167_a_142__dup_2247), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_2247), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6905 (.Q (
                         modgen_ram_ix167_a_141__dup_2248), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_2248), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6909 (.Q (
                         modgen_ram_ix167_a_140__dup_2249), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_2249), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6913 (.Q (
                         modgen_ram_ix167_a_139__dup_2250), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_2250), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6917 (.Q (
                         modgen_ram_ix167_a_138__dup_2251), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_2251), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6921 (.Q (
                         modgen_ram_ix167_a_137__dup_2252), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_2252), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6925 (.Q (
                         modgen_ram_ix167_a_136__dup_2253), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_2253), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6929 (.Q (
                         modgen_ram_ix167_a_135__dup_2254), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_2254), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6933 (.Q (
                         modgen_ram_ix167_a_134__dup_2255), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_2255), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6937 (.Q (
                         modgen_ram_ix167_a_133__dup_2256), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_2256), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6941 (.Q (
                         modgen_ram_ix167_a_132__dup_2257), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_2257), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6945 (.Q (
                         modgen_ram_ix167_a_131__dup_2258), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_2258), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6949 (.Q (
                         modgen_ram_ix167_a_130__dup_2259), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_2259), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6953 (.Q (
                         modgen_ram_ix167_a_129__dup_2260), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_2260), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6957 (.Q (
                         modgen_ram_ix167_a_128__dup_2261), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_2261), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6961 (.Q (
                         modgen_ram_ix167_a_127__dup_2262), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_2262), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6965 (.Q (
                         modgen_ram_ix167_a_126__dup_2263), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_2263), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6969 (.Q (
                         modgen_ram_ix167_a_125__dup_2264), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_2264), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6973 (.Q (
                         modgen_ram_ix167_a_124__dup_2265), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_2265), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6977 (.Q (
                         modgen_ram_ix167_a_123__dup_2266), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_2266), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6981 (.Q (
                         modgen_ram_ix167_a_122__dup_2267), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_2267), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6985 (.Q (
                         modgen_ram_ix167_a_121__dup_2268), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_2268), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6989 (.Q (
                         modgen_ram_ix167_a_120__dup_2269), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_2269), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6993 (.Q (
                         modgen_ram_ix167_a_119__dup_2270), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_2270), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix6997 (.Q (
                         modgen_ram_ix167_a_118__dup_2271), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_2271), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7001 (.Q (
                         modgen_ram_ix167_a_117__dup_2272), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_2272), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7005 (.Q (
                         modgen_ram_ix167_a_116__dup_2273), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_2273), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7009 (.Q (
                         modgen_ram_ix167_a_115__dup_2274), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_2274), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7013 (.Q (
                         modgen_ram_ix167_a_114__dup_2275), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_2275), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7017 (.Q (
                         modgen_ram_ix167_a_113__dup_2276), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_2276), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7021 (.Q (
                         modgen_ram_ix167_a_112__dup_2277), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_2277), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7025 (.Q (
                         modgen_ram_ix167_a_111__dup_2278), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_2278), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7029 (.Q (
                         modgen_ram_ix167_a_110__dup_2279), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_2279), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7033 (.Q (
                         modgen_ram_ix167_a_109__dup_2280), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_2280), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7037 (.Q (
                         modgen_ram_ix167_a_108__dup_2281), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_2281), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7041 (.Q (
                         modgen_ram_ix167_a_107__dup_2282), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_2282), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7045 (.Q (
                         modgen_ram_ix167_a_106__dup_2283), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_2283), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7049 (.Q (
                         modgen_ram_ix167_a_105__dup_2284), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_2284), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7053 (.Q (
                         modgen_ram_ix167_a_104__dup_2285), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_2285), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7057 (.Q (
                         modgen_ram_ix167_a_103__dup_2286), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_2286), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7061 (.Q (
                         modgen_ram_ix167_a_102__dup_2287), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_2287), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7065 (.Q (
                         modgen_ram_ix167_a_101__dup_2288), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_2288), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7069 (.Q (
                         modgen_ram_ix167_a_100__dup_2289), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_2289), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7073 (.Q (
                         modgen_ram_ix167_a_99__dup_2290), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_2290), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7077 (.Q (
                         modgen_ram_ix167_a_98__dup_2291), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_2291), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7081 (.Q (
                         modgen_ram_ix167_a_97__dup_2292), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_2292), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7085 (.Q (
                         modgen_ram_ix167_a_96__dup_2293), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_2293), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7089 (.Q (
                         modgen_ram_ix167_a_95__dup_2294), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_2294), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7093 (.Q (
                         modgen_ram_ix167_a_94__dup_2295), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_2295), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7097 (.Q (
                         modgen_ram_ix167_a_93__dup_2296), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_2296), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7101 (.Q (
                         modgen_ram_ix167_a_92__dup_2297), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_2297), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7105 (.Q (
                         modgen_ram_ix167_a_91__dup_2298), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_2298), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7109 (.Q (
                         modgen_ram_ix167_a_90__dup_2299), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_2299), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7113 (.Q (
                         modgen_ram_ix167_a_89__dup_2300), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_2300), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7117 (.Q (
                         modgen_ram_ix167_a_88__dup_2301), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_2301), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7121 (.Q (
                         modgen_ram_ix167_a_87__dup_2302), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_2302), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7125 (.Q (
                         modgen_ram_ix167_a_86__dup_2303), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_2303), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7129 (.Q (
                         modgen_ram_ix167_a_85__dup_2304), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_2304), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7133 (.Q (
                         modgen_ram_ix167_a_84__dup_2305), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_2305), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7137 (.Q (
                         modgen_ram_ix167_a_83__dup_2306), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_2306), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7141 (.Q (
                         modgen_ram_ix167_a_82__dup_2307), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_2307), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7145 (.Q (
                         modgen_ram_ix167_a_81__dup_2308), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_2308), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7149 (.Q (
                         modgen_ram_ix167_a_80__dup_2309), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_2309), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7153 (.Q (
                         modgen_ram_ix167_a_79__dup_2310), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_2310), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7157 (.Q (
                         modgen_ram_ix167_a_78__dup_2311), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_2311), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7161 (.Q (
                         modgen_ram_ix167_a_77__dup_2312), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_2312), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7165 (.Q (
                         modgen_ram_ix167_a_76__dup_2313), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_2313), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7169 (.Q (
                         modgen_ram_ix167_a_75__dup_2314), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_2314), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7173 (.Q (
                         modgen_ram_ix167_a_74__dup_2315), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_2315), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7177 (.Q (
                         modgen_ram_ix167_a_73__dup_2316), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_2316), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7181 (.Q (
                         modgen_ram_ix167_a_72__dup_2317), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_2317), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7185 (.Q (
                         modgen_ram_ix167_a_71__dup_2318), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_2318), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7189 (.Q (
                         modgen_ram_ix167_a_70__dup_2319), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_2319), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7193 (.Q (
                         modgen_ram_ix167_a_69__dup_2320), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_2320), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7197 (.Q (
                         modgen_ram_ix167_a_68__dup_2321), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_2321), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7201 (.Q (
                         modgen_ram_ix167_a_67__dup_2322), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_2322), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7205 (.Q (
                         modgen_ram_ix167_a_66__dup_2323), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_2323), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7209 (.Q (
                         modgen_ram_ix167_a_65__dup_2324), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_2324), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7213 (.Q (
                         modgen_ram_ix167_a_64__dup_2325), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_2325), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7217 (.Q (
                         modgen_ram_ix167_a_63__dup_2326), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_2326), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7221 (.Q (
                         modgen_ram_ix167_a_62__dup_2327), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_2327), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7225 (.Q (
                         modgen_ram_ix167_a_61__dup_2328), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_2328), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7229 (.Q (
                         modgen_ram_ix167_a_60__dup_2329), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_2329), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7233 (.Q (
                         modgen_ram_ix167_a_59__dup_2330), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_2330), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7237 (.Q (
                         modgen_ram_ix167_a_58__dup_2331), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_2331), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7241 (.Q (
                         modgen_ram_ix167_a_57__dup_2332), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_2332), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7245 (.Q (
                         modgen_ram_ix167_a_56__dup_2333), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_2333), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7249 (.Q (
                         modgen_ram_ix167_a_55__dup_2334), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_2334), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7253 (.Q (
                         modgen_ram_ix167_a_54__dup_2335), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_2335), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7257 (.Q (
                         modgen_ram_ix167_a_53__dup_2336), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_2336), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7261 (.Q (
                         modgen_ram_ix167_a_52__dup_2337), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_2337), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7265 (.Q (
                         modgen_ram_ix167_a_51__dup_2338), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_2338), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7269 (.Q (
                         modgen_ram_ix167_a_50__dup_2339), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_2339), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7273 (.Q (
                         modgen_ram_ix167_a_49__dup_2340), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_2340), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7277 (.Q (
                         modgen_ram_ix167_a_48__dup_2341), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_2341), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7281 (.Q (
                         modgen_ram_ix167_a_47__dup_2342), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_2342), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7285 (.Q (
                         modgen_ram_ix167_a_46__dup_2343), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_2343), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7289 (.Q (
                         modgen_ram_ix167_a_45__dup_2344), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_2344), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7293 (.Q (
                         modgen_ram_ix167_a_44__dup_2345), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_2345), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7297 (.Q (
                         modgen_ram_ix167_a_43__dup_2346), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_2346), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7301 (.Q (
                         modgen_ram_ix167_a_42__dup_2347), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_2347), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7305 (.Q (
                         modgen_ram_ix167_a_41__dup_2348), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_2348), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7309 (.Q (
                         modgen_ram_ix167_a_40__dup_2349), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_2349), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7313 (.Q (
                         modgen_ram_ix167_a_39__dup_2350), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_2350), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7317 (.Q (
                         modgen_ram_ix167_a_38__dup_2351), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_2351), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7321 (.Q (
                         modgen_ram_ix167_a_37__dup_2352), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_2352), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7325 (.Q (
                         modgen_ram_ix167_a_36__dup_2353), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_2353), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7329 (.Q (
                         modgen_ram_ix167_a_35__dup_2354), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_2354), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7333 (.Q (
                         modgen_ram_ix167_a_34__dup_2355), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_2355), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7337 (.Q (
                         modgen_ram_ix167_a_33__dup_2356), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_2356), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7341 (.Q (
                         modgen_ram_ix167_a_32__dup_2357), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_2357), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7345 (.Q (
                         modgen_ram_ix167_a_31__dup_2358), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_2358), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7349 (.Q (
                         modgen_ram_ix167_a_30__dup_2359), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_2359), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7353 (.Q (
                         modgen_ram_ix167_a_29__dup_2360), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_2360), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7357 (.Q (
                         modgen_ram_ix167_a_28__dup_2361), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_2361), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7361 (.Q (
                         modgen_ram_ix167_a_27__dup_2362), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_2362), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7365 (.Q (
                         modgen_ram_ix167_a_26__dup_2363), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_2363), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7369 (.Q (
                         modgen_ram_ix167_a_25__dup_2364), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_2364), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7373 (.Q (
                         modgen_ram_ix167_a_24__dup_2365), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_2365), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7377 (.Q (
                         modgen_ram_ix167_a_23__dup_2366), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_2366), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7381 (.Q (
                         modgen_ram_ix167_a_22__dup_2367), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_2367), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7385 (.Q (
                         modgen_ram_ix167_a_21__dup_2368), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_2368), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7389 (.Q (
                         modgen_ram_ix167_a_20__dup_2369), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_2369), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7393 (.Q (
                         modgen_ram_ix167_a_19__dup_2370), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_2370), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7397 (.Q (
                         modgen_ram_ix167_a_18__dup_2371), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_2371), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7401 (.Q (
                         modgen_ram_ix167_a_17__dup_2372), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_2372), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7405 (.Q (
                         modgen_ram_ix167_a_16__dup_2373), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_2373), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7409 (.Q (
                         modgen_ram_ix167_a_15__dup_2374), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_2374), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7413 (.Q (
                         modgen_ram_ix167_a_14__dup_2375), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_2375), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7417 (.Q (
                         modgen_ram_ix167_a_13__dup_2376), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_2376), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7421 (.Q (
                         modgen_ram_ix167_a_12__dup_2377), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_2377), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7425 (.Q (
                         modgen_ram_ix167_a_11__dup_2378), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_2378), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7429 (.Q (
                         modgen_ram_ix167_a_10__dup_2379), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_2379), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7433 (.Q (
                         modgen_ram_ix167_a_9__dup_2380), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_2380), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7437 (.Q (
                         modgen_ram_ix167_a_8__dup_2381), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_2381), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7441 (.Q (
                         modgen_ram_ix167_a_7__dup_2382), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_2382), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7445 (.Q (
                         modgen_ram_ix167_a_6__dup_2383), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_2383), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7449 (.Q (
                         modgen_ram_ix167_a_5__dup_2384), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_2384), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7453 (.Q (
                         modgen_ram_ix167_a_4__dup_2385), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_2385), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7457 (.Q (
                         modgen_ram_ix167_a_3__dup_2386), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_2386), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7461 (.Q (
                         modgen_ram_ix167_a_2__dup_2387), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_2387), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7465 (.Q (
                         modgen_ram_ix167_a_1__dup_2388), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_2388), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7469 (.Q (
                         modgen_ram_ix167_a_0__dup_2389), .CK (wb_clk_i), .D (
                         nx28521), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_2389), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7474 (.Q (
                         modgen_ram_ix167_a_255__dup_2398), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5764), .SI (
                         modgen_ram_ix167_a_255__dup_2398), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7478 (.Q (
                         modgen_ram_ix167_a_254__dup_2399), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5746), .SI (
                         modgen_ram_ix167_a_254__dup_2399), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7482 (.Q (
                         modgen_ram_ix167_a_253__dup_2400), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5724), .SI (
                         modgen_ram_ix167_a_253__dup_2400), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7486 (.Q (
                         modgen_ram_ix167_a_252__dup_2401), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5706), .SI (
                         modgen_ram_ix167_a_252__dup_2401), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7490 (.Q (
                         modgen_ram_ix167_a_251__dup_2402), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5680), .SI (
                         modgen_ram_ix167_a_251__dup_2402), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7494 (.Q (
                         modgen_ram_ix167_a_250__dup_2403), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5662), .SI (
                         modgen_ram_ix167_a_250__dup_2403), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7498 (.Q (
                         modgen_ram_ix167_a_249__dup_2404), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5640), .SI (
                         modgen_ram_ix167_a_249__dup_2404), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7502 (.Q (
                         modgen_ram_ix167_a_248__dup_2405), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5622), .SI (
                         modgen_ram_ix167_a_248__dup_2405), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7506 (.Q (
                         modgen_ram_ix167_a_247__dup_2406), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5592), .SI (
                         modgen_ram_ix167_a_247__dup_2406), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7510 (.Q (
                         modgen_ram_ix167_a_246__dup_2407), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5574), .SI (
                         modgen_ram_ix167_a_246__dup_2407), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7514 (.Q (
                         modgen_ram_ix167_a_245__dup_2408), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5552), .SI (
                         modgen_ram_ix167_a_245__dup_2408), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7518 (.Q (
                         modgen_ram_ix167_a_244__dup_2409), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5534), .SI (
                         modgen_ram_ix167_a_244__dup_2409), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7522 (.Q (
                         modgen_ram_ix167_a_243__dup_2410), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5508), .SI (
                         modgen_ram_ix167_a_243__dup_2410), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7526 (.Q (
                         modgen_ram_ix167_a_242__dup_2411), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5490), .SI (
                         modgen_ram_ix167_a_242__dup_2411), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7530 (.Q (
                         modgen_ram_ix167_a_241__dup_2412), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5468), .SI (
                         modgen_ram_ix167_a_241__dup_2412), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7534 (.Q (
                         modgen_ram_ix167_a_240__dup_2413), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5450), .SI (
                         modgen_ram_ix167_a_240__dup_2413), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7538 (.Q (
                         modgen_ram_ix167_a_239__dup_2414), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5414), .SI (
                         modgen_ram_ix167_a_239__dup_2414), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7542 (.Q (
                         modgen_ram_ix167_a_238__dup_2415), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5396), .SI (
                         modgen_ram_ix167_a_238__dup_2415), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7546 (.Q (
                         modgen_ram_ix167_a_237__dup_2416), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5374), .SI (
                         modgen_ram_ix167_a_237__dup_2416), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7550 (.Q (
                         modgen_ram_ix167_a_236__dup_2417), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5356), .SI (
                         modgen_ram_ix167_a_236__dup_2417), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7554 (.Q (
                         modgen_ram_ix167_a_235__dup_2418), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5330), .SI (
                         modgen_ram_ix167_a_235__dup_2418), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7558 (.Q (
                         modgen_ram_ix167_a_234__dup_2419), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5312), .SI (
                         modgen_ram_ix167_a_234__dup_2419), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7562 (.Q (
                         modgen_ram_ix167_a_233__dup_2420), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5290), .SI (
                         modgen_ram_ix167_a_233__dup_2420), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7566 (.Q (
                         modgen_ram_ix167_a_232__dup_2421), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5272), .SI (
                         modgen_ram_ix167_a_232__dup_2421), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7570 (.Q (
                         modgen_ram_ix167_a_231__dup_2422), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5242), .SI (
                         modgen_ram_ix167_a_231__dup_2422), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7574 (.Q (
                         modgen_ram_ix167_a_230__dup_2423), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5224), .SI (
                         modgen_ram_ix167_a_230__dup_2423), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7578 (.Q (
                         modgen_ram_ix167_a_229__dup_2424), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5202), .SI (
                         modgen_ram_ix167_a_229__dup_2424), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7582 (.Q (
                         modgen_ram_ix167_a_228__dup_2425), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5184), .SI (
                         modgen_ram_ix167_a_228__dup_2425), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7586 (.Q (
                         modgen_ram_ix167_a_227__dup_2426), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5158), .SI (
                         modgen_ram_ix167_a_227__dup_2426), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7590 (.Q (
                         modgen_ram_ix167_a_226__dup_2427), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5140), .SI (
                         modgen_ram_ix167_a_226__dup_2427), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7594 (.Q (
                         modgen_ram_ix167_a_225__dup_2428), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5118), .SI (
                         modgen_ram_ix167_a_225__dup_2428), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7598 (.Q (
                         modgen_ram_ix167_a_224__dup_2429), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5100), .SI (
                         modgen_ram_ix167_a_224__dup_2429), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7602 (.Q (
                         modgen_ram_ix167_a_223__dup_2430), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5060), .SI (
                         modgen_ram_ix167_a_223__dup_2430), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7606 (.Q (
                         modgen_ram_ix167_a_222__dup_2431), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5042), .SI (
                         modgen_ram_ix167_a_222__dup_2431), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7610 (.Q (
                         modgen_ram_ix167_a_221__dup_2432), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5020), .SI (
                         modgen_ram_ix167_a_221__dup_2432), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7614 (.Q (
                         modgen_ram_ix167_a_220__dup_2433), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx5002), .SI (
                         modgen_ram_ix167_a_220__dup_2433), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7618 (.Q (
                         modgen_ram_ix167_a_219__dup_2434), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4976), .SI (
                         modgen_ram_ix167_a_219__dup_2434), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7622 (.Q (
                         modgen_ram_ix167_a_218__dup_2435), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4958), .SI (
                         modgen_ram_ix167_a_218__dup_2435), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7626 (.Q (
                         modgen_ram_ix167_a_217__dup_2436), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4936), .SI (
                         modgen_ram_ix167_a_217__dup_2436), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7630 (.Q (
                         modgen_ram_ix167_a_216__dup_2437), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4918), .SI (
                         modgen_ram_ix167_a_216__dup_2437), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7634 (.Q (
                         modgen_ram_ix167_a_215__dup_2438), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4888), .SI (
                         modgen_ram_ix167_a_215__dup_2438), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7638 (.Q (
                         modgen_ram_ix167_a_214__dup_2439), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4870), .SI (
                         modgen_ram_ix167_a_214__dup_2439), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7642 (.Q (
                         modgen_ram_ix167_a_213__dup_2440), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4848), .SI (
                         modgen_ram_ix167_a_213__dup_2440), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7646 (.Q (
                         modgen_ram_ix167_a_212__dup_2441), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4830), .SI (
                         modgen_ram_ix167_a_212__dup_2441), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7650 (.Q (
                         modgen_ram_ix167_a_211__dup_2442), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4804), .SI (
                         modgen_ram_ix167_a_211__dup_2442), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7654 (.Q (
                         modgen_ram_ix167_a_210__dup_2443), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4786), .SI (
                         modgen_ram_ix167_a_210__dup_2443), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7658 (.Q (
                         modgen_ram_ix167_a_209__dup_2444), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4764), .SI (
                         modgen_ram_ix167_a_209__dup_2444), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7662 (.Q (
                         modgen_ram_ix167_a_208__dup_2445), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4746), .SI (
                         modgen_ram_ix167_a_208__dup_2445), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7666 (.Q (
                         modgen_ram_ix167_a_207__dup_2446), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4710), .SI (
                         modgen_ram_ix167_a_207__dup_2446), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7670 (.Q (
                         modgen_ram_ix167_a_206__dup_2447), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4692), .SI (
                         modgen_ram_ix167_a_206__dup_2447), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7674 (.Q (
                         modgen_ram_ix167_a_205__dup_2448), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4670), .SI (
                         modgen_ram_ix167_a_205__dup_2448), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7678 (.Q (
                         modgen_ram_ix167_a_204__dup_2449), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4652), .SI (
                         modgen_ram_ix167_a_204__dup_2449), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7682 (.Q (
                         modgen_ram_ix167_a_203__dup_2450), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4626), .SI (
                         modgen_ram_ix167_a_203__dup_2450), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7686 (.Q (
                         modgen_ram_ix167_a_202__dup_2451), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4608), .SI (
                         modgen_ram_ix167_a_202__dup_2451), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7690 (.Q (
                         modgen_ram_ix167_a_201__dup_2452), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4586), .SI (
                         modgen_ram_ix167_a_201__dup_2452), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7694 (.Q (
                         modgen_ram_ix167_a_200__dup_2453), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4568), .SI (
                         modgen_ram_ix167_a_200__dup_2453), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7698 (.Q (
                         modgen_ram_ix167_a_199__dup_2454), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4538), .SI (
                         modgen_ram_ix167_a_199__dup_2454), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7702 (.Q (
                         modgen_ram_ix167_a_198__dup_2455), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4520), .SI (
                         modgen_ram_ix167_a_198__dup_2455), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7706 (.Q (
                         modgen_ram_ix167_a_197__dup_2456), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4498), .SI (
                         modgen_ram_ix167_a_197__dup_2456), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7710 (.Q (
                         modgen_ram_ix167_a_196__dup_2457), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4480), .SI (
                         modgen_ram_ix167_a_196__dup_2457), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7714 (.Q (
                         modgen_ram_ix167_a_195__dup_2458), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4454), .SI (
                         modgen_ram_ix167_a_195__dup_2458), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7718 (.Q (
                         modgen_ram_ix167_a_194__dup_2459), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4436), .SI (
                         modgen_ram_ix167_a_194__dup_2459), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7722 (.Q (
                         modgen_ram_ix167_a_193__dup_2460), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4414), .SI (
                         modgen_ram_ix167_a_193__dup_2460), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7726 (.Q (
                         modgen_ram_ix167_a_192__dup_2461), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4396), .SI (
                         modgen_ram_ix167_a_192__dup_2461), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7730 (.Q (
                         modgen_ram_ix167_a_191__dup_2462), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4346), .SI (
                         modgen_ram_ix167_a_191__dup_2462), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7734 (.Q (
                         modgen_ram_ix167_a_190__dup_2463), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4328), .SI (
                         modgen_ram_ix167_a_190__dup_2463), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7738 (.Q (
                         modgen_ram_ix167_a_189__dup_2464), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4306), .SI (
                         modgen_ram_ix167_a_189__dup_2464), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7742 (.Q (
                         modgen_ram_ix167_a_188__dup_2465), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4288), .SI (
                         modgen_ram_ix167_a_188__dup_2465), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7746 (.Q (
                         modgen_ram_ix167_a_187__dup_2466), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4262), .SI (
                         modgen_ram_ix167_a_187__dup_2466), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7750 (.Q (
                         modgen_ram_ix167_a_186__dup_2467), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4244), .SI (
                         modgen_ram_ix167_a_186__dup_2467), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7754 (.Q (
                         modgen_ram_ix167_a_185__dup_2468), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4222), .SI (
                         modgen_ram_ix167_a_185__dup_2468), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7758 (.Q (
                         modgen_ram_ix167_a_184__dup_2469), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4204), .SI (
                         modgen_ram_ix167_a_184__dup_2469), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7762 (.Q (
                         modgen_ram_ix167_a_183__dup_2470), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4174), .SI (
                         modgen_ram_ix167_a_183__dup_2470), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7766 (.Q (
                         modgen_ram_ix167_a_182__dup_2471), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4156), .SI (
                         modgen_ram_ix167_a_182__dup_2471), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7770 (.Q (
                         modgen_ram_ix167_a_181__dup_2472), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4134), .SI (
                         modgen_ram_ix167_a_181__dup_2472), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7774 (.Q (
                         modgen_ram_ix167_a_180__dup_2473), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4116), .SI (
                         modgen_ram_ix167_a_180__dup_2473), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7778 (.Q (
                         modgen_ram_ix167_a_179__dup_2474), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4090), .SI (
                         modgen_ram_ix167_a_179__dup_2474), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7782 (.Q (
                         modgen_ram_ix167_a_178__dup_2475), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4072), .SI (
                         modgen_ram_ix167_a_178__dup_2475), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7786 (.Q (
                         modgen_ram_ix167_a_177__dup_2476), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4050), .SI (
                         modgen_ram_ix167_a_177__dup_2476), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7790 (.Q (
                         modgen_ram_ix167_a_176__dup_2477), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx4032), .SI (
                         modgen_ram_ix167_a_176__dup_2477), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7794 (.Q (
                         modgen_ram_ix167_a_175__dup_2478), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3996), .SI (
                         modgen_ram_ix167_a_175__dup_2478), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7798 (.Q (
                         modgen_ram_ix167_a_174__dup_2479), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3978), .SI (
                         modgen_ram_ix167_a_174__dup_2479), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7802 (.Q (
                         modgen_ram_ix167_a_173__dup_2480), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3956), .SI (
                         modgen_ram_ix167_a_173__dup_2480), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7806 (.Q (
                         modgen_ram_ix167_a_172__dup_2481), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3938), .SI (
                         modgen_ram_ix167_a_172__dup_2481), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7810 (.Q (
                         modgen_ram_ix167_a_171__dup_2482), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3912), .SI (
                         modgen_ram_ix167_a_171__dup_2482), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7814 (.Q (
                         modgen_ram_ix167_a_170__dup_2483), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3894), .SI (
                         modgen_ram_ix167_a_170__dup_2483), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7818 (.Q (
                         modgen_ram_ix167_a_169__dup_2484), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3872), .SI (
                         modgen_ram_ix167_a_169__dup_2484), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7822 (.Q (
                         modgen_ram_ix167_a_168__dup_2485), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3854), .SI (
                         modgen_ram_ix167_a_168__dup_2485), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7826 (.Q (
                         modgen_ram_ix167_a_167__dup_2486), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3824), .SI (
                         modgen_ram_ix167_a_167__dup_2486), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7830 (.Q (
                         modgen_ram_ix167_a_166__dup_2487), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3806), .SI (
                         modgen_ram_ix167_a_166__dup_2487), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7834 (.Q (
                         modgen_ram_ix167_a_165__dup_2488), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3784), .SI (
                         modgen_ram_ix167_a_165__dup_2488), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7838 (.Q (
                         modgen_ram_ix167_a_164__dup_2489), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3766), .SI (
                         modgen_ram_ix167_a_164__dup_2489), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7842 (.Q (
                         modgen_ram_ix167_a_163__dup_2490), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3740), .SI (
                         modgen_ram_ix167_a_163__dup_2490), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7846 (.Q (
                         modgen_ram_ix167_a_162__dup_2491), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3722), .SI (
                         modgen_ram_ix167_a_162__dup_2491), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7850 (.Q (
                         modgen_ram_ix167_a_161__dup_2492), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3700), .SI (
                         modgen_ram_ix167_a_161__dup_2492), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7854 (.Q (
                         modgen_ram_ix167_a_160__dup_2493), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3682), .SI (
                         modgen_ram_ix167_a_160__dup_2493), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7858 (.Q (
                         modgen_ram_ix167_a_159__dup_2494), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3642), .SI (
                         modgen_ram_ix167_a_159__dup_2494), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7862 (.Q (
                         modgen_ram_ix167_a_158__dup_2495), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3624), .SI (
                         modgen_ram_ix167_a_158__dup_2495), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7866 (.Q (
                         modgen_ram_ix167_a_157__dup_2496), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3602), .SI (
                         modgen_ram_ix167_a_157__dup_2496), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7870 (.Q (
                         modgen_ram_ix167_a_156__dup_2497), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3584), .SI (
                         modgen_ram_ix167_a_156__dup_2497), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7874 (.Q (
                         modgen_ram_ix167_a_155__dup_2498), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3558), .SI (
                         modgen_ram_ix167_a_155__dup_2498), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7878 (.Q (
                         modgen_ram_ix167_a_154__dup_2499), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3540), .SI (
                         modgen_ram_ix167_a_154__dup_2499), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7882 (.Q (
                         modgen_ram_ix167_a_153__dup_2500), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3518), .SI (
                         modgen_ram_ix167_a_153__dup_2500), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7886 (.Q (
                         modgen_ram_ix167_a_152__dup_2501), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3500), .SI (
                         modgen_ram_ix167_a_152__dup_2501), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7890 (.Q (
                         modgen_ram_ix167_a_151__dup_2502), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3470), .SI (
                         modgen_ram_ix167_a_151__dup_2502), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7894 (.Q (
                         modgen_ram_ix167_a_150__dup_2503), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3452), .SI (
                         modgen_ram_ix167_a_150__dup_2503), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7898 (.Q (
                         modgen_ram_ix167_a_149__dup_2504), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3430), .SI (
                         modgen_ram_ix167_a_149__dup_2504), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7902 (.Q (
                         modgen_ram_ix167_a_148__dup_2505), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3412), .SI (
                         modgen_ram_ix167_a_148__dup_2505), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7906 (.Q (
                         modgen_ram_ix167_a_147__dup_2506), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3386), .SI (
                         modgen_ram_ix167_a_147__dup_2506), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7910 (.Q (
                         modgen_ram_ix167_a_146__dup_2507), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3368), .SI (
                         modgen_ram_ix167_a_146__dup_2507), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7914 (.Q (
                         modgen_ram_ix167_a_145__dup_2508), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3346), .SI (
                         modgen_ram_ix167_a_145__dup_2508), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7918 (.Q (
                         modgen_ram_ix167_a_144__dup_2509), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3328), .SI (
                         modgen_ram_ix167_a_144__dup_2509), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7922 (.Q (
                         modgen_ram_ix167_a_143__dup_2510), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3292), .SI (
                         modgen_ram_ix167_a_143__dup_2510), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7926 (.Q (
                         modgen_ram_ix167_a_142__dup_2511), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3274), .SI (
                         modgen_ram_ix167_a_142__dup_2511), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7930 (.Q (
                         modgen_ram_ix167_a_141__dup_2512), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3252), .SI (
                         modgen_ram_ix167_a_141__dup_2512), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7934 (.Q (
                         modgen_ram_ix167_a_140__dup_2513), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3234), .SI (
                         modgen_ram_ix167_a_140__dup_2513), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7938 (.Q (
                         modgen_ram_ix167_a_139__dup_2514), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3208), .SI (
                         modgen_ram_ix167_a_139__dup_2514), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7942 (.Q (
                         modgen_ram_ix167_a_138__dup_2515), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3190), .SI (
                         modgen_ram_ix167_a_138__dup_2515), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7946 (.Q (
                         modgen_ram_ix167_a_137__dup_2516), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3168), .SI (
                         modgen_ram_ix167_a_137__dup_2516), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7950 (.Q (
                         modgen_ram_ix167_a_136__dup_2517), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3150), .SI (
                         modgen_ram_ix167_a_136__dup_2517), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7954 (.Q (
                         modgen_ram_ix167_a_135__dup_2518), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3120), .SI (
                         modgen_ram_ix167_a_135__dup_2518), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7958 (.Q (
                         modgen_ram_ix167_a_134__dup_2519), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3102), .SI (
                         modgen_ram_ix167_a_134__dup_2519), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7962 (.Q (
                         modgen_ram_ix167_a_133__dup_2520), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3080), .SI (
                         modgen_ram_ix167_a_133__dup_2520), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7966 (.Q (
                         modgen_ram_ix167_a_132__dup_2521), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3062), .SI (
                         modgen_ram_ix167_a_132__dup_2521), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7970 (.Q (
                         modgen_ram_ix167_a_131__dup_2522), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3036), .SI (
                         modgen_ram_ix167_a_131__dup_2522), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7974 (.Q (
                         modgen_ram_ix167_a_130__dup_2523), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx3018), .SI (
                         modgen_ram_ix167_a_130__dup_2523), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7978 (.Q (
                         modgen_ram_ix167_a_129__dup_2524), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2996), .SI (
                         modgen_ram_ix167_a_129__dup_2524), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7982 (.Q (
                         modgen_ram_ix167_a_128__dup_2525), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2978), .SI (
                         modgen_ram_ix167_a_128__dup_2525), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7986 (.Q (
                         modgen_ram_ix167_a_127__dup_2526), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2926), .SI (
                         modgen_ram_ix167_a_127__dup_2526), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7990 (.Q (
                         modgen_ram_ix167_a_126__dup_2527), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2908), .SI (
                         modgen_ram_ix167_a_126__dup_2527), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7994 (.Q (
                         modgen_ram_ix167_a_125__dup_2528), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2886), .SI (
                         modgen_ram_ix167_a_125__dup_2528), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix7998 (.Q (
                         modgen_ram_ix167_a_124__dup_2529), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2868), .SI (
                         modgen_ram_ix167_a_124__dup_2529), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8002 (.Q (
                         modgen_ram_ix167_a_123__dup_2530), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2842), .SI (
                         modgen_ram_ix167_a_123__dup_2530), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8006 (.Q (
                         modgen_ram_ix167_a_122__dup_2531), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2824), .SI (
                         modgen_ram_ix167_a_122__dup_2531), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8010 (.Q (
                         modgen_ram_ix167_a_121__dup_2532), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2802), .SI (
                         modgen_ram_ix167_a_121__dup_2532), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8014 (.Q (
                         modgen_ram_ix167_a_120__dup_2533), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2784), .SI (
                         modgen_ram_ix167_a_120__dup_2533), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8018 (.Q (
                         modgen_ram_ix167_a_119__dup_2534), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2754), .SI (
                         modgen_ram_ix167_a_119__dup_2534), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8022 (.Q (
                         modgen_ram_ix167_a_118__dup_2535), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2736), .SI (
                         modgen_ram_ix167_a_118__dup_2535), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8026 (.Q (
                         modgen_ram_ix167_a_117__dup_2536), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2714), .SI (
                         modgen_ram_ix167_a_117__dup_2536), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8030 (.Q (
                         modgen_ram_ix167_a_116__dup_2537), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2696), .SI (
                         modgen_ram_ix167_a_116__dup_2537), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8034 (.Q (
                         modgen_ram_ix167_a_115__dup_2538), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2670), .SI (
                         modgen_ram_ix167_a_115__dup_2538), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8038 (.Q (
                         modgen_ram_ix167_a_114__dup_2539), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2652), .SI (
                         modgen_ram_ix167_a_114__dup_2539), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8042 (.Q (
                         modgen_ram_ix167_a_113__dup_2540), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2630), .SI (
                         modgen_ram_ix167_a_113__dup_2540), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8046 (.Q (
                         modgen_ram_ix167_a_112__dup_2541), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2612), .SI (
                         modgen_ram_ix167_a_112__dup_2541), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8050 (.Q (
                         modgen_ram_ix167_a_111__dup_2542), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2576), .SI (
                         modgen_ram_ix167_a_111__dup_2542), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8054 (.Q (
                         modgen_ram_ix167_a_110__dup_2543), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2558), .SI (
                         modgen_ram_ix167_a_110__dup_2543), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8058 (.Q (
                         modgen_ram_ix167_a_109__dup_2544), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2536), .SI (
                         modgen_ram_ix167_a_109__dup_2544), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8062 (.Q (
                         modgen_ram_ix167_a_108__dup_2545), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2518), .SI (
                         modgen_ram_ix167_a_108__dup_2545), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8066 (.Q (
                         modgen_ram_ix167_a_107__dup_2546), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2492), .SI (
                         modgen_ram_ix167_a_107__dup_2546), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8070 (.Q (
                         modgen_ram_ix167_a_106__dup_2547), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2474), .SI (
                         modgen_ram_ix167_a_106__dup_2547), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8074 (.Q (
                         modgen_ram_ix167_a_105__dup_2548), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2452), .SI (
                         modgen_ram_ix167_a_105__dup_2548), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8078 (.Q (
                         modgen_ram_ix167_a_104__dup_2549), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2434), .SI (
                         modgen_ram_ix167_a_104__dup_2549), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8082 (.Q (
                         modgen_ram_ix167_a_103__dup_2550), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2404), .SI (
                         modgen_ram_ix167_a_103__dup_2550), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8086 (.Q (
                         modgen_ram_ix167_a_102__dup_2551), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2386), .SI (
                         modgen_ram_ix167_a_102__dup_2551), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8090 (.Q (
                         modgen_ram_ix167_a_101__dup_2552), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2364), .SI (
                         modgen_ram_ix167_a_101__dup_2552), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8094 (.Q (
                         modgen_ram_ix167_a_100__dup_2553), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2346), .SI (
                         modgen_ram_ix167_a_100__dup_2553), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8098 (.Q (
                         modgen_ram_ix167_a_99__dup_2554), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2320), .SI (
                         modgen_ram_ix167_a_99__dup_2554), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8102 (.Q (
                         modgen_ram_ix167_a_98__dup_2555), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2302), .SI (
                         modgen_ram_ix167_a_98__dup_2555), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8106 (.Q (
                         modgen_ram_ix167_a_97__dup_2556), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2280), .SI (
                         modgen_ram_ix167_a_97__dup_2556), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8110 (.Q (
                         modgen_ram_ix167_a_96__dup_2557), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2262), .SI (
                         modgen_ram_ix167_a_96__dup_2557), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8114 (.Q (
                         modgen_ram_ix167_a_95__dup_2558), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2222), .SI (
                         modgen_ram_ix167_a_95__dup_2558), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8118 (.Q (
                         modgen_ram_ix167_a_94__dup_2559), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2204), .SI (
                         modgen_ram_ix167_a_94__dup_2559), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8122 (.Q (
                         modgen_ram_ix167_a_93__dup_2560), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2182), .SI (
                         modgen_ram_ix167_a_93__dup_2560), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8126 (.Q (
                         modgen_ram_ix167_a_92__dup_2561), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2164), .SI (
                         modgen_ram_ix167_a_92__dup_2561), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8130 (.Q (
                         modgen_ram_ix167_a_91__dup_2562), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2138), .SI (
                         modgen_ram_ix167_a_91__dup_2562), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8134 (.Q (
                         modgen_ram_ix167_a_90__dup_2563), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2120), .SI (
                         modgen_ram_ix167_a_90__dup_2563), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8138 (.Q (
                         modgen_ram_ix167_a_89__dup_2564), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2098), .SI (
                         modgen_ram_ix167_a_89__dup_2564), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8142 (.Q (
                         modgen_ram_ix167_a_88__dup_2565), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2080), .SI (
                         modgen_ram_ix167_a_88__dup_2565), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8146 (.Q (
                         modgen_ram_ix167_a_87__dup_2566), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2050), .SI (
                         modgen_ram_ix167_a_87__dup_2566), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8150 (.Q (
                         modgen_ram_ix167_a_86__dup_2567), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2032), .SI (
                         modgen_ram_ix167_a_86__dup_2567), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8154 (.Q (
                         modgen_ram_ix167_a_85__dup_2568), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx2010), .SI (
                         modgen_ram_ix167_a_85__dup_2568), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8158 (.Q (
                         modgen_ram_ix167_a_84__dup_2569), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1992), .SI (
                         modgen_ram_ix167_a_84__dup_2569), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8162 (.Q (
                         modgen_ram_ix167_a_83__dup_2570), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1966), .SI (
                         modgen_ram_ix167_a_83__dup_2570), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8166 (.Q (
                         modgen_ram_ix167_a_82__dup_2571), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1948), .SI (
                         modgen_ram_ix167_a_82__dup_2571), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8170 (.Q (
                         modgen_ram_ix167_a_81__dup_2572), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1926), .SI (
                         modgen_ram_ix167_a_81__dup_2572), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8174 (.Q (
                         modgen_ram_ix167_a_80__dup_2573), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1908), .SI (
                         modgen_ram_ix167_a_80__dup_2573), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8178 (.Q (
                         modgen_ram_ix167_a_79__dup_2574), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1872), .SI (
                         modgen_ram_ix167_a_79__dup_2574), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8182 (.Q (
                         modgen_ram_ix167_a_78__dup_2575), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1854), .SI (
                         modgen_ram_ix167_a_78__dup_2575), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8186 (.Q (
                         modgen_ram_ix167_a_77__dup_2576), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1832), .SI (
                         modgen_ram_ix167_a_77__dup_2576), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8190 (.Q (
                         modgen_ram_ix167_a_76__dup_2577), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1814), .SI (
                         modgen_ram_ix167_a_76__dup_2577), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8194 (.Q (
                         modgen_ram_ix167_a_75__dup_2578), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1788), .SI (
                         modgen_ram_ix167_a_75__dup_2578), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8198 (.Q (
                         modgen_ram_ix167_a_74__dup_2579), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1770), .SI (
                         modgen_ram_ix167_a_74__dup_2579), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8202 (.Q (
                         modgen_ram_ix167_a_73__dup_2580), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1748), .SI (
                         modgen_ram_ix167_a_73__dup_2580), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8206 (.Q (
                         modgen_ram_ix167_a_72__dup_2581), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1730), .SI (
                         modgen_ram_ix167_a_72__dup_2581), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8210 (.Q (
                         modgen_ram_ix167_a_71__dup_2582), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1700), .SI (
                         modgen_ram_ix167_a_71__dup_2582), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8214 (.Q (
                         modgen_ram_ix167_a_70__dup_2583), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1682), .SI (
                         modgen_ram_ix167_a_70__dup_2583), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8218 (.Q (
                         modgen_ram_ix167_a_69__dup_2584), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1660), .SI (
                         modgen_ram_ix167_a_69__dup_2584), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8222 (.Q (
                         modgen_ram_ix167_a_68__dup_2585), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1642), .SI (
                         modgen_ram_ix167_a_68__dup_2585), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8226 (.Q (
                         modgen_ram_ix167_a_67__dup_2586), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1616), .SI (
                         modgen_ram_ix167_a_67__dup_2586), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8230 (.Q (
                         modgen_ram_ix167_a_66__dup_2587), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1598), .SI (
                         modgen_ram_ix167_a_66__dup_2587), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8234 (.Q (
                         modgen_ram_ix167_a_65__dup_2588), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1576), .SI (
                         modgen_ram_ix167_a_65__dup_2588), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8238 (.Q (
                         modgen_ram_ix167_a_64__dup_2589), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1558), .SI (
                         modgen_ram_ix167_a_64__dup_2589), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8242 (.Q (
                         modgen_ram_ix167_a_63__dup_2590), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1510), .SI (
                         modgen_ram_ix167_a_63__dup_2590), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8246 (.Q (
                         modgen_ram_ix167_a_62__dup_2591), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1492), .SI (
                         modgen_ram_ix167_a_62__dup_2591), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8250 (.Q (
                         modgen_ram_ix167_a_61__dup_2592), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1470), .SI (
                         modgen_ram_ix167_a_61__dup_2592), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8254 (.Q (
                         modgen_ram_ix167_a_60__dup_2593), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1452), .SI (
                         modgen_ram_ix167_a_60__dup_2593), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8258 (.Q (
                         modgen_ram_ix167_a_59__dup_2594), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1426), .SI (
                         modgen_ram_ix167_a_59__dup_2594), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8262 (.Q (
                         modgen_ram_ix167_a_58__dup_2595), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1408), .SI (
                         modgen_ram_ix167_a_58__dup_2595), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8266 (.Q (
                         modgen_ram_ix167_a_57__dup_2596), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1386), .SI (
                         modgen_ram_ix167_a_57__dup_2596), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8270 (.Q (
                         modgen_ram_ix167_a_56__dup_2597), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1368), .SI (
                         modgen_ram_ix167_a_56__dup_2597), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8274 (.Q (
                         modgen_ram_ix167_a_55__dup_2598), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1338), .SI (
                         modgen_ram_ix167_a_55__dup_2598), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8278 (.Q (
                         modgen_ram_ix167_a_54__dup_2599), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1320), .SI (
                         modgen_ram_ix167_a_54__dup_2599), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8282 (.Q (
                         modgen_ram_ix167_a_53__dup_2600), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1298), .SI (
                         modgen_ram_ix167_a_53__dup_2600), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8286 (.Q (
                         modgen_ram_ix167_a_52__dup_2601), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1280), .SI (
                         modgen_ram_ix167_a_52__dup_2601), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8290 (.Q (
                         modgen_ram_ix167_a_51__dup_2602), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1254), .SI (
                         modgen_ram_ix167_a_51__dup_2602), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8294 (.Q (
                         modgen_ram_ix167_a_50__dup_2603), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1236), .SI (
                         modgen_ram_ix167_a_50__dup_2603), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8298 (.Q (
                         modgen_ram_ix167_a_49__dup_2604), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1214), .SI (
                         modgen_ram_ix167_a_49__dup_2604), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8302 (.Q (
                         modgen_ram_ix167_a_48__dup_2605), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1196), .SI (
                         modgen_ram_ix167_a_48__dup_2605), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8306 (.Q (
                         modgen_ram_ix167_a_47__dup_2606), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1154), .SI (
                         modgen_ram_ix167_a_47__dup_2606), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8310 (.Q (
                         modgen_ram_ix167_a_46__dup_2607), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1136), .SI (
                         modgen_ram_ix167_a_46__dup_2607), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8314 (.Q (
                         modgen_ram_ix167_a_45__dup_2608), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1114), .SI (
                         modgen_ram_ix167_a_45__dup_2608), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8318 (.Q (
                         modgen_ram_ix167_a_44__dup_2609), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1096), .SI (
                         modgen_ram_ix167_a_44__dup_2609), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8322 (.Q (
                         modgen_ram_ix167_a_43__dup_2610), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1070), .SI (
                         modgen_ram_ix167_a_43__dup_2610), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8326 (.Q (
                         modgen_ram_ix167_a_42__dup_2611), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1052), .SI (
                         modgen_ram_ix167_a_42__dup_2611), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8330 (.Q (
                         modgen_ram_ix167_a_41__dup_2612), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1030), .SI (
                         modgen_ram_ix167_a_41__dup_2612), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8334 (.Q (
                         modgen_ram_ix167_a_40__dup_2613), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx1012), .SI (
                         modgen_ram_ix167_a_40__dup_2613), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8338 (.Q (
                         modgen_ram_ix167_a_39__dup_2614), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx982), .SI (
                         modgen_ram_ix167_a_39__dup_2614), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8342 (.Q (
                         modgen_ram_ix167_a_38__dup_2615), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx964), .SI (
                         modgen_ram_ix167_a_38__dup_2615), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8346 (.Q (
                         modgen_ram_ix167_a_37__dup_2616), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx942), .SI (
                         modgen_ram_ix167_a_37__dup_2616), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8350 (.Q (
                         modgen_ram_ix167_a_36__dup_2617), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx924), .SI (
                         modgen_ram_ix167_a_36__dup_2617), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8354 (.Q (
                         modgen_ram_ix167_a_35__dup_2618), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx898), .SI (
                         modgen_ram_ix167_a_35__dup_2618), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8358 (.Q (
                         modgen_ram_ix167_a_34__dup_2619), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx880), .SI (
                         modgen_ram_ix167_a_34__dup_2619), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8362 (.Q (
                         modgen_ram_ix167_a_33__dup_2620), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx858), .SI (
                         modgen_ram_ix167_a_33__dup_2620), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8366 (.Q (
                         modgen_ram_ix167_a_32__dup_2621), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx840), .SI (
                         modgen_ram_ix167_a_32__dup_2621), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8370 (.Q (
                         modgen_ram_ix167_a_31__dup_2622), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx796), .SI (
                         modgen_ram_ix167_a_31__dup_2622), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8374 (.Q (
                         modgen_ram_ix167_a_30__dup_2623), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx778), .SI (
                         modgen_ram_ix167_a_30__dup_2623), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8378 (.Q (
                         modgen_ram_ix167_a_29__dup_2624), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx756), .SI (
                         modgen_ram_ix167_a_29__dup_2624), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8382 (.Q (
                         modgen_ram_ix167_a_28__dup_2625), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx738), .SI (
                         modgen_ram_ix167_a_28__dup_2625), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8386 (.Q (
                         modgen_ram_ix167_a_27__dup_2626), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx712), .SI (
                         modgen_ram_ix167_a_27__dup_2626), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8390 (.Q (
                         modgen_ram_ix167_a_26__dup_2627), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx694), .SI (
                         modgen_ram_ix167_a_26__dup_2627), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8394 (.Q (
                         modgen_ram_ix167_a_25__dup_2628), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx672), .SI (
                         modgen_ram_ix167_a_25__dup_2628), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8398 (.Q (
                         modgen_ram_ix167_a_24__dup_2629), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx654), .SI (
                         modgen_ram_ix167_a_24__dup_2629), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8402 (.Q (
                         modgen_ram_ix167_a_23__dup_2630), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx624), .SI (
                         modgen_ram_ix167_a_23__dup_2630), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8406 (.Q (
                         modgen_ram_ix167_a_22__dup_2631), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx606), .SI (
                         modgen_ram_ix167_a_22__dup_2631), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8410 (.Q (
                         modgen_ram_ix167_a_21__dup_2632), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx584), .SI (
                         modgen_ram_ix167_a_21__dup_2632), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8414 (.Q (
                         modgen_ram_ix167_a_20__dup_2633), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx566), .SI (
                         modgen_ram_ix167_a_20__dup_2633), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8418 (.Q (
                         modgen_ram_ix167_a_19__dup_2634), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx540), .SI (
                         modgen_ram_ix167_a_19__dup_2634), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8422 (.Q (
                         modgen_ram_ix167_a_18__dup_2635), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx522), .SI (
                         modgen_ram_ix167_a_18__dup_2635), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8426 (.Q (
                         modgen_ram_ix167_a_17__dup_2636), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx500), .SI (
                         modgen_ram_ix167_a_17__dup_2636), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8430 (.Q (
                         modgen_ram_ix167_a_16__dup_2637), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx482), .SI (
                         modgen_ram_ix167_a_16__dup_2637), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8434 (.Q (
                         modgen_ram_ix167_a_15__dup_2638), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx442), .SI (
                         modgen_ram_ix167_a_15__dup_2638), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8438 (.Q (
                         modgen_ram_ix167_a_14__dup_2639), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx422), .SI (
                         modgen_ram_ix167_a_14__dup_2639), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8442 (.Q (
                         modgen_ram_ix167_a_13__dup_2640), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx398), .SI (
                         modgen_ram_ix167_a_13__dup_2640), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8446 (.Q (
                         modgen_ram_ix167_a_12__dup_2641), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx378), .SI (
                         modgen_ram_ix167_a_12__dup_2641), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8450 (.Q (
                         modgen_ram_ix167_a_11__dup_2642), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx344), .SI (
                         modgen_ram_ix167_a_11__dup_2642), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8454 (.Q (
                         modgen_ram_ix167_a_10__dup_2643), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx324), .SI (
                         modgen_ram_ix167_a_10__dup_2643), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8458 (.Q (
                         modgen_ram_ix167_a_9__dup_2644), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx340), .SI (
                         modgen_ram_ix167_a_9__dup_2644), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8462 (.Q (
                         modgen_ram_ix167_a_8__dup_2645), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx280), .SI (
                         modgen_ram_ix167_a_8__dup_2645), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8466 (.Q (
                         modgen_ram_ix167_a_7__dup_2646), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx244), .SI (
                         modgen_ram_ix167_a_7__dup_2646), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8470 (.Q (
                         modgen_ram_ix167_a_6__dup_2647), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx224), .SI (
                         modgen_ram_ix167_a_6__dup_2647), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8474 (.Q (
                         modgen_ram_ix167_a_5__dup_2648), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx200), .SI (
                         modgen_ram_ix167_a_5__dup_2648), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8478 (.Q (
                         modgen_ram_ix167_a_4__dup_2649), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx180), .SI (
                         modgen_ram_ix167_a_4__dup_2649), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8482 (.Q (
                         modgen_ram_ix167_a_3__dup_2650), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx148), .SI (
                         modgen_ram_ix167_a_3__dup_2650), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8486 (.Q (
                         modgen_ram_ix167_a_2__dup_2651), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (nx3519), .SI (
                         modgen_ram_ix167_a_2__dup_2651), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8490 (.Q (
                         modgen_ram_ix167_a_1__dup_2652), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (nx3520), .SI (
                         modgen_ram_ix167_a_1__dup_2652), .SN (nx28503)) ;
    SDFFSRPQ_X0P5M_A12TS modgen_ram_ix167_ix8494 (.Q (
                         modgen_ram_ix167_a_0__dup_2653), .CK (wb_clk_i), .D (
                         nx28523), .R (nx3204), .SE (NOT_nx70), .SI (
                         modgen_ram_ix167_a_0__dup_2653), .SN (nx28503)) ;
    INV_X13M_A12TS ix28496 (.Y (nx28497), .A (nx3204)) ;
    INV_X13M_A12TS ix28498 (.Y (nx28499), .A (nx3204)) ;
    INV_X13M_A12TS ix28500 (.Y (nx28501), .A (nx3204)) ;
    INV_X13M_A12TS ix28502 (.Y (nx28503), .A (nx3204)) ;
    OR3_X0P5M_A12TS ix5765 (.Y (NOT_nx5764), .A (nx3225), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5747 (.Y (NOT_nx5746), .A (nx3224), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix3038 (.Y (NOT_nx5724), .A (nx390), .B (nx3286), .C (nx5442
                    )) ;
    OR3_X0P5M_A12TS ix5707 (.Y (NOT_nx5706), .A (nx3223), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5681 (.Y (NOT_nx5680), .A (nx336), .B (nx3286), .C (nx5442
                    )) ;
    OR3_X0P5M_A12TS ix5663 (.Y (NOT_nx5662), .A (nx316), .B (nx3286), .C (nx5442
                    )) ;
    OR3_X0P5M_A12TS ix5641 (.Y (NOT_nx5640), .A (nx292), .B (nx3286), .C (nx5442
                    )) ;
    OR3_X0P5M_A12TS ix5623 (.Y (NOT_nx5622), .A (nx3220), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5593 (.Y (NOT_nx5592), .A (nx3218), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5575 (.Y (NOT_nx5574), .A (nx3217), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5553 (.Y (NOT_nx5552), .A (nx3216), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5535 (.Y (NOT_nx5534), .A (nx172), .B (nx3286), .C (nx5442
                    )) ;
    OR3_X0P5M_A12TS ix5509 (.Y (NOT_nx5508), .A (nx140), .B (nx3286), .C (nx5442
                    )) ;
    OR3_X0P5M_A12TS ix5491 (.Y (NOT_nx5490), .A (nx3215), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5469 (.Y (NOT_nx5468), .A (nx3214), .B (nx3286), .C (
                    nx5442)) ;
    OR3_X0P5M_A12TS ix5451 (.Y (NOT_nx5450), .A (nx62), .B (nx3286), .C (nx5442)
                    ) ;
    OR3_X0P5M_A12TS ix5415 (.Y (NOT_nx5414), .A (nx5092), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix5397 (.Y (NOT_nx5396), .A (nx5092), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix5375 (.Y (NOT_nx5374), .A (nx5092), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix5357 (.Y (NOT_nx5356), .A (nx5092), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix5331 (.Y (NOT_nx5330), .A (nx5092), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix5313 (.Y (NOT_nx5312), .A (nx5092), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix5291 (.Y (NOT_nx5290), .A (nx5092), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix5273 (.Y (NOT_nx5272), .A (nx5092), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix5243 (.Y (NOT_nx5242), .A (nx5092), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix5225 (.Y (NOT_nx5224), .A (nx5092), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix5203 (.Y (NOT_nx5202), .A (nx5092), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix5185 (.Y (NOT_nx5184), .A (nx5092), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix5159 (.Y (NOT_nx5158), .A (nx5092), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix5141 (.Y (NOT_nx5140), .A (nx5092), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix5119 (.Y (NOT_nx5118), .A (nx5092), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix5101 (.Y (NOT_nx5100), .A (nx5092), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix5061 (.Y (NOT_nx5060), .A (nx4738), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix5043 (.Y (NOT_nx5042), .A (nx4738), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix5021 (.Y (NOT_nx5020), .A (nx4738), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix5003 (.Y (NOT_nx5002), .A (nx4738), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix4977 (.Y (NOT_nx4976), .A (nx4738), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix4959 (.Y (NOT_nx4958), .A (nx4738), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix4937 (.Y (NOT_nx4936), .A (nx4738), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3039 (.Y (NOT_nx4918), .A (nx4738), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix4889 (.Y (NOT_nx4888), .A (nx4738), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix4871 (.Y (NOT_nx4870), .A (nx4738), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix4849 (.Y (NOT_nx4848), .A (nx4738), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3040 (.Y (NOT_nx4830), .A (nx4738), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix4805 (.Y (NOT_nx4804), .A (nx4738), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix4787 (.Y (NOT_nx4786), .A (nx4738), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix4765 (.Y (NOT_nx4764), .A (nx4738), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix4747 (.Y (NOT_nx4746), .A (nx4738), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3041 (.Y (NOT_nx4710), .A (nx3263), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3042 (.Y (NOT_nx4692), .A (nx3263), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3044 (.Y (NOT_nx4670), .A (nx3263), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix4653 (.Y (NOT_nx4652), .A (nx3263), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3045 (.Y (NOT_nx4626), .A (nx3263), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3046 (.Y (NOT_nx4608), .A (nx3263), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix4587 (.Y (NOT_nx4586), .A (nx3263), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix4569 (.Y (NOT_nx4568), .A (nx3263), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3047 (.Y (NOT_nx4538), .A (nx3263), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix4521 (.Y (NOT_nx4520), .A (nx3263), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3048 (.Y (NOT_nx4498), .A (nx3263), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix4481 (.Y (NOT_nx4480), .A (nx3263), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix4455 (.Y (NOT_nx4454), .A (nx3263), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3049 (.Y (NOT_nx4436), .A (nx3263), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix4415 (.Y (NOT_nx4414), .A (nx3263), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix4397 (.Y (NOT_nx4396), .A (nx3263), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3050 (.Y (NOT_nx4346), .A (nx4024), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix4329 (.Y (NOT_nx4328), .A (nx4024), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3051 (.Y (NOT_nx4306), .A (nx4024), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3052 (.Y (NOT_nx4288), .A (nx4024), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix4263 (.Y (NOT_nx4262), .A (nx4024), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix4245 (.Y (NOT_nx4244), .A (nx4024), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix4223 (.Y (NOT_nx4222), .A (nx4024), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3053 (.Y (NOT_nx4204), .A (nx4024), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix4175 (.Y (NOT_nx4174), .A (nx4024), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix4157 (.Y (NOT_nx4156), .A (nx4024), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix4135 (.Y (NOT_nx4134), .A (nx4024), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix4117 (.Y (NOT_nx4116), .A (nx4024), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix4091 (.Y (NOT_nx4090), .A (nx4024), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3054 (.Y (NOT_nx4072), .A (nx4024), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix4051 (.Y (NOT_nx4050), .A (nx4024), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix4033 (.Y (NOT_nx4032), .A (nx4024), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3997 (.Y (NOT_nx3996), .A (nx3674), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3979 (.Y (NOT_nx3978), .A (nx3674), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3957 (.Y (NOT_nx3956), .A (nx3674), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3939 (.Y (NOT_nx3938), .A (nx3674), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3913 (.Y (NOT_nx3912), .A (nx3674), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3056 (.Y (NOT_nx3894), .A (nx3674), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3057 (.Y (NOT_nx3872), .A (nx3674), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3855 (.Y (NOT_nx3854), .A (nx3674), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3825 (.Y (NOT_nx3824), .A (nx3674), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3807 (.Y (NOT_nx3806), .A (nx3674), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3785 (.Y (NOT_nx3784), .A (nx3674), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3767 (.Y (NOT_nx3766), .A (nx3674), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3058 (.Y (NOT_nx3740), .A (nx3674), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3723 (.Y (NOT_nx3722), .A (nx3674), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3060 (.Y (NOT_nx3700), .A (nx3674), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3683 (.Y (NOT_nx3682), .A (nx3674), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3643 (.Y (NOT_nx3642), .A (nx3320), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3061 (.Y (NOT_nx3624), .A (nx3320), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3603 (.Y (NOT_nx3602), .A (nx3320), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3585 (.Y (NOT_nx3584), .A (nx3320), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3559 (.Y (NOT_nx3558), .A (nx3320), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3541 (.Y (NOT_nx3540), .A (nx3320), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3519 (.Y (NOT_nx3518), .A (nx3320), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3501 (.Y (NOT_nx3500), .A (nx3320), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3471 (.Y (NOT_nx3470), .A (nx3320), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3453 (.Y (NOT_nx3452), .A (nx3320), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3431 (.Y (NOT_nx3430), .A (nx3320), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3413 (.Y (NOT_nx3412), .A (nx3320), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3387 (.Y (NOT_nx3386), .A (nx3320), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3062 (.Y (NOT_nx3368), .A (nx3320), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3347 (.Y (NOT_nx3346), .A (nx3320), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3329 (.Y (NOT_nx3328), .A (nx3320), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3293 (.Y (NOT_nx3292), .A (nx2970), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3063 (.Y (NOT_nx3274), .A (nx2970), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3253 (.Y (NOT_nx3252), .A (nx2970), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3064 (.Y (NOT_nx3234), .A (nx2970), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3209 (.Y (NOT_nx3208), .A (nx2970), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3191 (.Y (NOT_nx3190), .A (nx2970), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3065 (.Y (NOT_nx3168), .A (nx2970), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3151 (.Y (NOT_nx3150), .A (nx2970), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3121 (.Y (NOT_nx3120), .A (nx2970), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3103 (.Y (NOT_nx3102), .A (nx2970), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3081 (.Y (NOT_nx3080), .A (nx2970), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3066 (.Y (NOT_nx3062), .A (nx2970), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3067 (.Y (NOT_nx3036), .A (nx2970), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3068 (.Y (NOT_nx3018), .A (nx2970), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3070 (.Y (NOT_nx2996), .A (nx2970), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3071 (.Y (NOT_nx2978), .A (nx2970), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3072 (.Y (NOT_nx2926), .A (nx3257), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3073 (.Y (NOT_nx2908), .A (nx3257), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3074 (.Y (NOT_nx2886), .A (nx3257), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3075 (.Y (NOT_nx2868), .A (nx3257), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3076 (.Y (NOT_nx2842), .A (nx3257), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3078 (.Y (NOT_nx2824), .A (nx3257), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3079 (.Y (NOT_nx2802), .A (nx3257), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3080 (.Y (NOT_nx2784), .A (nx3257), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3082 (.Y (NOT_nx2754), .A (nx3257), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3084 (.Y (NOT_nx2736), .A (nx3257), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3085 (.Y (NOT_nx2714), .A (nx3257), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3086 (.Y (NOT_nx2696), .A (nx3257), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3087 (.Y (NOT_nx2670), .A (nx3257), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3088 (.Y (NOT_nx2652), .A (nx3257), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3090 (.Y (NOT_nx2630), .A (nx3257), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3091 (.Y (NOT_nx2612), .A (nx3257), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3092 (.Y (NOT_nx2576), .A (nx3250), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3093 (.Y (NOT_nx2558), .A (nx3250), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3094 (.Y (NOT_nx2536), .A (nx3250), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3095 (.Y (NOT_nx2518), .A (nx3250), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3096 (.Y (NOT_nx2492), .A (nx3250), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3097 (.Y (NOT_nx2474), .A (nx3250), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3098 (.Y (NOT_nx2452), .A (nx3250), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3099 (.Y (NOT_nx2434), .A (nx3250), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix2405 (.Y (NOT_nx2404), .A (nx3250), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix2387 (.Y (NOT_nx2386), .A (nx3250), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix2365 (.Y (NOT_nx2364), .A (nx3250), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix2347 (.Y (NOT_nx2346), .A (nx3250), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3100 (.Y (NOT_nx2320), .A (nx3250), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3102 (.Y (NOT_nx2302), .A (nx3250), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3104 (.Y (NOT_nx2280), .A (nx3250), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3105 (.Y (NOT_nx2262), .A (nx3250), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3106 (.Y (NOT_nx2222), .A (nx3247), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3107 (.Y (NOT_nx2204), .A (nx3247), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3108 (.Y (NOT_nx2182), .A (nx3247), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix3109 (.Y (NOT_nx2164), .A (nx3247), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix2139 (.Y (NOT_nx2138), .A (nx3247), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3110 (.Y (NOT_nx2120), .A (nx3247), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3111 (.Y (NOT_nx2098), .A (nx3247), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix2081 (.Y (NOT_nx2080), .A (nx3247), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix2051 (.Y (NOT_nx2050), .A (nx3247), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3112 (.Y (NOT_nx2032), .A (nx3247), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3113 (.Y (NOT_nx2010), .A (nx3247), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3114 (.Y (NOT_nx1992), .A (nx3247), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3115 (.Y (NOT_nx1966), .A (nx3247), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3116 (.Y (NOT_nx1948), .A (nx3247), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3118 (.Y (NOT_nx1926), .A (nx3247), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix1909 (.Y (NOT_nx1908), .A (nx3247), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3119 (.Y (NOT_nx1872), .A (nx1550), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3120 (.Y (NOT_nx1854), .A (nx1550), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix1833 (.Y (NOT_nx1832), .A (nx1550), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix1815 (.Y (NOT_nx1814), .A (nx1550), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix1789 (.Y (NOT_nx1788), .A (nx1550), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3122 (.Y (NOT_nx1770), .A (nx1550), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3124 (.Y (NOT_nx1748), .A (nx1550), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3125 (.Y (NOT_nx1730), .A (nx1550), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3126 (.Y (NOT_nx1700), .A (nx1550), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3127 (.Y (NOT_nx1682), .A (nx1550), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3128 (.Y (NOT_nx1660), .A (nx1550), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3129 (.Y (NOT_nx1642), .A (nx1550), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3130 (.Y (NOT_nx1616), .A (nx1550), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix3131 (.Y (NOT_nx1598), .A (nx1550), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3132 (.Y (NOT_nx1576), .A (nx1550), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3133 (.Y (NOT_nx1558), .A (nx1550), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3134 (.Y (NOT_nx1510), .A (nx3239), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix1493 (.Y (NOT_nx1492), .A (nx3239), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix1471 (.Y (NOT_nx1470), .A (nx3239), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix1453 (.Y (NOT_nx1452), .A (nx3239), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix1427 (.Y (NOT_nx1426), .A (nx3239), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3136 (.Y (NOT_nx1408), .A (nx3239), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3137 (.Y (NOT_nx1386), .A (nx3239), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix1369 (.Y (NOT_nx1368), .A (nx3239), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix3138 (.Y (NOT_nx1338), .A (nx3239), .B (nx3286), .C (
                    nx3218)) ;
    OR3_X0P5M_A12TS ix3140 (.Y (NOT_nx1320), .A (nx3239), .B (nx3286), .C (
                    nx3217)) ;
    OR3_X0P5M_A12TS ix3141 (.Y (NOT_nx1298), .A (nx3239), .B (nx3286), .C (
                    nx3216)) ;
    OR3_X0P5M_A12TS ix3142 (.Y (NOT_nx1280), .A (nx3239), .B (nx3286), .C (nx172
                    )) ;
    OR3_X0P5M_A12TS ix3143 (.Y (NOT_nx1254), .A (nx3239), .B (nx3286), .C (nx140
                    )) ;
    OR3_X0P5M_A12TS ix1237 (.Y (NOT_nx1236), .A (nx3239), .B (nx3286), .C (
                    nx3215)) ;
    OR3_X0P5M_A12TS ix3144 (.Y (NOT_nx1214), .A (nx3239), .B (nx3286), .C (
                    nx3214)) ;
    OR3_X0P5M_A12TS ix3145 (.Y (NOT_nx1196), .A (nx3239), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix1155 (.Y (NOT_nx1154), .A (nx3231), .B (nx3286), .C (
                    nx3225)) ;
    OR3_X0P5M_A12TS ix3146 (.Y (NOT_nx1136), .A (nx3231), .B (nx3286), .C (
                    nx3224)) ;
    OR3_X0P5M_A12TS ix3148 (.Y (NOT_nx1114), .A (nx3231), .B (nx3286), .C (nx390
                    )) ;
    OR3_X0P5M_A12TS ix1097 (.Y (NOT_nx1096), .A (nx3231), .B (nx3286), .C (
                    nx3223)) ;
    OR3_X0P5M_A12TS ix3149 (.Y (NOT_nx1070), .A (nx3231), .B (nx3286), .C (nx336
                    )) ;
    OR3_X0P5M_A12TS ix3150 (.Y (NOT_nx1052), .A (nx3231), .B (nx3286), .C (nx316
                    )) ;
    OR3_X0P5M_A12TS ix3152 (.Y (NOT_nx1030), .A (nx3231), .B (nx3286), .C (nx292
                    )) ;
    OR3_X0P5M_A12TS ix3153 (.Y (NOT_nx1012), .A (nx3231), .B (nx3286), .C (
                    nx3220)) ;
    OR3_X0P5M_A12TS ix983 (.Y (NOT_nx982), .A (nx3231), .B (nx3286), .C (nx3218)
                    ) ;
    OR3_X0P5M_A12TS ix3154 (.Y (NOT_nx964), .A (nx3231), .B (nx3286), .C (nx3217
                    )) ;
    OR3_X0P5M_A12TS ix3155 (.Y (NOT_nx942), .A (nx3231), .B (nx3286), .C (nx3216
                    )) ;
    OR3_X0P5M_A12TS ix3156 (.Y (NOT_nx924), .A (nx3231), .B (nx3286), .C (nx172)
                    ) ;
    OR3_X0P5M_A12TS ix3158 (.Y (NOT_nx898), .A (nx3231), .B (nx3286), .C (nx140)
                    ) ;
    OR3_X0P5M_A12TS ix3160 (.Y (NOT_nx880), .A (nx3231), .B (nx3286), .C (nx3215
                    )) ;
    OR3_X0P5M_A12TS ix3161 (.Y (NOT_nx858), .A (nx3231), .B (nx3286), .C (nx3214
                    )) ;
    OR3_X0P5M_A12TS ix841 (.Y (NOT_nx840), .A (nx3231), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3162 (.Y (NOT_nx796), .A (nx3227), .B (nx3286), .C (nx3225
                    )) ;
    OR3_X0P5M_A12TS ix3163 (.Y (NOT_nx778), .A (nx3227), .B (nx3286), .C (nx3224
                    )) ;
    OR3_X0P5M_A12TS ix3164 (.Y (NOT_nx756), .A (nx3227), .B (nx3286), .C (nx390)
                    ) ;
    OR3_X0P5M_A12TS ix739 (.Y (NOT_nx738), .A (nx3227), .B (nx3286), .C (nx3223)
                    ) ;
    OR3_X0P5M_A12TS ix713 (.Y (NOT_nx712), .A (nx3227), .B (nx3286), .C (nx336)
                    ) ;
    OR3_X0P5M_A12TS ix3165 (.Y (NOT_nx694), .A (nx3227), .B (nx3286), .C (nx316)
                    ) ;
    OR3_X0P5M_A12TS ix673 (.Y (NOT_nx672), .A (nx3227), .B (nx3286), .C (nx292)
                    ) ;
    OR3_X0P5M_A12TS ix655 (.Y (NOT_nx654), .A (nx3227), .B (nx3286), .C (nx3220)
                    ) ;
    OR3_X0P5M_A12TS ix3166 (.Y (NOT_nx624), .A (nx3227), .B (nx3286), .C (nx3218
                    )) ;
    OR3_X0P5M_A12TS ix607 (.Y (NOT_nx606), .A (nx3227), .B (nx3286), .C (nx3217)
                    ) ;
    OR3_X0P5M_A12TS ix585 (.Y (NOT_nx584), .A (nx3227), .B (nx3286), .C (nx3216)
                    ) ;
    OR3_X0P5M_A12TS ix567 (.Y (NOT_nx566), .A (nx3227), .B (nx3286), .C (nx172)
                    ) ;
    OR3_X0P5M_A12TS ix3167 (.Y (NOT_nx540), .A (nx3227), .B (nx3286), .C (nx140)
                    ) ;
    OR3_X0P5M_A12TS ix523 (.Y (NOT_nx522), .A (nx3227), .B (nx3286), .C (nx3215)
                    ) ;
    OR3_X0P5M_A12TS ix3168 (.Y (NOT_nx500), .A (nx3227), .B (nx3286), .C (nx3214
                    )) ;
    OR3_X0P5M_A12TS ix3170 (.Y (NOT_nx482), .A (nx3227), .B (nx3286), .C (nx62)
                    ) ;
    OR3_X0P5M_A12TS ix3171 (.Y (NOT_nx442), .A (nx3213), .B (nx3286), .C (nx3225
                    )) ;
    OR3_X0P5M_A12TS ix3172 (.Y (NOT_nx422), .A (nx3213), .B (nx3286), .C (nx3224
                    )) ;
    OR3_X0P5M_A12TS ix3173 (.Y (NOT_nx398), .A (nx3213), .B (nx3286), .C (nx390)
                    ) ;
    OR3_X0P5M_A12TS ix3174 (.Y (NOT_nx378), .A (nx3213), .B (nx3286), .C (nx3223
                    )) ;
    OR3_X0P5M_A12TS ix345 (.Y (NOT_nx344), .A (nx3213), .B (nx3286), .C (nx336)
                    ) ;
    OR3_X0P5M_A12TS ix3175 (.Y (NOT_nx324), .A (nx3213), .B (nx3286), .C (nx316)
                    ) ;
    OR3_X0P5M_A12TS ix3176 (.Y (NOT_nx340), .A (nx3213), .B (nx3286), .C (nx292)
                    ) ;
    OR3_X0P5M_A12TS ix3177 (.Y (NOT_nx280), .A (nx3213), .B (nx3286), .C (nx3220
                    )) ;
    OR3_X0P5M_A12TS ix3178 (.Y (NOT_nx244), .A (nx3213), .B (nx3286), .C (nx3218
                    )) ;
    OR3_X0P5M_A12TS ix3179 (.Y (NOT_nx224), .A (nx3213), .B (nx3286), .C (nx3217
                    )) ;
    OR3_X0P5M_A12TS ix3180 (.Y (NOT_nx200), .A (nx3213), .B (nx3286), .C (nx3216
                    )) ;
    OR3_X0P5M_A12TS ix3181 (.Y (NOT_nx180), .A (nx3213), .B (nx3286), .C (nx172)
                    ) ;
    OR3_X0P5M_A12TS ix3182 (.Y (NOT_nx148), .A (nx3213), .B (nx3286), .C (nx140)
                    ) ;
    OR3_X0P5M_A12TS ix3183 (.Y (nx3519), .A (nx3213), .B (nx3286), .C (nx3215)
                    ) ;
    OR3_X0P5M_A12TS ix3184 (.Y (nx3520), .A (nx3213), .B (nx3286), .C (nx3214)
                    ) ;
    OR3_X0P5M_A12TS ix3186 (.Y (NOT_nx70), .A (nx3213), .B (nx3286), .C (nx62)
                    ) ;
    INV_X3P5B_A12TS ix28508 (.Y (nx28509), .A (nx2755)) ;
    INV_X3P5B_A12TS ix28510 (.Y (nx28511), .A (nx2493)) ;
    INV_X3P5B_A12TS ix28512 (.Y (nx28513), .A (nx3454)) ;
    INV_X3P5B_A12TS ix28514 (.Y (nx28515), .A (nx3415)) ;
    INV_X3P5B_A12TS ix28516 (.Y (nx28517), .A (nx3374)) ;
    INV_X3P5B_A12TS ix28518 (.Y (nx28519), .A (nx1423)) ;
    INV_X3P5B_A12TS ix28520 (.Y (nx28521), .A (nx3326)) ;
    INV_X3P5B_A12TS ix28522 (.Y (nx28523), .A (nx863)) ;
    XOR2_X0P5M_A12TS ix3521 (.Y (p), .A (nx3597), .B (nx3614)) ;
    XNOR3_X0P5M_A12TS ix3522 (.Y (nx3597), .A (nx3590), .B (nx422), .C (nx3592)
                      ) ;
    XOR2_X0P5M_A12TS ix3523 (.Y (nx3590), .A (nx3581), .B (nx421)) ;
    OAI211_X0P5M_A12TS ix3524 (.Y (nx3581), .A0 (nx3587), .A1 (nx3598), .B0 (
                       nx477), .C0 (nx3608)) ;
    NAND2_X0P5A_A12TS ix75 (.Y (nx3587), .A (wr_addr_0), .B (wr_addr_1)) ;
    NAND3_X0P5A_A12TS ix3525 (.Y (nx3598), .A (nx3588), .B (desCy), .C (nx3606)
                      ) ;
    INV_X0P5B_A12TS ix3526 (.Y (nx3600), .A (wr_addr_3)) ;
    INV_X0P5B_A12TS ix3527 (.Y (nx3601), .A (wr_addr_2)) ;
    OAI22_X0P5M_A12TS ix3528 (.Y (nx3585), .A0 (wr_sfr_1), .A1 (nx457), .B0 (
                      nx3602), .B1 (nx3603)) ;
    INV_X0P5B_A12TS ix458 (.Y (nx457), .A (wr_sfr_0)) ;
    NAND4_X0P5A_A12TS ix3530 (.Y (nx3602), .A (wr_addr_7), .B (wr_addr_5), .C (
                      wr_addr_6), .D (nx3583)) ;
    NOR2_X0P5A_A12TS ix3531 (.Y (nx3583), .A (wr_addr_4), .B (wr_addr_3)) ;
    NOR2_X0P5A_A12TS ix3532 (.Y (nx3604), .A (wr_addr_0), .B (wr_addr_1)) ;
    OAI21_X0P5M_A12TS ix3533 (.Y (nx3606), .A0 (nx3607), .A1 (nx3601), .B0 (
                      nx3586)) ;
    NAND4B_X0P5M_A12TS ix3534 (.Y (nx3607), .AN (nx3599), .B (wr_bit_r_dup_1790)
                       , .C (nx3600), .D (we)) ;
    NOR2_X0P5A_A12TS ix3535 (.Y (nx3586), .A (nx3585), .B (nx3605)) ;
    AOI22_X0P5M_A12TS ix478 (.Y (nx477), .A0 (des2_7), .A1 (nx3605), .B0 (
                      des_acc_7), .B1 (nx100)) ;
    NOR2B_X0P7M_A12TS ix101 (.Y (nx100), .AN (nx3585), .B (nx3605)) ;
    AO21A1AI2_X0P5M_A12TS ix3536 (.Y (nx3608), .A0 (nx3587), .A1 (nx3586), .B0 (
                          nx68), .C0 (acc_7)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_7 (.Q (acc_7), .CK (wb_clk_i), .D (nx3581), 
                       .R (wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix3537 (.Y (nx421), .A0 (nx3589), .A1 (nx3598), .B0 (
                       nx3609), .C0 (nx3611)) ;
    AOI22_X0P5M_A12TS ix3538 (.Y (nx3609), .A0 (des2_6), .A1 (nx3605), .B0 (
                      des_acc_6), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix3539 (.Y (nx3611), .A0 (nx3589), .A1 (nx3586), .B0 (
                          nx68), .C0 (acc_6)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_6 (.Q (acc_6), .CK (wb_clk_i), .D (nx421), .R (
                       wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix3540 (.Y (nx422), .A0 (nx3591), .A1 (nx3598), .B0 (
                       nx497), .C0 (nx499)) ;
    AOI22_X0P5M_A12TS ix498 (.Y (nx497), .A0 (des2_5), .A1 (nx3605), .B0 (
                      des_acc_5), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix500 (.Y (nx499), .A0 (nx3591), .A1 (nx3586), .B0 (
                          nx68), .C0 (acc_5)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_5 (.Q (acc_5), .CK (wb_clk_i), .D (nx422), .R (
                       wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix3542 (.Y (nx3592), .A0 (nx3584), .A1 (nx3598), .B0 (
                       nx3612), .C0 (nx3613)) ;
    AOI22_X0P5M_A12TS ix3544 (.Y (nx3612), .A0 (des2_4), .A1 (nx3605), .B0 (
                      des_acc_4), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix3545 (.Y (nx3613), .A0 (nx3584), .A1 (nx3586), .B0 (
                          nx68), .C0 (acc_4)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_4 (.Q (acc_4), .CK (wb_clk_i), .D (nx3592), 
                       .R (wb_rst_i)) ;
    XNOR3_X0P5M_A12TS ix3546 (.Y (nx3614), .A (nx3594), .B (nx3595), .C (nx3596)
                      ) ;
    XOR2_X0P5M_A12TS ix3547 (.Y (nx3594), .A (nx3593), .B (nx425)) ;
    OAI211_X0P5M_A12TS ix3548 (.Y (nx3593), .A0 (nx3587), .A1 (nx3615), .B0 (
                       nx3617), .C0 (nx3618)) ;
    NAND3_X0P5A_A12TS ix3550 (.Y (nx3615), .A (nx3616), .B (desCy), .C (nx68)) ;
    OAI21_X0P5M_A12TS ix3551 (.Y (nx3616), .A0 (nx3607), .A1 (wr_addr_2), .B0 (
                      nx3586)) ;
    AOI22_X0P5M_A12TS ix3552 (.Y (nx3617), .A0 (des2_3), .A1 (nx3605), .B0 (
                      des_acc_3), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix3553 (.Y (nx3618), .A0 (nx3587), .A1 (nx3586), .B0 (
                          nx3588), .C0 (acc_3)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_3 (.Q (acc_3), .CK (wb_clk_i), .D (nx3593), 
                       .R (wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix3554 (.Y (nx425), .A0 (nx3589), .A1 (nx3615), .B0 (
                       nx523), .C0 (nx525)) ;
    AOI22_X0P5M_A12TS ix524 (.Y (nx523), .A0 (des2_2), .A1 (nx3605), .B0 (
                      des_acc_2), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix526 (.Y (nx525), .A0 (nx3589), .A1 (nx3586), .B0 (
                          nx3588), .C0 (acc_2)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_2 (.Q (acc_2), .CK (wb_clk_i), .D (nx425), .R (
                       wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix3555 (.Y (nx3595), .A0 (nx3591), .A1 (nx3615), .B0 (
                       nx3619), .C0 (nx3620)) ;
    AOI22_X0P5M_A12TS ix3556 (.Y (nx3619), .A0 (des2_1), .A1 (nx3605), .B0 (
                      des_acc_1), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix3557 (.Y (nx3620), .A0 (nx3591), .A1 (nx3586), .B0 (
                          nx3588), .C0 (acc_1)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_1 (.Q (acc_1), .CK (wb_clk_i), .D (nx3595), 
                       .R (wb_rst_i)) ;
    OAI211_X0P5M_A12TS ix315 (.Y (nx3596), .A0 (nx3584), .A1 (nx3615), .B0 (
                       nx3621), .C0 (nx3622)) ;
    AOI22_X0P5M_A12TS ix3558 (.Y (nx3621), .A0 (des2_0), .A1 (nx3605), .B0 (
                      des_acc_0), .B1 (nx100)) ;
    AO21A1AI2_X0P5M_A12TS ix3560 (.Y (nx3622), .A0 (nx3584), .A1 (nx3586), .B0 (
                          nx3588), .C0 (acc_0)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_0 (.Q (acc_0), .CK (wb_clk_i), .D (nx3596), 
                       .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix3561 (.Y (nx3588), .A (nx3616)) ;
    INV_X0P5B_A12TS ix69 (.Y (nx68), .A (nx3606)) ;
    INV_X0P5B_A12TS ix3562 (.Y (nx3584), .A (nx3604)) ;
    NAND4B_X0P5M_A12TS ix3563 (.Y (nx3599), .AN (wr_addr_4), .B (wr_addr_5), .C (
                       wr_addr_6), .D (wr_addr_7)) ;
    NAND4B_X0P5M_A12TS ix3564 (.Y (nx3603), .AN (wr_bit_r_dup_1790), .B (nx3601)
                       , .C (we), .D (nx3604)) ;
    NOR2B_X0P7M_A12TS ix3566 (.Y (nx3605), .AN (wr_sfr_1), .B (wr_sfr_0)) ;
    NAND2B_X0P7M_A12TS ix3567 (.Y (nx3589), .AN (wr_addr_0), .B (wr_addr_1)) ;
    NAND2B_X0P7M_A12TS ix3568 (.Y (nx3591), .AN (wr_addr_1), .B (wr_addr_0)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_0__dup_70485 (.Q (b_reg_0), .CK (wb_clk_i), 
                       .D (nx3683), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3623 (.Y (nx3683), .A (nx534), .B (nx3691), .S0 (nx3692)
                      ) ;
    AOI21_X0P5M_A12TS ix535 (.Y (nx534), .A0 (des_acc_0), .A1 (nx3690), .B0 (
                      nx3676)) ;
    INV_X0P5B_A12TS ix3624 (.Y (nx3690), .A (wr_bit_r_dup_1790)) ;
    AND2_X0P5M_A12TS ix3626 (.Y (nx3676), .A (wr_bit_r_dup_1790), .B (desCy)) ;
    INV_X0P5B_A12TS ix3627 (.Y (nx3691), .A (b_reg_0)) ;
    INV_X0P5B_A12TS ix3628 (.Y (nx3693), .A (wr_addr_0)) ;
    INV_X0P5B_A12TS ix3629 (.Y (nx3695), .A (wr_addr_2)) ;
    NAND3_X0P5A_A12TS ix3630 (.Y (nx3696), .A (wr_addr_6), .B (wr_addr_4), .C (
                      wr_addr_5)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_1__dup_70494 (.Q (b_reg_1), .CK (wb_clk_i), 
                       .D (nx3684), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3632 (.Y (nx3684), .A (nx3697), .B (nx3698), .S0 (nx3699
                      )) ;
    AOI21_X0P5M_A12TS ix3633 (.Y (nx3697), .A0 (des_acc_1), .A1 (nx3690), .B0 (
                      nx3676)) ;
    INV_X0P5B_A12TS ix3634 (.Y (nx3698), .A (b_reg_1)) ;
    AOI31_X0P5M_A12TS ix3635 (.Y (nx3699), .A0 (nx3677), .A1 (wr_addr_0), .A2 (
                      nx3695), .B0 (nx38)) ;
    NOR3_X0P5A_A12TS ix3636 (.Y (nx3677), .A (nx3701), .B (wr_addr_1), .C (
                     nx3690)) ;
    NAND4B_X0P5M_A12TS ix3638 (.Y (nx3701), .AN (wr_addr_3), .B (nx3675), .C (we
                       ), .D (wr_addr_7)) ;
    NOR2_X0P5A_A12TS ix3639 (.Y (nx38), .A (wr_bit_r_dup_1790), .B (nx3692)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_2__dup_70502 (.Q (b_reg_2), .CK (wb_clk_i), 
                       .D (nx3685), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3640 (.Y (nx3685), .A (nx569), .B (nx571), .S0 (nx3680)
                      ) ;
    INV_X0P5B_A12TS ix570 (.Y (nx569), .A (b_reg_2)) ;
    AOI21_X0P5M_A12TS ix572 (.Y (nx571), .A0 (des_acc_2), .A1 (nx3690), .B0 (
                      nx3676)) ;
    OAI31_X0P5M_A12TS ix3641 (.Y (nx3680), .A0 (nx574), .A1 (wr_addr_0), .A2 (
                      wr_addr_2), .B0 (nx3702)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_3__dup_70507 (.Q (b_reg_3), .CK (wb_clk_i), 
                       .D (nx3686), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3642 (.Y (nx3686), .A (nx3703), .B (nx3704), .S0 (nx3681
                      )) ;
    INV_X0P5B_A12TS ix3644 (.Y (nx3703), .A (b_reg_3)) ;
    AOI21_X0P5M_A12TS ix3645 (.Y (nx3704), .A0 (des_acc_3), .A1 (nx3690), .B0 (
                      nx3676)) ;
    OAI31_X0P5M_A12TS ix3646 (.Y (nx3681), .A0 (nx574), .A1 (nx3693), .A2 (
                      wr_addr_2), .B0 (nx3702)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_4__dup_70512 (.Q (b_reg_4), .CK (wb_clk_i), 
                       .D (nx3687), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3647 (.Y (nx3687), .A (nx3705), .B (nx3706), .S0 (nx592)
                      ) ;
    AOI21_X0P5M_A12TS ix3648 (.Y (nx3705), .A0 (des_acc_4), .A1 (nx3690), .B0 (
                      nx3676)) ;
    INV_X0P5B_A12TS ix3650 (.Y (nx3706), .A (b_reg_4)) ;
    AOI31_X0P5M_A12TS ix593 (.Y (nx592), .A0 (nx3677), .A1 (nx3693), .A2 (
                      wr_addr_2), .B0 (nx38)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_5__dup_70517 (.Q (b_reg_5), .CK (wb_clk_i), 
                       .D (nx3689), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3651 (.Y (nx3689), .A (nx3707), .B (nx3708), .S0 (nx600)
                      ) ;
    AOI21_X0P5M_A12TS ix3652 (.Y (nx3707), .A0 (des_acc_5), .A1 (nx3690), .B0 (
                      nx3676)) ;
    INV_X0P5B_A12TS ix3653 (.Y (nx3708), .A (b_reg_5)) ;
    AOI31_X0P5M_A12TS ix601 (.Y (nx600), .A0 (nx3677), .A1 (wr_addr_0), .A2 (
                      wr_addr_2), .B0 (nx38)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_6__dup_70522 (.Q (b_reg_6), .CK (wb_clk_i), 
                       .D (nx512), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3654 (.Y (nx512), .A (nx604), .B (nx606), .S0 (nx3682)
                      ) ;
    INV_X0P5B_A12TS ix605 (.Y (nx604), .A (b_reg_6)) ;
    AOI21_X0P5M_A12TS ix3655 (.Y (nx606), .A0 (des_acc_6), .A1 (nx3690), .B0 (
                      nx3676)) ;
    OAI31_X0P5M_A12TS ix3656 (.Y (nx3682), .A0 (nx574), .A1 (wr_addr_0), .A2 (
                      nx3695), .B0 (nx3702)) ;
    DFFRPQ_X0P5M_A12TS reg_data_out_7__dup_70527 (.Q (b_reg_7), .CK (wb_clk_i), 
                       .D (nx522), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix3658 (.Y (nx522), .A (nx3709), .B (nx3710), .S0 (nx615)
                      ) ;
    AOI21_X0P5M_A12TS ix3659 (.Y (nx3709), .A0 (nx3690), .A1 (des_acc_7), .B0 (
                      nx3676)) ;
    INV_X0P5B_A12TS ix3660 (.Y (nx3710), .A (b_reg_7)) ;
    AOI31_X0P5M_A12TS ix616 (.Y (nx615), .A0 (nx3679), .A1 (wr_addr_0), .A2 (
                      wr_addr_2), .B0 (nx38)) ;
    INV_X0P5B_A12TS ix3661 (.Y (nx3679), .A (nx574)) ;
    INV_X0P5B_A12TS ix3662 (.Y (nx3702), .A (nx38)) ;
    INV_X0P5B_A12TS ix3663 (.Y (nx3675), .A (nx3696)) ;
    OR4_X0P5M_A12TS ix3664 (.Y (nx3692), .A (wr_addr_1), .B (wr_addr_0), .C (
                    wr_addr_2), .D (nx3701)) ;
    NAND3B_X0P5M_A12TS ix575 (.Y (nx574), .AN (nx3701), .B (wr_addr_1), .C (
                       wr_bit_r_dup_1790)) ;
    AOI21_X0P5M_A12TS ix3711 (.Y (sp_w_0), .A0 (nx3803), .A1 (nx323), .B0 (
                      nx3819)) ;
    NAND3B_X0P5M_A12TS ix3712 (.Y (nx3803), .AN (ram_wr_sel_2), .B (ram_wr_sel_1
                       ), .C (ram_wr_sel_0)) ;
    INV_X0P5B_A12TS ix324 (.Y (nx323), .A (sp_0__dup_3810)) ;
    SDFFSQ_X0P5M_A12TS reg_sp_0 (.Q (sp_0__dup_3810), .CK (wb_clk_i), .D (des1_0
                       ), .SE (NOT_nx30), .SI (sp_0), .SN (nx359)) ;
    NAND4XXXB_X1M_A12TS ix328 (.Y (NOT_nx30), .DN (wr_bit_r_dup_1790), .A (
                        nx3800), .B (nx3801), .C (we)) ;
    NOR3_X0P5A_A12TS ix3713 (.Y (nx3800), .A (nx331), .B (wr_addr_5), .C (
                     wr_addr_4)) ;
    NAND3B_X0P5M_A12TS ix332 (.Y (nx331), .AN (wr_addr_6), .B (wr_addr_0), .C (
                       wr_addr_7)) ;
    NOR3_X0P5A_A12TS ix3714 (.Y (nx3801), .A (wr_addr_1), .B (wr_addr_3), .C (
                     wr_addr_2)) ;
    OAI21_X0P5M_A12TS ix3715 (.Y (sp_0), .A0 (nx30), .A1 (nx345), .B0 (nx357)) ;
    XOR2_X0P5M_A12TS ix346 (.Y (nx345), .A (nx3812), .B (nx3825)) ;
    NAND2_X0P5A_A12TS ix3716 (.Y (nx3812), .A (nx3803), .B (pop)) ;
    DFFRPQ_X0P5M_A12TS reg_pop (.Q (pop), .CK (wb_clk_i), .D (nx3811), .R (
                       wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix3717 (.Y (nx3811), .A (ram_rd_sel_2), .B (nx3824)) ;
    NAND2_X0P5A_A12TS ix3718 (.Y (nx3824), .A (ram_rd_sel_0), .B (ram_rd_sel_1)
                      ) ;
    XOR2_X0P5M_A12TS ix3719 (.Y (nx3825), .A (nx3803), .B (nx355)) ;
    MXIT2_X0P5M_A12TS ix356 (.Y (nx355), .A (des1_0), .B (sp_0__dup_3810), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix358 (.Y (nx357), .A (nx30), .B (des1_0)) ;
    INV_X0P5B_A12TS ix3720 (.Y (nx359), .A (wb_rst_i)) ;
    AOI21_X0P5M_A12TS ix3722 (.Y (sp_w_1), .A0 (nx3826), .A1 (nx3829), .B0 (
                      nx3820)) ;
    NAND2_X0P5A_A12TS ix3724 (.Y (nx3826), .A (sp_0__dup_3810), .B (nx3827)) ;
    INV_X0P5B_A12TS ix3725 (.Y (nx3829), .A (sp_1__dup_3809)) ;
    SDFFSQ_X0P5M_A12TS reg_sp_1 (.Q (sp_1__dup_3809), .CK (wb_clk_i), .D (des1_1
                       ), .SE (NOT_nx30), .SI (sp_1), .SN (nx359)) ;
    OAI21_X0P5M_A12TS ix3726 (.Y (sp_1), .A0 (nx30), .A1 (nx377), .B0 (nx385)) ;
    XOR2_X0P5M_A12TS ix378 (.Y (nx377), .A (nx3813), .B (nx381)) ;
    OAI21_X0P5M_A12TS ix3727 (.Y (nx3813), .A0 (nx3827), .A1 (pop), .B0 (nx355)
                      ) ;
    XOR2_X0P5M_A12TS ix382 (.Y (nx381), .A (nx3803), .B (nx3830)) ;
    MXIT2_X0P5M_A12TS ix3728 (.Y (nx3830), .A (des1_1), .B (sp_1__dup_3809), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix386 (.Y (nx385), .A (nx30), .B (des1_1)) ;
    AOI21_X0P5M_A12TS ix3729 (.Y (sp_w_2), .A0 (nx3831), .A1 (nx393), .B0 (
                      nx3821)) ;
    NAND3_X0P5A_A12TS ix3730 (.Y (nx3831), .A (sp_1__dup_3809), .B (
                      sp_0__dup_3810), .C (nx3827)) ;
    INV_X0P5B_A12TS ix394 (.Y (nx393), .A (sp_2__dup_3808)) ;
    SDFFSQ_X0P5M_A12TS reg_sp_2 (.Q (sp_2__dup_3808), .CK (wb_clk_i), .D (des1_2
                       ), .SE (NOT_nx30), .SI (sp_2), .SN (nx359)) ;
    OAI21_X0P5M_A12TS ix3731 (.Y (sp_2), .A0 (nx30), .A1 (nx399), .B0 (nx3833)
                      ) ;
    XNOR2_X0P5M_A12TS ix400 (.Y (nx399), .A (nx3832), .B (nx405)) ;
    CGENI_X1M_A12TS ix3732 (.CON (nx3832), .A (nx3813), .B (nx3803), .CI (nx303)
                    ) ;
    XOR2_X0P5M_A12TS ix406 (.Y (nx405), .A (nx3803), .B (nx407)) ;
    MXIT2_X0P5M_A12TS ix408 (.Y (nx407), .A (des1_2), .B (sp_2__dup_3808), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix3734 (.Y (nx3833), .A (nx30), .B (des1_2)) ;
    NOR2_X0P5A_A12TS ix3736 (.Y (nx3821), .A (nx393), .B (nx3831)) ;
    SDFFRPQ_X0P5M_A12TS reg_sp_3 (.Q (sp_3__dup_3807), .CK (wb_clk_i), .D (
                        des1_3), .R (wb_rst_i), .SE (NOT_nx30), .SI (sp_3)) ;
    OAI21_X0P5M_A12TS ix187 (.Y (sp_3), .A0 (nx30), .A1 (nx3834), .B0 (nx431)) ;
    XOR2_X0P5M_A12TS ix3737 (.Y (nx3834), .A (nx3814), .B (nx3835)) ;
    CGENI_X1M_A12TS ix3738 (.CON (nx3814), .A (nx3832), .B (nx3827), .CI (nx407)
                    ) ;
    XOR2_X0P5M_A12TS ix3739 (.Y (nx3835), .A (nx3803), .B (nx429)) ;
    MXIT2_X0P5M_A12TS ix430 (.Y (nx429), .A (des1_3), .B (sp_3__dup_3807), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix432 (.Y (nx431), .A (nx30), .B (des1_3)) ;
    AOI21_X0P5M_A12TS ix3740 (.Y (sp_w_4), .A0 (nx3836), .A1 (nx3837), .B0 (
                      nx3823)) ;
    NAND2_X0P5A_A12TS ix3742 (.Y (nx3836), .A (sp_3__dup_3807), .B (nx3821)) ;
    INV_X0P5B_A12TS ix3743 (.Y (nx3837), .A (sp_4__dup_3806)) ;
    SDFFRPQ_X0P5M_A12TS reg_sp_4 (.Q (sp_4__dup_3806), .CK (wb_clk_i), .D (
                        des1_4), .R (wb_rst_i), .SE (NOT_nx30), .SI (sp_4)) ;
    OAI21_X0P5M_A12TS ix3744 (.Y (sp_4), .A0 (nx30), .A1 (nx441), .B0 (nx3842)
                      ) ;
    XNOR2_X0P5M_A12TS ix442 (.Y (nx441), .A (nx3839), .B (nx3841)) ;
    CGENI_X1M_A12TS ix3745 (.CON (nx3839), .A (nx3814), .B (nx3803), .CI (nx305)
                    ) ;
    XOR2_X0P5M_A12TS ix3746 (.Y (nx3841), .A (nx3803), .B (nx448)) ;
    MXIT2_X0P5M_A12TS ix449 (.Y (nx448), .A (des1_4), .B (sp_4__dup_3806), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix3747 (.Y (nx3842), .A (nx30), .B (des1_4)) ;
    NOR2_X0P5A_A12TS ix3748 (.Y (nx3823), .A (nx3837), .B (nx3836)) ;
    SDFFRPQ_X0P5M_A12TS reg_sp_5 (.Q (sp_5__dup_3805), .CK (wb_clk_i), .D (
                        des1_5), .R (wb_rst_i), .SE (NOT_nx30), .SI (sp_5)) ;
    OAI21_X0P5M_A12TS ix3749 (.Y (sp_5), .A0 (nx30), .A1 (nx3843), .B0 (nx3845)
                      ) ;
    XOR2_X0P5M_A12TS ix3750 (.Y (nx3843), .A (nx3815), .B (nx3844)) ;
    CGENI_X1M_A12TS ix3751 (.CON (nx3815), .A (nx3839), .B (nx3827), .CI (nx448)
                    ) ;
    XOR2_X0P5M_A12TS ix3752 (.Y (nx3844), .A (nx3803), .B (nx465)) ;
    MXIT2_X0P5M_A12TS ix466 (.Y (nx465), .A (des1_5), .B (sp_5__dup_3805), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix3753 (.Y (nx3845), .A (nx30), .B (des1_5)) ;
    AOI21_X0P5M_A12TS ix3754 (.Y (sp_w_6), .A0 (nx3846), .A1 (nx473), .B0 (nx382
                      )) ;
    NAND2_X0P5A_A12TS ix3755 (.Y (nx3846), .A (sp_5__dup_3805), .B (nx3823)) ;
    INV_X0P5B_A12TS ix474 (.Y (nx473), .A (sp_6__dup_3804)) ;
    SDFFRPQ_X0P5M_A12TS reg_sp_6 (.Q (sp_6__dup_3804), .CK (wb_clk_i), .D (
                        des1_6), .R (wb_rst_i), .SE (NOT_nx30), .SI (sp_6)) ;
    OAI21_X0P5M_A12TS ix3756 (.Y (sp_6), .A0 (nx30), .A1 (nx3847), .B0 (nx486)
                      ) ;
    XNOR2_X0P5M_A12TS ix3758 (.Y (nx3847), .A (nx479), .B (nx3849)) ;
    CGENI_X1M_A12TS ix480 (.CON (nx479), .A (nx3815), .B (nx3803), .CI (nx309)
                    ) ;
    XOR2_X0P5M_A12TS ix3760 (.Y (nx3849), .A (nx3850), .B (nx3803)) ;
    MXIT2_X0P5M_A12TS ix3761 (.Y (nx3850), .A (des1_6), .B (sp_6__dup_3804), .S0 (
                      NOT_nx30)) ;
    NAND2_X0P5A_A12TS ix3762 (.Y (nx486), .A (nx30), .B (des1_6)) ;
    NOR2_X0P5A_A12TS ix383 (.Y (nx382), .A (nx473), .B (nx3846)) ;
    XOR2_X0P5M_A12TS ix385 (.Y (sp_w_7), .A (sp_7__dup_3799), .B (nx382)) ;
    SDFFRPQ_X0P5M_A12TS reg_sp_7 (.Q (sp_7__dup_3799), .CK (wb_clk_i), .D (
                        des1_7), .R (wb_rst_i), .SE (NOT_nx30), .SI (sp_7)) ;
    MXT2_X0P5M_A12TS ix3763 (.Y (sp_7), .A (des1_7), .B (nx3818), .S0 (NOT_nx30)
                     ) ;
    XNOR3_X0P5M_A12TS ix3764 (.Y (nx3818), .A (nx3817), .B (nx3803), .C (nx3851)
                      ) ;
    CGENI_X1M_A12TS ix3765 (.CON (nx3817), .A (nx479), .B (nx3850), .CI (nx3827)
                    ) ;
    MXIT2_X0P5M_A12TS ix3766 (.Y (nx3851), .A (des1_7), .B (sp_7__dup_3799), .S0 (
                      NOT_nx30)) ;
    INV_X0P5B_A12TS ix3768 (.Y (nx3820), .A (nx3831)) ;
    INV_X0P5B_A12TS ix3769 (.Y (nx3819), .A (nx3826)) ;
    INV_X0P5B_A12TS ix287 (.Y (nx309), .A (nx465)) ;
    INV_X0P5B_A12TS ix3770 (.Y (nx305), .A (nx429)) ;
    INV_X0P5B_A12TS ix3771 (.Y (nx303), .A (nx3830)) ;
    INV_X0P5B_A12TS ix3772 (.Y (nx3827), .A (nx3803)) ;
    INV_X0P5B_A12TS ix3773 (.Y (nx30), .A (NOT_nx30)) ;
    OA21_X0P5M_A12TS ix3774 (.Y (sp_w_3), .A0 (nx3821), .A1 (sp_3__dup_3807), .B0 (
                     nx3836)) ;
    OA21_X0P5M_A12TS ix3775 (.Y (sp_w_5), .A0 (nx3823), .A1 (sp_5__dup_3805), .B0 (
                     nx3846)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_0 (.Q (dptr_lo_0), .CK (wb_clk_i), .D (
                        des_acc_0), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_0)) ;
    AND2_X0P5M_A12TS ix651 (.Y (NOT_nx158), .A (nx652), .B (nx3880)) ;
    NAND4_X0P5A_A12TS ix653 (.Y (nx652), .A (nx3885), .B (nx659), .C (we), .D (
                      nx3898)) ;
    NOR3_X0P5A_A12TS ix3852 (.Y (nx3885), .A (nx655), .B (wr_addr_2), .C (
                     wr_bit_r_dup_1790)) ;
    NAND2_X0P5A_A12TS ix656 (.Y (nx655), .A (wr_addr_1), .B (nx657)) ;
    INV_X0P5B_A12TS ix658 (.Y (nx657), .A (wr_addr_3)) ;
    AOI31_X0P5M_A12TS ix660 (.Y (nx659), .A0 (nx3881), .A1 (nx3898), .A2 (nx3884
                      ), .B0 (nx670)) ;
    AND4_X0P5M_A12TS ix3853 (.Y (nx3881), .A (wr_addr_1), .B (nx657), .C (nx3896
                     ), .D (wr_addr_0)) ;
    INV_X0P5B_A12TS ix3854 (.Y (nx3896), .A (wr_addr_2)) ;
    NOR3_X0P5A_A12TS ix3856 (.Y (nx3898), .A (wr_addr_4), .B (wr_addr_5), .C (
                     nx3883)) ;
    NAND2B_X0P7M_A12TS ix3857 (.Y (nx3883), .AN (wr_addr_6), .B (wr_addr_7)) ;
    NAND2_X0P5A_A12TS ix3858 (.Y (nx3880), .A (wr_sfr_1), .B (wr_sfr_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_1 (.Q (dptr_lo_1), .CK (wb_clk_i), .D (
                        des_acc_1), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_2 (.Q (dptr_lo_2), .CK (wb_clk_i), .D (
                        des_acc_2), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_3 (.Q (dptr_lo_3), .CK (wb_clk_i), .D (
                        des_acc_3), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_4 (.Q (dptr_lo_4), .CK (wb_clk_i), .D (
                        des_acc_4), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_5 (.Q (dptr_lo_5), .CK (wb_clk_i), .D (
                        des_acc_5), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_6 (.Q (dptr_lo_6), .CK (wb_clk_i), .D (
                        des_acc_6), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_data_lo_7 (.Q (dptr_lo_7), .CK (wb_clk_i), .D (
                        des_acc_7), .R (wb_rst_i), .SE (NOT_nx158), .SI (
                        dptr_lo_7)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_0 (.Q (dptr_hi_0), .CK (wb_clk_i), .D (nx3888
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3859 (.Y (nx3888), .A0 (nx3899), .A1 (nx659), .B0 (
                      nx3900)) ;
    AOI32_X0P5M_A12TS ix3860 (.Y (nx3899), .A0 (des2_0), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_0), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix3861 (.Y (nx3900), .A (dptr_hi_0), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_1 (.Q (dptr_hi_1), .CK (wb_clk_i), .D (nx3889
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3862 (.Y (nx3889), .A0 (nx3901), .A1 (nx659), .B0 (nx690
                      )) ;
    AOI32_X0P5M_A12TS ix3863 (.Y (nx3901), .A0 (des2_1), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_1), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix691 (.Y (nx690), .A (dptr_hi_1), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_2 (.Q (dptr_hi_2), .CK (wb_clk_i), .D (nx3890
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3864 (.Y (nx3890), .A0 (nx3902), .A1 (nx659), .B0 (
                      nx3903)) ;
    AOI32_X0P5M_A12TS ix3865 (.Y (nx3902), .A0 (des2_2), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_2), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix3866 (.Y (nx3903), .A (dptr_hi_2), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_3 (.Q (dptr_hi_3), .CK (wb_clk_i), .D (nx3891
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3867 (.Y (nx3891), .A0 (nx700), .A1 (nx659), .B0 (nx702)
                      ) ;
    AOI32_X0P5M_A12TS ix701 (.Y (nx700), .A0 (des2_3), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_3), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix703 (.Y (nx702), .A (dptr_hi_3), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_4 (.Q (dptr_hi_4), .CK (wb_clk_i), .D (nx3892
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3868 (.Y (nx3892), .A0 (nx706), .A1 (nx659), .B0 (nx708)
                      ) ;
    AOI32_X0P5M_A12TS ix707 (.Y (nx706), .A0 (des2_4), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_4), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix709 (.Y (nx708), .A (dptr_hi_4), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_5 (.Q (dptr_hi_5), .CK (wb_clk_i), .D (nx3893
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3869 (.Y (nx3893), .A0 (nx712), .A1 (nx659), .B0 (nx3905
                      )) ;
    AOI32_X0P5M_A12TS ix3870 (.Y (nx712), .A0 (des2_5), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_5), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix3871 (.Y (nx3905), .A (dptr_hi_5), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_6 (.Q (dptr_hi_6), .CK (wb_clk_i), .D (nx549)
                       , .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix550 (.Y (nx549), .A0 (nx718), .A1 (nx659), .B0 (nx720)
                      ) ;
    AOI32_X0P5M_A12TS ix719 (.Y (nx718), .A0 (des2_6), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_6), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix3872 (.Y (nx720), .A (dptr_hi_6), .B (nx659)) ;
    DFFRPQ_X0P5M_A12TS reg_data_hi_7 (.Q (dptr_hi_7), .CK (wb_clk_i), .D (nx3895
                       ), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix3874 (.Y (nx3895), .A0 (nx724), .A1 (nx659), .B0 (nx3906
                      )) ;
    AOI32_X0P5M_A12TS ix725 (.Y (nx724), .A0 (des2_7), .A1 (wr_sfr_1), .A2 (
                      wr_sfr_0), .B0 (des_acc_7), .B1 (nx3880)) ;
    NAND2_X0P5A_A12TS ix3875 (.Y (nx3906), .A (dptr_hi_7), .B (nx659)) ;
    INV_X0P5B_A12TS ix671 (.Y (nx670), .A (nx3880)) ;
    NOR2B_X0P7M_A12TS ix3876 (.Y (nx3884), .AN (we), .B (wr_bit_r_dup_1790)) ;
    MXT2_X0P5M_A12TS ix3907 (.Y (bank_sel_0), .A (des1_3), .B (psw_3), .S0 (
                     nx3996)) ;
    DFFRPQ_X0P5M_A12TS reg_data_3 (.Q (psw_3), .CK (wb_clk_i), .D (nx3994), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3908 (.Y (nx3994), .A (psw_3), .B (nx3988), .S0 (nx3986)
                     ) ;
    OAI21_X0P5M_A12TS ix3910 (.Y (nx3988), .A0 (nx478), .A1 (nx3996), .B0 (
                      nx3997)) ;
    INV_X0P5B_A12TS ix479 (.Y (nx478), .A (des1_3)) ;
    NOR3_X0P5A_A12TS ix3911 (.Y (nx3973), .A (nx483), .B (wr_addr_5), .C (
                     wr_addr_3)) ;
    NAND3_X0P5A_A12TS ix484 (.Y (nx483), .A (wr_addr_7), .B (wr_addr_4), .C (
                      wr_addr_6)) ;
    NOR3_X0P5A_A12TS ix3912 (.Y (nx3974), .A (wr_addr_0), .B (wr_addr_2), .C (
                     wr_addr_1)) ;
    NAND2_X0P5A_A12TS ix3914 (.Y (nx3997), .A (desCy), .B (nx3996)) ;
    NAND2_X0P5A_A12TS ix3915 (.Y (nx3986), .A (nx3998), .B (nx505)) ;
    NAND4_X0P5A_A12TS ix3916 (.Y (nx3998), .A (nx493), .B (wr_addr_1), .C (
                      wr_addr_0), .D (nx3999)) ;
    INV_X0P5B_A12TS ix494 (.Y (nx493), .A (wr_addr_2)) ;
    NAND2_X0P5A_A12TS ix3917 (.Y (nx3999), .A (nx4000), .B (nx3996)) ;
    NAND4B_X0P5M_A12TS ix3918 (.Y (nx4000), .AN (nx4001), .B (we), .C (nx4002), 
                       .D (wr_bit_r_dup_1790)) ;
    INV_X0P5B_A12TS ix3919 (.Y (nx4002), .A (wr_addr_3)) ;
    NAND2_X0P5A_A12TS ix506 (.Y (nx505), .A (nx4000), .B (nx3999)) ;
    MXT2_X0P5M_A12TS ix3920 (.Y (bank_sel_1), .A (des1_4), .B (psw_4), .S0 (
                     nx3996)) ;
    DFFRPQ_X0P5M_A12TS reg_data_4 (.Q (psw_4), .CK (wb_clk_i), .D (nx3995), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3921 (.Y (nx3995), .A (nx3989), .B (psw_4), .S0 (nx4003)
                     ) ;
    OAI21_X0P5M_A12TS ix3922 (.Y (nx3989), .A0 (nx511), .A1 (nx3996), .B0 (
                      nx3997)) ;
    INV_X0P5B_A12TS ix512 (.Y (nx511), .A (des1_4)) ;
    AOI31_X0P5M_A12TS ix3923 (.Y (nx4003), .A0 (nx3979), .A1 (wr_addr_2), .A2 (
                      nx521), .B0 (nx3978)) ;
    NOR2_X0P5A_A12TS ix3924 (.Y (nx3979), .A (wr_addr_1), .B (nx3977)) ;
    INV_X0P5B_A12TS ix522 (.Y (nx521), .A (wr_addr_0)) ;
    DFFRPQ_X0P5M_A12TS reg_data_1 (.Q (psw_1), .CK (wb_clk_i), .D (nx404), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3926 (.Y (nx404), .A (nx3980), .B (psw_1), .S0 (nx4004)
                     ) ;
    AOI31_X0P5M_A12TS ix3927 (.Y (nx4004), .A0 (nx3979), .A1 (nx493), .A2 (
                      wr_addr_0), .B0 (nx3978)) ;
    DFFRPQ_X0P5M_A12TS reg_data_2 (.Q (psw_2), .CK (wb_clk_i), .D (nx3990), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3928 (.Y (nx3990), .A (psw_2), .B (nx3982), .S0 (nx3981)
                     ) ;
    NAND2_X0P5A_A12TS ix3929 (.Y (nx3982), .A (nx4005), .B (nx4006)) ;
    AOI22_X0P5M_A12TS ix3930 (.Y (nx4005), .A0 (des1_2), .A1 (nx3975), .B0 (
                      desOv), .B1 (nx3977)) ;
    NAND2_X0P5A_A12TS ix3932 (.Y (nx4006), .A (desCy), .B (nx3972)) ;
    AO21A1AI2_X0P5M_A12TS ix3933 (.Y (nx3981), .A0 (nx3996), .A1 (nx4008), .B0 (
                          nx3972), .C0 (nx4009)) ;
    INV_X0P5B_A12TS ix3934 (.Y (nx4008), .A (psw_set_1)) ;
    NAND4_X0P5A_A12TS ix3935 (.Y (nx4009), .A (nx493), .B (wr_addr_1), .C (nx521
                      ), .D (nx3972)) ;
    DFFRPQ_X0P5M_A12TS reg_data_5 (.Q (psw_5), .CK (wb_clk_i), .D (nx3991), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3936 (.Y (nx3991), .A (nx3983), .B (psw_5), .S0 (nx4011)
                     ) ;
    AOI31_X0P5M_A12TS ix3937 (.Y (nx4011), .A0 (nx3979), .A1 (wr_addr_2), .A2 (
                      wr_addr_0), .B0 (nx3978)) ;
    DFFRPQ_X0P5M_A12TS reg_data_6 (.Q (srcAc), .CK (wb_clk_i), .D (nx3992), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3938 (.Y (nx3992), .A (srcAc), .B (nx3985), .S0 (nx3984)
                     ) ;
    NAND2_X0P5A_A12TS ix3940 (.Y (nx3985), .A (nx4012), .B (nx4006)) ;
    AOI22_X0P5M_A12TS ix3941 (.Y (nx4012), .A0 (des1_6), .A1 (nx3975), .B0 (
                      desAc), .B1 (nx3977)) ;
    OAI211_X0P5M_A12TS ix3942 (.Y (nx3984), .A0 (nx4013), .A1 (nx4014), .B0 (
                       nx4015), .C0 (nx505)) ;
    NAND2_X0P5A_A12TS ix3943 (.Y (nx4013), .A (wr_addr_2), .B (wr_addr_1)) ;
    AO21A1AI2_X0P5M_A12TS ix3944 (.Y (nx4014), .A0 (psw_set_0), .A1 (psw_set_1)
                          , .B0 (nx3999), .C0 (nx521)) ;
    NAND3_X0P5A_A12TS ix3946 (.Y (nx4015), .A (nx4000), .B (psw_set_0), .C (
                      psw_set_1)) ;
    DFFRPQ_X0P5M_A12TS reg_data_7 (.Q (cy), .CK (wb_clk_i), .D (nx3993), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3947 (.Y (nx3993), .A (nx180), .B (cy), .S0 (nx4018)) ;
    NAND2_X0P5A_A12TS ix3948 (.Y (nx180), .A (nx4016), .B (nx4006)) ;
    AOI22_X0P5M_A12TS ix3949 (.Y (nx4016), .A0 (des1_7), .A1 (nx3975), .B0 (
                      desCy), .B1 (nx3977)) ;
    AOI31_X0P5M_A12TS ix3950 (.Y (nx4018), .A0 (wr_addr_0), .A1 (wr_addr_2), .A2 (
                      wr_addr_1), .B0 (nx4000)) ;
    INV_X0P5B_A12TS ix3951 (.Y (nx3978), .A (nx505)) ;
    INV_X0P5B_A12TS ix3952 (.Y (nx3977), .A (nx3999)) ;
    INV_X0P5B_A12TS ix3953 (.Y (nx3975), .A (nx3996)) ;
    INV_X0P5B_A12TS ix3954 (.Y (nx3972), .A (nx4000)) ;
    NAND4B_X0P5M_A12TS ix3955 (.Y (nx3996), .AN (wr_bit_r_dup_1790), .B (nx3973)
                       , .C (nx3974), .D (we)) ;
    NAND4B_X0P5M_A12TS ix3956 (.Y (nx4001), .AN (wr_addr_5), .B (wr_addr_4), .C (
                       wr_addr_6), .D (wr_addr_7)) ;
    OAI2XB1_X0P5M_A12TS ix3958 (.Y (nx3980), .A0 (nx3996), .A1N (des1_1), .B0 (
                        nx3997)) ;
    OAI2XB1_X0P5M_A12TS ix3960 (.Y (nx3983), .A0 (nx3996), .A1N (des1_5), .B0 (
                        nx3997)) ;
    MXT2_X0P5M_A12TS ix4019 (.Y (p3_data_0), .A (p3_i[0]), .B (p3_o[0]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_0 (.Q (p3_o[0]), .CK (wb_clk_i), .D (nx4237), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4020 (.Y (nx4237), .A (nx4208), .B (p3_o[0]), .S0 (nx4270
                     )) ;
    NAND2_X0P5A_A12TS ix1908 (.Y (nx4269), .A (wr_bit_r_dup_1790), .B (desCy)) ;
    NAND2_X0P5A_A12TS ix4021 (.Y (nx4270), .A (nx4272), .B (nx4206)) ;
    OAI31_X0P5M_A12TS ix4022 (.Y (nx4206), .A0 (nx4274), .A1 (wr_addr_1), .A2 (
                      wr_addr_0), .B0 (nx4277)) ;
    INV_X1M_A12TS ix4024 (.Y (nx4279), .A (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4026 (.Y (p3_data_1), .A (p3_i[1]), .B (p3_o[1]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_1 (.Q (p3_o[1]), .CK (wb_clk_i), .D (nx4238), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4027 (.Y (nx4238), .A (p3_o[1]), .B (nx4211), .S0 (nx4209
                     )) ;
    NOR2_X0P5A_A12TS ix4028 (.Y (nx4209), .A (nx4203), .B (nx1934)) ;
    NAND2_X0P5A_A12TS ix4029 (.Y (nx4203), .A (wr_addr_5), .B (wr_addr_4)) ;
    AOI31_X0P5M_A12TS ix4030 (.Y (nx1934), .A0 (nx16), .A1 (nx4280), .A2 (
                      wr_addr_0), .B0 (nx4205)) ;
    INV_X0P5B_A12TS ix4031 (.Y (nx4280), .A (wr_addr_1)) ;
    MXT2_X0P5M_A12TS ix4032 (.Y (p3_data_2), .A (p3_i[2]), .B (p3_o[2]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_2 (.Q (p3_o[2]), .CK (wb_clk_i), .D (nx4239), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4034 (.Y (nx4239), .A (p3_o[2]), .B (nx4213), .S0 (nx92)
                     ) ;
    NOR2_X0P5A_A12TS ix4035 (.Y (nx92), .A (nx4203), .B (nx4282)) ;
    AOI31_X0P5M_A12TS ix4036 (.Y (nx4282), .A0 (nx16), .A1 (wr_addr_1), .A2 (
                      nx1949), .B0 (nx4205)) ;
    INV_X0P5B_A12TS ix4039 (.Y (nx1949), .A (wr_addr_0)) ;
    MXT2_X0P5M_A12TS ix4040 (.Y (p3_data_3), .A (p3_i[3]), .B (p3_o[3]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_3 (.Q (p3_o[3]), .CK (wb_clk_i), .D (nx4241), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4041 (.Y (nx4241), .A (p3_o[3]), .B (nx4217), .S0 (nx4215
                     )) ;
    NOR2_X0P5A_A12TS ix4042 (.Y (nx4215), .A (nx4203), .B (nx1956)) ;
    AOI31_X0P5M_A12TS ix4043 (.Y (nx1956), .A0 (nx16), .A1 (wr_addr_1), .A2 (
                      wr_addr_0), .B0 (nx4205)) ;
    MXT2_X0P5M_A12TS ix4044 (.Y (p3_data_4), .A (p3_i[4]), .B (p3_o[4]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_4 (.Q (p3_o[4]), .CK (wb_clk_i), .D (nx4242), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4045 (.Y (nx4242), .A (nx4219), .B (p3_o[4]), .S0 (nx1962
                     )) ;
    NAND2_X0P5A_A12TS ix4046 (.Y (nx1962), .A (nx4272), .B (nx4218)) ;
    OAI31_X0P5M_A12TS ix4047 (.Y (nx4218), .A0 (nx4284), .A1 (wr_addr_1), .A2 (
                      wr_addr_0), .B0 (nx4277)) ;
    NAND2_X0P5A_A12TS ix4050 (.Y (nx4284), .A (wr_addr_2), .B (we)) ;
    MXT2_X0P5M_A12TS ix4052 (.Y (p3_data_5), .A (p3_i[5]), .B (p3_o[5]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_5 (.Q (p3_o[5]), .CK (wb_clk_i), .D (nx4243), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4053 (.Y (nx4243), .A (nx4222), .B (p3_o[5]), .S0 (nx1971
                     )) ;
    NAND2_X0P5A_A12TS ix4054 (.Y (nx1971), .A (nx4272), .B (nx4220)) ;
    OAI31_X0P5M_A12TS ix4055 (.Y (nx4220), .A0 (nx4284), .A1 (wr_addr_1), .A2 (
                      nx1949), .B0 (nx4277)) ;
    MXT2_X0P5M_A12TS ix229 (.Y (p3_data_6), .A (p3_i[6]), .B (p3_o[6]), .S0 (rmw
                     )) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_6 (.Q (p3_o[6]), .CK (wb_clk_i), .D (nx4244), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4056 (.Y (nx4244), .A (nx220), .B (p3_o[6]), .S0 (nx4286)
                     ) ;
    NAND2_X0P5A_A12TS ix4057 (.Y (nx4286), .A (nx4272), .B (nx4223)) ;
    OAI31_X0P5M_A12TS ix4059 (.Y (nx4223), .A0 (nx4284), .A1 (nx4280), .A2 (
                      wr_addr_0), .B0 (nx4277)) ;
    MXT2_X0P5M_A12TS ix4060 (.Y (p3_data_7), .A (p3_i[7]), .B (p3_o[7]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p3_out_7 (.Q (p3_o[7]), .CK (wb_clk_i), .D (nx4245), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4062 (.Y (nx4245), .A (nx248), .B (p3_o[7]), .S0 (nx4287)
                     ) ;
    NAND2_X0P5A_A12TS ix4063 (.Y (nx4287), .A (nx4272), .B (nx4224)) ;
    OAI31_X0P5M_A12TS ix4064 (.Y (nx4224), .A0 (nx4284), .A1 (nx4280), .A2 (
                      nx1949), .B0 (nx4277)) ;
    MXT2_X0P5M_A12TS ix4065 (.Y (p2_data_0), .A (p2_i[0]), .B (p2_o[0]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_0 (.Q (p2_o[0]), .CK (wb_clk_i), .D (nx4247), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4066 (.Y (nx4247), .A (nx4208), .B (p2_o[0]), .S0 (nx4289
                     )) ;
    NAND2_X0P5A_A12TS ix4067 (.Y (nx4289), .A (nx1993), .B (nx4206)) ;
    MXT2_X0P5M_A12TS ix4068 (.Y (p2_data_1), .A (p2_i[1]), .B (p2_o[1]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_1 (.Q (p2_o[1]), .CK (wb_clk_i), .D (nx1673), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4069 (.Y (nx1673), .A (p2_o[1]), .B (nx4211), .S0 (nx4227
                     )) ;
    NOR2_X0P5A_A12TS ix4070 (.Y (nx4227), .A (nx4225), .B (nx1934)) ;
    MXT2_X0P5M_A12TS ix4071 (.Y (p2_data_2), .A (p2_i[2]), .B (p2_o[2]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_2 (.Q (p2_o[2]), .CK (wb_clk_i), .D (nx1683), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4072 (.Y (nx1683), .A (p2_o[2]), .B (nx4213), .S0 (nx4228
                     )) ;
    NOR2_X0P5A_A12TS ix4074 (.Y (nx4228), .A (nx4225), .B (nx4282)) ;
    MXT2_X0P5M_A12TS ix4075 (.Y (p2_data_3), .A (p2_i[3]), .B (p2_o[3]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_3 (.Q (p2_o[3]), .CK (wb_clk_i), .D (nx4248), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4076 (.Y (nx4248), .A (p2_o[3]), .B (nx4217), .S0 (nx4229
                     )) ;
    NOR2_X0P5A_A12TS ix4077 (.Y (nx4229), .A (nx4225), .B (nx1956)) ;
    MXT2_X0P5M_A12TS ix341 (.Y (p2_data_4), .A (p2_i[4]), .B (p2_o[4]), .S0 (rmw
                     )) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_4 (.Q (p2_o[4]), .CK (wb_clk_i), .D (nx1703), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4079 (.Y (nx1703), .A (nx4219), .B (p2_o[4]), .S0 (nx4290
                     )) ;
    NAND2_X0P5A_A12TS ix4080 (.Y (nx4290), .A (nx1993), .B (nx4218)) ;
    MXT2_X0P5M_A12TS ix4081 (.Y (p2_data_5), .A (p2_i[5]), .B (p2_o[5]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_5 (.Q (p2_o[5]), .CK (wb_clk_i), .D (nx1713), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix1714 (.Y (nx1713), .A (nx4222), .B (p2_o[5]), .S0 (nx4291
                     )) ;
    NAND2_X0P5A_A12TS ix4082 (.Y (nx4291), .A (nx1993), .B (nx4220)) ;
    MXT2_X0P5M_A12TS ix4083 (.Y (p2_data_6), .A (p2_i[6]), .B (p2_o[6]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_6 (.Q (p2_o[6]), .CK (wb_clk_i), .D (nx1723), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix1724 (.Y (nx1723), .A (nx220), .B (p2_o[6]), .S0 (nx4292)
                     ) ;
    NAND2_X0P5A_A12TS ix4084 (.Y (nx4292), .A (nx1993), .B (nx4223)) ;
    MXT2_X0P5M_A12TS ix4086 (.Y (p2_data_7), .A (p2_i[7]), .B (p2_o[7]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p2_out_7 (.Q (p2_o[7]), .CK (wb_clk_i), .D (nx4249), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4087 (.Y (nx4249), .A (nx248), .B (p2_o[7]), .S0 (nx4293)
                     ) ;
    NAND2_X0P5A_A12TS ix4088 (.Y (nx4293), .A (nx1993), .B (nx4224)) ;
    MXT2_X0P5M_A12TS ix4089 (.Y (p1_data_0), .A (p1_i[0]), .B (p1_o[0]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_0 (.Q (p1_o[0]), .CK (wb_clk_i), .D (nx4250), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4090 (.Y (nx4250), .A (nx4208), .B (p1_o[0]), .S0 (nx4295
                     )) ;
    NAND2_X0P5A_A12TS ix4092 (.Y (nx4295), .A (nx4296), .B (nx4206)) ;
    MXT2_X0P5M_A12TS ix4093 (.Y (p1_data_1), .A (p1_i[1]), .B (p1_o[1]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_1 (.Q (p1_o[1]), .CK (wb_clk_i), .D (nx1753), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix1754 (.Y (nx1753), .A (p1_o[1]), .B (nx4211), .S0 (nx4232
                     )) ;
    NOR2_X0P5A_A12TS ix4094 (.Y (nx4232), .A (nx4231), .B (nx1934)) ;
    MXT2_X0P5M_A12TS ix4095 (.Y (p1_data_2), .A (p1_i[2]), .B (p1_o[2]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_2 (.Q (p1_o[2]), .CK (wb_clk_i), .D (nx4251), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4096 (.Y (nx4251), .A (p1_o[2]), .B (nx4213), .S0 (nx432)
                     ) ;
    NOR2_X0P5A_A12TS ix4099 (.Y (nx432), .A (nx4231), .B (nx4282)) ;
    MXT2_X0P5M_A12TS ix4100 (.Y (p1_data_3), .A (p1_i[3]), .B (p1_o[3]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_3 (.Q (p1_o[3]), .CK (wb_clk_i), .D (nx4252), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4101 (.Y (nx4252), .A (p1_o[3]), .B (nx4217), .S0 (nx4233
                     )) ;
    NOR2_X0P5A_A12TS ix4102 (.Y (nx4233), .A (nx4231), .B (nx1956)) ;
    MXT2_X0P5M_A12TS ix4103 (.Y (p1_data_4), .A (p1_i[4]), .B (p1_o[4]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_4 (.Q (p1_o[4]), .CK (wb_clk_i), .D (nx4253), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4104 (.Y (nx4253), .A (nx4219), .B (p1_o[4]), .S0 (nx4298
                     )) ;
    NAND2_X0P5A_A12TS ix4106 (.Y (nx4298), .A (nx4296), .B (nx4218)) ;
    MXT2_X0P5M_A12TS ix4107 (.Y (p1_data_5), .A (p1_i[5]), .B (p1_o[5]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_5 (.Q (p1_o[5]), .CK (wb_clk_i), .D (nx4254), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4108 (.Y (nx4254), .A (nx4222), .B (p1_o[5]), .S0 (nx4300
                     )) ;
    NAND2_X0P5A_A12TS ix4110 (.Y (nx4300), .A (nx4296), .B (nx4220)) ;
    MXT2_X0P5M_A12TS ix4111 (.Y (p1_data_6), .A (p1_i[6]), .B (p1_o[6]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_6 (.Q (p1_o[6]), .CK (wb_clk_i), .D (nx4256), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4112 (.Y (nx4256), .A (nx220), .B (p1_o[6]), .S0 (nx4301)
                     ) ;
    NAND2_X0P5A_A12TS ix4113 (.Y (nx4301), .A (nx4296), .B (nx4223)) ;
    MXT2_X0P5M_A12TS ix4114 (.Y (p1_data_7), .A (p1_i[7]), .B (p1_o[7]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p1_out_7 (.Q (p1_o[7]), .CK (wb_clk_i), .D (nx4258), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4115 (.Y (nx4258), .A (nx248), .B (p1_o[7]), .S0 (nx4303)
                     ) ;
    NAND2_X0P5A_A12TS ix4116 (.Y (nx4303), .A (nx4296), .B (nx4224)) ;
    MXT2_X0P5M_A12TS ix539 (.Y (p0_data_0), .A (p0_i[0]), .B (p0_o[0]), .S0 (rmw
                     )) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_0 (.Q (p0_o[0]), .CK (wb_clk_i), .D (nx4260), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4119 (.Y (nx4260), .A (nx4208), .B (p0_o[0]), .S0 (nx4304
                     )) ;
    NAND2_X0P5A_A12TS ix4120 (.Y (nx4304), .A (nx4305), .B (nx4206)) ;
    NOR2_X0P5A_A12TS ix4122 (.Y (nx4305), .A (wr_addr_5), .B (wr_addr_4)) ;
    MXT2_X0P5M_A12TS ix4123 (.Y (p0_data_1), .A (p0_i[1]), .B (p0_o[1]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_1 (.Q (p0_o[1]), .CK (wb_clk_i), .D (nx4261), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4124 (.Y (nx4261), .A (p0_o[1]), .B (nx4211), .S0 (nx4235
                     )) ;
    NOR2_X0P5A_A12TS ix4125 (.Y (nx4235), .A (nx4234), .B (nx1934)) ;
    MXT2_X0P5M_A12TS ix4126 (.Y (p0_data_2), .A (p0_i[2]), .B (p0_o[2]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_2 (.Q (p0_o[2]), .CK (wb_clk_i), .D (nx4262), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix1844 (.Y (nx4262), .A (p0_o[2]), .B (nx4213), .S0 (nx562)
                     ) ;
    NOR2_X0P5A_A12TS ix4127 (.Y (nx562), .A (nx4234), .B (nx4282)) ;
    MXT2_X0P5M_A12TS ix4129 (.Y (p0_data_3), .A (p0_i[3]), .B (p0_o[3]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_3 (.Q (p0_o[3]), .CK (wb_clk_i), .D (nx4263), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4130 (.Y (nx4263), .A (p0_o[3]), .B (nx4217), .S0 (nx4236
                     )) ;
    NOR2_X0P5A_A12TS ix4131 (.Y (nx4236), .A (nx4234), .B (nx1956)) ;
    MXT2_X0P5M_A12TS ix603 (.Y (p0_data_4), .A (p0_i[4]), .B (p0_o[4]), .S0 (rmw
                     )) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_4 (.Q (p0_o[4]), .CK (wb_clk_i), .D (nx4264), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4132 (.Y (nx4264), .A (nx4219), .B (p0_o[4]), .S0 (nx4307
                     )) ;
    NAND2_X0P5A_A12TS ix4133 (.Y (nx4307), .A (nx4305), .B (nx4218)) ;
    MXT2_X0P5M_A12TS ix4134 (.Y (p0_data_5), .A (p0_i[5]), .B (p0_o[5]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_5 (.Q (p0_o[5]), .CK (wb_clk_i), .D (nx4265), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4136 (.Y (nx4265), .A (nx4222), .B (p0_o[5]), .S0 (nx4309
                     )) ;
    NAND2_X0P5A_A12TS ix2097 (.Y (nx4309), .A (nx4305), .B (nx4220)) ;
    MXT2_X0P5M_A12TS ix4137 (.Y (p0_data_6), .A (p0_i[6]), .B (p0_o[6]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_6 (.Q (p0_o[6]), .CK (wb_clk_i), .D (nx4266), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix4139 (.Y (nx4266), .A (nx220), .B (p0_o[6]), .S0 (nx4311)
                     ) ;
    NAND2_X0P5A_A12TS ix4140 (.Y (nx4311), .A (nx4305), .B (nx4223)) ;
    MXT2_X0P5M_A12TS ix4141 (.Y (p0_data_7), .A (p0_i[7]), .B (p0_o[7]), .S0 (
                     rmw)) ;
    DFFSQ_X0P5M_A12TS reg_p0_out_7 (.Q (p0_o[7]), .CK (wb_clk_i), .D (nx4268), .SN (
                      nx4279)) ;
    MXT2_X0P5M_A12TS ix1894 (.Y (nx4268), .A (nx248), .B (p0_o[7]), .S0 (nx4312)
                     ) ;
    NAND2_X0P5A_A12TS ix2107 (.Y (nx4312), .A (nx4305), .B (nx4224)) ;
    INV_X0P5B_A12TS ix4142 (.Y (nx4234), .A (nx4305)) ;
    INV_X0P5B_A12TS ix4143 (.Y (nx4231), .A (nx4296)) ;
    INV_X0P5B_A12TS ix4144 (.Y (nx4225), .A (nx1993)) ;
    INV_X0P5B_A12TS ix4145 (.Y (nx4274), .A (nx16)) ;
    INV_X0P5B_A12TS ix4146 (.Y (nx4205), .A (nx4277)) ;
    INV_X0P5B_A12TS ix4147 (.Y (nx4272), .A (nx4203)) ;
    OAI2XB1_X0P5M_A12TS ix4149 (.Y (nx4208), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_0), .B0 (nx4269)) ;
    OAI2XB1_X0P5M_A12TS ix4150 (.Y (nx4211), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_1), .B0 (nx4269)) ;
    NOR2B_X0P7M_A12TS ix4151 (.Y (nx16), .AN (we), .B (wr_addr_2)) ;
    OAI2XB1_X0P5M_A12TS ix4152 (.Y (nx4213), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_2), .B0 (nx4269)) ;
    OAI2XB1_X0P5M_A12TS ix4153 (.Y (nx4217), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_3), .B0 (nx4269)) ;
    OAI2XB1_X0P5M_A12TS ix4154 (.Y (nx4219), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_4), .B0 (nx4269)) ;
    OAI2XB1_X0P5M_A12TS ix4155 (.Y (nx4222), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_5), .B0 (nx4269)) ;
    OAI2XB1_X0P5M_A12TS ix4156 (.Y (nx220), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_6), .B0 (nx4269)) ;
    OAI2XB1_X0P5M_A12TS ix4159 (.Y (nx248), .A0 (wr_bit_r_dup_1790), .A1N (
                        des1_7), .B0 (nx4269)) ;
    NOR2B_X0P7M_A12TS ix4160 (.Y (nx1993), .AN (wr_addr_5), .B (wr_addr_4)) ;
    NOR2B_X0P7M_A12TS ix4161 (.Y (nx4296), .AN (wr_addr_4), .B (wr_addr_5)) ;
    NAND2B_X0P7M_A12TS ix4162 (.Y (nx4277), .AN (wr_bit_r_dup_1790), .B (we)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_0 (.Q (sbuf_0), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_3), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_0)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_3 (.Q (sbuf_rxd_tmp_3), .CK (wb_clk_i), 
                       .D (nx4730), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4313 (.Y (nx4730), .A0 (nx4690), .A1 (nx4816), .B0 (
                          nx4799), .C0 (nx4839)) ;
    OAI21_X0P5M_A12TS ix4314 (.Y (nx4690), .A0 (nx2994), .A1 (nx3102), .B0 (
                      nx4793)) ;
    INV_X0P5B_A12TS ix4315 (.Y (nx2994), .A (rx_done)) ;
    DFFSQ_X0P5M_A12TS reg_rx_done (.Q (rx_done), .CK (wb_clk_i), .D (nx2800), .SN (
                      nx3094)) ;
    MXIT2_X0P5M_A12TS ix4316 (.Y (nx2800), .A (nx2994), .B (nx2998), .S0 (nx4669
                      )) ;
    NOR2_X0P5A_A12TS ix4317 (.Y (nx2998), .A (nx3000), .B (sbuf_rxd_tmp_0)) ;
    NOR2_X0P5A_A12TS ix4319 (.Y (nx3003), .A (scon_6), .B (scon_7)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_6 (.Q (scon_6), .CK (wb_clk_i), .D (nx4697), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4320 (.Y (nx4697), .A (nx4634), .B (scon_6), .S0 (nx4740)
                     ) ;
    OAI21_X0P5M_A12TS ix4322 (.Y (nx4634), .A0 (nx3008), .A1 (nx4735), .B0 (
                      nx3024)) ;
    INV_X0P5B_A12TS ix4324 (.Y (nx3008), .A (des1_6)) ;
    NAND4_X0P5A_A12TS ix4325 (.Y (nx4735), .A (nx3012), .B (nx3014), .C (nx4622)
                      , .D (nx4624)) ;
    INV_X0P5B_A12TS ix4327 (.Y (nx3012), .A (wr_addr_2)) ;
    INV_X0P5B_A12TS ix4328 (.Y (nx3014), .A (wr_bit_r_dup_1790)) ;
    NAND4B_X0P5M_A12TS ix4330 (.Y (nx4739), .AN (wr_addr_6), .B (wr_addr_7), .C (
                       nx3019), .D (we)) ;
    INV_X0P5B_A12TS ix4331 (.Y (nx3019), .A (wr_addr_5)) ;
    NOR2_X0P5A_A12TS ix4332 (.Y (nx4624), .A (wr_addr_1), .B (wr_addr_0)) ;
    NAND2_X0P5A_A12TS ix4334 (.Y (nx3024), .A (desCy), .B (nx4623)) ;
    NOR2_X0P5A_A12TS ix4336 (.Y (nx4623), .A (nx3014), .B (nx3027)) ;
    AOI31_X0P5M_A12TS ix4337 (.Y (nx4740), .A0 (nx4631), .A1 (wr_addr_1), .A2 (
                      nx3040), .B0 (nx4627)) ;
    NOR2_X0P5A_A12TS ix4338 (.Y (nx4631), .A (nx3012), .B (nx3037)) ;
    NOR2_X0P5A_A12TS ix4340 (.Y (nx3037), .A (nx4625), .B (nx4623)) ;
    INV_X0P5B_A12TS ix4342 (.Y (nx3040), .A (wr_addr_0)) ;
    NOR2_X0P5A_A12TS ix4343 (.Y (nx4627), .A (nx4623), .B (nx3037)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_7 (.Q (scon_7), .CK (wb_clk_i), .D (nx4695), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4344 (.Y (nx4695), .A (nx4632), .B (scon_7), .S0 (nx3048)
                     ) ;
    OAI21_X0P5M_A12TS ix4346 (.Y (nx4632), .A0 (nx3046), .A1 (nx4735), .B0 (
                      nx3024)) ;
    INV_X0P5B_A12TS ix4348 (.Y (nx3046), .A (des1_7)) ;
    AOI31_X0P5M_A12TS ix4350 (.Y (nx3048), .A0 (wr_addr_0), .A1 (wr_addr_1), .A2 (
                      nx4631), .B0 (nx4627)) ;
    DFFRPQ_X0P5M_A12TS reg_receive (.Q (receive), .CK (wb_clk_i), .D (nx2680), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4352 (.Y (nx2680), .A (nx3052), .B (nx4742), .S0 (nx4687
                      )) ;
    INV_X0P5B_A12TS ix4353 (.Y (nx3052), .A (receive)) ;
    AOI31_X0P5M_A12TS ix4354 (.Y (nx4742), .A0 (nx644), .A1 (nx3085), .A2 (rxd_r
                      ), .B0 (nx4636)) ;
    AOI211_X0P5M_A12TS ix4356 (.Y (nx3057), .A0 (receive), .A1 (shift_re), .B0 (
                       nx3003), .C0 (nx2994)) ;
    DFFRPQ_X0P5M_A12TS reg_shift_re (.Q (shift_re), .CK (wb_clk_i), .D (nx4676)
                       , .R (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix4358 (.Y (nx4676), .A (nx3061), .B (nx3069)) ;
    AOI221_X0P5M_A12TS ix4359 (.Y (nx3061), .A0 (scon_7), .A1 (nx3063), .B0 (
                       rclk), .B1 (brate2), .C0 (nx4672)) ;
    INV_X0P5B_A12TS ix4360 (.Y (nx3063), .A (scon_6)) ;
    NOR3_X0P5A_A12TS ix4363 (.Y (nx4672), .A (t1_ow_buf), .B (rclk), .C (nx3067)
                     ) ;
    DFFRPQ_X0P5M_A12TS reg_t1_ow_buf (.Q (t1_ow_buf), .CK (wb_clk_i), .D (tf1), 
                       .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix4364 (.Y (nx3067), .A (tf1)) ;
    NOR2_X0P5A_A12TS ix4366 (.Y (nx3069), .A (smod_clk_re), .B (pcon_7)) ;
    DFFRPQ_X0P5M_A12TS reg_smod_clk_re (.Q (smod_clk_re), .CK (wb_clk_i), .D (
                       nx4717), .R (wb_rst_i)) ;
    XOR2_X0P5M_A12TS ix4367 (.Y (nx4717), .A (smod_clk_re), .B (nx4674)) ;
    NOR2_X0P5A_A12TS ix4368 (.Y (nx4674), .A (pcon_7), .B (nx3061)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_7 (.Q (pcon_7), .CK (wb_clk_i), .D (des1_7), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_7)) ;
    OR6_X0P5M_A12TS ix4370 (.Y (NOT_nx444), .A (wr_addr_3), .B (nx3012), .C (
                    wr_addr_4), .D (nx4739), .E (wr_bit_r_dup_1790), .F (nx4629)
                    ) ;
    NAND2_X0P5A_A12TS ix4371 (.Y (nx4629), .A (wr_addr_0), .B (wr_addr_1)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_4 (.Q (scon_4), .CK (wb_clk_i), .D (nx4698), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4372 (.Y (nx4698), .A (nx4638), .B (scon_4), .S0 (nx3083)
                     ) ;
    OAI21_X0P5M_A12TS ix4374 (.Y (nx4638), .A0 (nx3081), .A1 (nx4735), .B0 (
                      nx3024)) ;
    INV_X0P5B_A12TS ix4375 (.Y (nx3081), .A (des1_4)) ;
    AOI21_X0P5M_A12TS ix4376 (.Y (nx3083), .A0 (nx4631), .A1 (nx4624), .B0 (
                      nx4627)) ;
    INV_X0P5B_A12TS ix4377 (.Y (nx3085), .A (rxd_i)) ;
    DFFSQ_X0P5M_A12TS reg_rxd_r (.Q (rxd_r), .CK (wb_clk_i), .D (nx4722), .SN (
                      nx3094)) ;
    MXT2_X0P5M_A12TS ix4379 (.Y (nx4722), .A (rxd_r), .B (rxd_i), .S0 (nx4689)
                     ) ;
    AOI21_X0P5M_A12TS ix4380 (.Y (nx4689), .A0 (scon_4), .A1 (nx3090), .B0 (
                      nx4677)) ;
    INV_X0P5B_A12TS ix4382 (.Y (nx3090), .A (shift_re)) ;
    INV_X0P5B_A12TS ix4384 (.Y (nx3094), .A (wb_rst_i)) ;
    AOI31_X0P5M_A12TS ix4385 (.Y (nx4687), .A0 (nx3098), .A1 (rx_done), .A2 (
                      nx4744), .B0 (nx4671)) ;
    NAND3_X0P5A_A12TS ix4386 (.Y (nx3098), .A (nx3057), .B (scon_4), .C (
                      shift_re)) ;
    NAND3_X0P5A_A12TS ix4388 (.Y (nx4744), .A (nx3102), .B (rx_done), .C (nx3003
                      )) ;
    NAND3_X0P5A_A12TS ix4390 (.Y (nx3102), .A (nx3003), .B (pres_ow), .C (
                      receive)) ;
    AOI31_X0P5M_A12TS ix775 (.Y (nx4671), .A0 (nx3105), .A1 (scon_4), .A2 (
                      nx3052), .B0 (nx4744)) ;
    INV_X0P5B_A12TS ix4392 (.Y (nx3105), .A (scon_0)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_0 (.Q (scon_0), .CK (wb_clk_i), .D (nx2660), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4393 (.Y (nx2660), .A (nx4686), .B (scon_0), .S0 (nx4776)
                     ) ;
    OAI211_X0P5M_A12TS ix4394 (.Y (nx4686), .A0 (nx3110), .A1 (nx4735), .B0 (
                       nx3112), .C0 (nx3024)) ;
    INV_X0P5B_A12TS ix4395 (.Y (nx3110), .A (des1_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tx_done (.Q (tx_done), .CK (wb_clk_i), .D (nx2560), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4398 (.Y (nx2560), .A (tx_done), .B (nx344), .S0 (nx4640)
                     ) ;
    OAI21_X0P5M_A12TS ix4400 (.Y (nx344), .A0 (nx3119), .A1 (nx4659), .B0 (
                      nx4775)) ;
    NAND4_X1M_A12TS ix4402 (.Y (nx3121), .A (nx3012), .B (nx3014), .C (nx3123), 
                    .D (nx4622)) ;
    NOR2_X0P5A_A12TS ix4404 (.Y (nx3123), .A (nx3040), .B (wr_addr_1)) ;
    DFFRPQ_X0P5M_A12TS reg_trans (.Q (trans), .CK (wb_clk_i), .D (nx4713), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4406 (.Y (nx4713), .A (nx3121), .B (nx3127), .S0 (nx3129
                      )) ;
    INV_X0P5B_A12TS ix4407 (.Y (nx3127), .A (trans)) ;
    NAND3_X0P5A_A12TS ix4408 (.Y (nx3129), .A (nx4640), .B (nx3132), .C (nx4660)
                      ) ;
    AOI32_X0P5M_A12TS ix549 (.Y (nx4640), .A0 (nx3132), .A1 (nx4746), .A2 (
                      nx3136), .B0 (nx3149), .B1 (nx4643)) ;
    NAND4_X0P5A_A12TS ix4410 (.Y (nx4746), .A (pres_ow), .B (trans), .C (nx3003)
                      , .D (nx3121)) ;
    DFFRPQ_X0P5M_A12TS reg_shift_tr (.Q (shift_tr), .CK (wb_clk_i), .D (nx4663)
                       , .R (wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix4411 (.Y (nx4663), .A (nx3140), .B (nx3143)) ;
    AOI221_X0P5M_A12TS ix4412 (.Y (nx3140), .A0 (scon_7), .A1 (nx3063), .B0 (
                       tclk), .B1 (brate2), .C0 (nx418)) ;
    NOR3_X0P5A_A12TS ix4413 (.Y (nx418), .A (t1_ow_buf), .B (tclk), .C (nx3067)
                     ) ;
    NOR2_X0P5A_A12TS ix4418 (.Y (nx3143), .A (smod_clk_tr), .B (pcon_7)) ;
    DFFRPQ_X0P5M_A12TS reg_smod_clk_tr (.Q (smod_clk_tr), .CK (wb_clk_i), .D (
                       nx4715), .R (wb_rst_i)) ;
    XOR2_X0P5M_A12TS ix4419 (.Y (nx4715), .A (smod_clk_tr), .B (nx4661)) ;
    NOR2_X0P5A_A12TS ix4420 (.Y (nx4661), .A (pcon_7), .B (nx3140)) ;
    INV_X0P5B_A12TS ix4422 (.Y (nx3151), .A (tr_count_3)) ;
    DFFRPQ_X0P5M_A12TS reg_tr_count_3 (.Q (tr_count_3), .CK (wb_clk_i), .D (
                       nx4716), .R (wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix4424 (.Y (nx4716), .A0 (nx3151), .A1 (nx4665), .B0 (
                      nx4748)) ;
    NAND2_X0P5A_A12TS ix4426 (.Y (nx4665), .A (nx4747), .B (nx3121)) ;
    NAND3_X0P5A_A12TS ix4427 (.Y (nx4747), .A (nx4635), .B (trans), .C (shift_tr
                      )) ;
    NAND3_X0P5A_A12TS ix4428 (.Y (nx4748), .A (nx3121), .B (nx4666), .C (nx4665)
                      ) ;
    XNOR2_X0P5M_A12TS ix4429 (.Y (nx4666), .A (tr_count_3), .B (nx3161)) ;
    NAND3_X0P5A_A12TS ix4431 (.Y (nx3161), .A (tr_count_2), .B (tr_count_1), .C (
                      tr_count_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tr_count_2 (.Q (tr_count_2), .CK (wb_clk_i), .D (
                       nx2540), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4432 (.Y (nx2540), .A (nx3165), .B (nx3167), .S0 (nx4665
                      )) ;
    INV_X0P5B_A12TS ix4434 (.Y (nx3165), .A (tr_count_2)) ;
    OAI211_X0P5M_A12TS ix4436 (.Y (nx3167), .A0 (nx2326), .A1 (tr_count_2), .B0 (
                       nx3121), .C0 (nx3161)) ;
    INV_X0P5B_A12TS ix4438 (.Y (nx3170), .A (tr_count_1)) ;
    DFFRPQ_X0P5M_A12TS reg_tr_count_1 (.Q (tr_count_1), .CK (wb_clk_i), .D (
                       nx2530), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4439 (.Y (nx2530), .A (nx3170), .B (nx3174), .S0 (nx4665
                      )) ;
    OAI211_X0P5M_A12TS ix4442 (.Y (nx3174), .A0 (tr_count_0), .A1 (tr_count_1), 
                       .B0 (nx3121), .C0 (nx3180)) ;
    DFFRPQ_X0P5M_A12TS reg_tr_count_0 (.Q (tr_count_0), .CK (wb_clk_i), .D (
                       nx2520), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4443 (.Y (nx2520), .A0 (tr_count_0), .A1 (nx4639), .A2 (
                      nx3136), .B0 (nx3178)) ;
    NAND2_X0P5A_A12TS ix4444 (.Y (nx3178), .A (tr_count_0), .B (nx3136)) ;
    NAND2_X0P5A_A12TS ix4446 (.Y (nx3180), .A (tr_count_1), .B (tr_count_0)) ;
    NOR2_X0P5A_A12TS ix4448 (.Y (nx4643), .A (nx4639), .B (nx4747)) ;
    AOI22_X0P5M_A12TS ix4450 (.Y (nx4660), .A0 (nx4659), .A1 (nx4643), .B0 (
                      nx4775), .B1 (nx4648)) ;
    NAND4_X0P5A_A12TS ix4451 (.Y (nx4659), .A (nx3187), .B (nx4767), .C (nx4769)
                      , .D (nx4772)) ;
    NOR2_X0P5A_A12TS ix3188 (.Y (nx3187), .A (nx4658), .B (nx4656)) ;
    INV_X0P5B_A12TS ix4453 (.Y (nx3190), .A (sbuf_txd_3)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_3 (.Q (sbuf_txd_3), .CK (wb_clk_i), .D (
                       nx4709), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4454 (.Y (nx4709), .A (nx3190), .B (nx3194), .S0 (nx4645
                      )) ;
    AOI222_X0P5M_A12TS ix3195 (.Y (nx3194), .A0 (sbuf_txd_4), .A1 (nx3121), .B0 (
                       des1_3), .B1 (nx4647), .C0 (des1_2), .C1 (nx4646)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_4 (.Q (sbuf_txd_4), .CK (wb_clk_i), .D (
                       nx4708), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4456 (.Y (nx4708), .A (nx3198), .B (nx4750), .S0 (nx4645
                      )) ;
    INV_X0P5B_A12TS ix3199 (.Y (nx3198), .A (sbuf_txd_4)) ;
    AOI222_X0P5M_A12TS ix4458 (.Y (nx4750), .A0 (sbuf_txd_5), .A1 (nx3121), .B0 (
                       des1_4), .B1 (nx4647), .C0 (des1_3), .C1 (nx4646)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_5 (.Q (sbuf_txd_5), .CK (wb_clk_i), .D (
                       nx4706), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4459 (.Y (nx4706), .A (nx4751), .B (nx4752), .S0 (nx4645
                      )) ;
    INV_X0P5B_A12TS ix3205 (.Y (nx4751), .A (sbuf_txd_5)) ;
    AOI222_X0P5M_A12TS ix4460 (.Y (nx4752), .A0 (sbuf_txd_6), .A1 (nx3121), .B0 (
                       des1_5), .B1 (nx4647), .C0 (des1_4), .C1 (nx4646)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_6 (.Q (sbuf_txd_6), .CK (wb_clk_i), .D (
                       nx4705), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4462 (.Y (nx4705), .A (nx4753), .B (nx4754), .S0 (nx4645
                      )) ;
    INV_X0P5B_A12TS ix3211 (.Y (nx4753), .A (sbuf_txd_6)) ;
    AOI222_X0P5M_A12TS ix3213 (.Y (nx4754), .A0 (sbuf_txd_7), .A1 (nx3121), .B0 (
                       des1_6), .B1 (nx4647), .C0 (des1_5), .C1 (nx4646)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_7 (.Q (sbuf_txd_7), .CK (wb_clk_i), .D (
                       nx4703), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4463 (.Y (nx4703), .A (nx4756), .B (nx4757), .S0 (nx4645
                      )) ;
    INV_X0P5B_A12TS ix3217 (.Y (nx4756), .A (sbuf_txd_7)) ;
    AOI222_X0P5M_A12TS ix3219 (.Y (nx4757), .A0 (sbuf_txd_8), .A1 (nx3121), .B0 (
                       des1_7), .B1 (nx4647), .C0 (des1_6), .C1 (nx4646)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_txd_8 (.Q (sbuf_txd_8), .CK (wb_clk_i), .D (
                        nx4655), .R (wb_rst_i), .SE (NOT_nx2324), .SI (
                        sbuf_txd_8)) ;
    OAI211_X0P5M_A12TS ix4464 (.Y (nx4655), .A0 (nx3046), .A1 (nx3121), .B0 (
                       nx4758), .C0 (nx4765)) ;
    NAND2_X0P5A_A12TS ix4466 (.Y (nx4758), .A (sbuf_txd_9), .B (nx3121)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_txd_9 (.Q (sbuf_txd_9), .CK (wb_clk_i), .D (
                        nx4654), .R (wb_rst_i), .SE (NOT_nx2324), .SI (
                        sbuf_txd_9)) ;
    INV_X0P5B_A12TS ix4468 (.Y (nx4759), .A (sbuf_txd_10)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_10 (.Q (sbuf_txd_10), .CK (wb_clk_i), .D (
                       nx4701), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4470 (.Y (nx4701), .A (nx4759), .B (nx4760), .S0 (nx4645
                      )) ;
    NAND2_X0P5A_A12TS ix3231 (.Y (nx4760), .A (scon_7), .B (nx4639)) ;
    NOR3_X0P5A_A12TS ix4471 (.Y (nx4645), .A (nx4641), .B (nx344), .C (nx4762)
                     ) ;
    NOR2_X0P5A_A12TS ix4474 (.Y (nx4641), .A (trans), .B (nx4639)) ;
    AO21A1AI2_X0P5M_A12TS ix3241 (.Y (nx4763), .A0 (scon_3), .A1 (scon_7), .B0 (
                          nx4650), .C0 (nx4639)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_3 (.Q (scon_3), .CK (wb_clk_i), .D (nx4702), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix2391 (.Y (nx4702), .A (scon_3), .B (nx4652), .S0 (nx4651)
                     ) ;
    OAI21_X0P5M_A12TS ix4475 (.Y (nx4652), .A0 (nx4764), .A1 (nx4735), .B0 (
                      nx3024)) ;
    INV_X0P5B_A12TS ix3246 (.Y (nx4764), .A (des1_3)) ;
    OA21A1OI2_X0P5M_A12TS ix4476 (.Y (nx4651), .A0 (nx4629), .A1 (wr_addr_2), .B0 (
                          nx4623), .C0 (nx3037)) ;
    NOR2B_X0P7M_A12TS ix4478 (.Y (nx4650), .AN (scon_6), .B (scon_7)) ;
    NAND2_X0P5A_A12TS ix3252 (.Y (nx4765), .A (nx3003), .B (nx4639)) ;
    NOR2_X0P5A_A12TS ix4480 (.Y (nx4646), .A (nx3003), .B (nx3121)) ;
    INV_X0P5B_A12TS ix3261 (.Y (nx4767), .A (sbuf_txd_0)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_0 (.Q (sbuf_txd_0), .CK (wb_clk_i), .D (
                       nx4711), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4482 (.Y (nx4711), .A (nx4767), .B (nx4768), .S0 (nx4645
                      )) ;
    AOI22_X0P5M_A12TS ix3265 (.Y (nx4768), .A0 (sbuf_txd_1), .A1 (nx3121), .B0 (
                      des1_0), .B1 (nx4647)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_1 (.Q (sbuf_txd_1), .CK (wb_clk_i), .D (
                       nx4700), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4484 (.Y (nx4700), .A (nx4769), .B (nx4770), .S0 (nx4645
                      )) ;
    INV_X0P5B_A12TS ix3269 (.Y (nx4769), .A (sbuf_txd_1)) ;
    AOI222_X0P5M_A12TS ix3271 (.Y (nx4770), .A0 (sbuf_txd_2), .A1 (nx3121), .B0 (
                       des1_1), .B1 (nx4647), .C0 (des1_0), .C1 (nx4646)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_txd_2 (.Q (sbuf_txd_2), .CK (wb_clk_i), .D (
                       nx2470), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4485 (.Y (nx2470), .A (nx4772), .B (nx4774), .S0 (nx4645
                      )) ;
    INV_X0P5B_A12TS ix4486 (.Y (nx4772), .A (sbuf_txd_2)) ;
    AOI222_X0P5M_A12TS ix3277 (.Y (nx4774), .A0 (sbuf_txd_3), .A1 (nx3121), .B0 (
                       des1_2), .B1 (nx4647), .C0 (des1_1), .C1 (nx4646)) ;
    NAND4_X0P5A_A12TS ix3279 (.Y (nx4775), .A (nx4772), .B (nx4769), .C (nx4648)
                      , .D (nx3187)) ;
    NAND3_X0P5A_A12TS ix3281 (.Y (nx4776), .A (nx112), .B (nx568), .C (nx752)) ;
    OAI31_X0P5M_A12TS ix4488 (.Y (nx112), .A0 (wr_addr_2), .A1 (wr_addr_1), .A2 (
                      wr_addr_0), .B0 (nx4623)) ;
    OAI21_X0P5M_A12TS ix569 (.Y (nx568), .A0 (tx_done), .A1 (rx_done), .B0 (
                      nx3037)) ;
    NAND4_X0P5A_A12TS ix753 (.Y (nx752), .A (nx4635), .B (nx4684), .C (nx4778), 
                      .D (scon_5)) ;
    NOR3_X0P5A_A12TS ix4490 (.Y (nx4684), .A (nx32), .B (tx_done), .C (rx_done)
                     ) ;
    INV_X0P5B_A12TS ix3290 (.Y (nx4778), .A (sbuf_rxd_tmp_11)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_11 (.Q (sbuf_rxd_tmp_11), .CK (wb_clk_i)
                       , .D (nx2650), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4492 (.Y (nx2650), .A0 (nx4780), .A1 (nx4795), .B0 (
                          nx4799), .C0 (nx4804)) ;
    AO21A1AI2_X0P5M_A12TS ix3294 (.Y (nx4780), .A0 (nx2331), .A1 (rx_sam_0), .B0 (
                          nx4682), .C0 (rxd_i)) ;
    NOR2_X0P5A_A12TS ix4494 (.Y (nx2331), .A (nx2994), .B (nx4781)) ;
    NAND3_X0P5A_A12TS ix4495 (.Y (nx4781), .A (nx4635), .B (receive), .C (
                      shift_re)) ;
    DFFRPQ_X0P5M_A12TS reg_rx_sam_0 (.Q (rx_sam_0), .CK (wb_clk_i), .D (nx2630)
                       , .R (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4497 (.Y (nx2630), .A (rx_sam_0), .B (rxd_i), .S0 (nx4681
                     )) ;
    NOR2_X0P5A_A12TS ix4498 (.Y (nx4681), .A (re_count_3), .B (nx4793)) ;
    DFFRPQ_X0P5M_A12TS reg_re_count_3 (.Q (re_count_3), .CK (wb_clk_i), .D (
                       nx2620), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix4500 (.Y (nx2620), .A (nx4782)) ;
    AOI32_X0P5M_A12TS ix3304 (.Y (nx4782), .A0 (nx3098), .A1 (nx4680), .A2 (
                      nx2331), .B0 (re_count_3), .B1 (nx4788)) ;
    XNOR2_X0P5M_A12TS ix4501 (.Y (nx4680), .A (re_count_3), .B (nx4783)) ;
    NAND3_X0P5A_A12TS ix4502 (.Y (nx4783), .A (re_count_2), .B (re_count_1), .C (
                      re_count_0)) ;
    DFFRPQ_X0P5M_A12TS reg_re_count_2 (.Q (re_count_2), .CK (wb_clk_i), .D (
                       nx4719), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4503 (.Y (nx4719), .A (nx4784), .B (nx4792), .S0 (nx4788
                      )) ;
    OAI211_X0P5M_A12TS ix3311 (.Y (nx4784), .A0 (nx4679), .A1 (re_count_2), .B0 (
                       nx3098), .C0 (nx4783)) ;
    INV_X0P5B_A12TS ix3314 (.Y (nx4786), .A (re_count_1)) ;
    DFFRPQ_X0P5M_A12TS reg_re_count_1 (.Q (re_count_1), .CK (wb_clk_i), .D (
                       nx2600), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4505 (.Y (nx2600), .A (nx4787), .B (nx4786), .S0 (nx4788
                      )) ;
    OAI211_X0P5M_A12TS ix3318 (.Y (nx4787), .A0 (re_count_0), .A1 (re_count_1), 
                       .B0 (nx3098), .C0 (nx4790)) ;
    DFFRPQ_X0P5M_A12TS reg_re_count_0 (.Q (re_count_0), .CK (wb_clk_i), .D (
                       nx4718), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4506 (.Y (nx4718), .A0 (re_count_0), .A1 (nx644), .A2 (
                      nx4788), .B0 (nx4789)) ;
    NOR2_X0P5A_A12TS ix3322 (.Y (nx4788), .A (nx644), .B (nx2331)) ;
    NAND2_X0P5A_A12TS ix3324 (.Y (nx4789), .A (re_count_0), .B (nx4788)) ;
    NAND2_X0P5A_A12TS ix3326 (.Y (nx4790), .A (re_count_1), .B (re_count_0)) ;
    INV_X0P5B_A12TS ix3330 (.Y (nx4792), .A (re_count_2)) ;
    NOR2_X0P5A_A12TS ix4507 (.Y (nx4682), .A (nx2994), .B (nx3102)) ;
    NAND3_X0P5A_A12TS ix3335 (.Y (nx4795), .A (nx4796), .B (rx_sam_1), .C (
                      nx2331)) ;
    XOR2_X0P5M_A12TS ix3337 (.Y (nx4796), .A (rxd_i), .B (rx_sam_0)) ;
    DFFRPQ_X0P5M_A12TS reg_rx_sam_1 (.Q (rx_sam_1), .CK (wb_clk_i), .D (nx4720)
                       , .R (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4509 (.Y (nx4720), .A (rxd_i), .B (rx_sam_1), .S0 (nx4797
                     )) ;
    NAND3_X0P5A_A12TS ix3343 (.Y (nx4799), .A (rx_done), .B (nx4669), .C (nx636)
                      ) ;
    AOI22_X0P5M_A12TS ix4510 (.Y (nx4669), .A0 (nx3057), .A1 (nx4801), .B0 (
                      nx4803), .B1 (nx2331)) ;
    INV_X0P5B_A12TS ix3346 (.Y (nx4801), .A (scon_4)) ;
    NAND4_X0P5A_A12TS ix3348 (.Y (nx4803), .A (re_count_3), .B (nx4792), .C (
                      nx4786), .D (re_count_0)) ;
    AOI21_X0P5M_A12TS ix637 (.Y (nx636), .A0 (nx3057), .A1 (nx3090), .B0 (nx4671
                      )) ;
    NAND2_X0P5A_A12TS ix3351 (.Y (nx4804), .A (sbuf_rxd_tmp_11), .B (nx4799)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_5 (.Q (scon_5), .CK (wb_clk_i), .D (nx2570), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4511 (.Y (nx2570), .A (nx4668), .B (scon_5), .S0 (nx4808)
                     ) ;
    OAI21_X0P5M_A12TS ix4513 (.Y (nx4668), .A0 (nx4806), .A1 (nx4735), .B0 (
                      nx3024)) ;
    INV_X0P5B_A12TS ix3356 (.Y (nx4806), .A (des1_5)) ;
    AOI21_X0P5M_A12TS ix3358 (.Y (nx4808), .A0 (nx3123), .A1 (nx4631), .B0 (
                      nx4627)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_0 (.Q (sbuf_rxd_tmp_0), .CK (wb_clk_i), 
                       .D (nx4732), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4514 (.Y (nx4732), .A0 (nx4690), .A1 (nx4809), .B0 (
                          nx4799), .C0 (nx4815)) ;
    INV_X0P5B_A12TS ix3362 (.Y (nx4809), .A (sbuf_rxd_tmp_1)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_1 (.Q (sbuf_rxd_tmp_1), .CK (wb_clk_i), 
                       .D (nx2780), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4516 (.Y (nx2780), .A0 (nx4690), .A1 (nx4810), .B0 (
                          nx4799), .C0 (nx4814)) ;
    INV_X0P5B_A12TS ix3366 (.Y (nx4810), .A (sbuf_rxd_tmp_2)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_2 (.Q (sbuf_rxd_tmp_2), .CK (wb_clk_i), 
                       .D (nx4731), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4518 (.Y (nx4731), .A0 (nx4690), .A1 (nx4811), .B0 (
                          nx4799), .C0 (nx4813)) ;
    INV_X0P5B_A12TS ix3370 (.Y (nx4811), .A (sbuf_rxd_tmp_3)) ;
    NAND2_X0P5A_A12TS ix3372 (.Y (nx4813), .A (sbuf_rxd_tmp_2), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix3374 (.Y (nx4814), .A (sbuf_rxd_tmp_1), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix3376 (.Y (nx4815), .A (sbuf_rxd_tmp_0), .B (nx4799)) ;
    INV_X0P5B_A12TS ix3378 (.Y (nx4816), .A (sbuf_rxd_tmp_4)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_4 (.Q (sbuf_rxd_tmp_4), .CK (wb_clk_i), 
                       .D (nx2750), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4519 (.Y (nx2750), .A0 (nx4690), .A1 (nx4820), .B0 (
                          nx4799), .C0 (nx4837)) ;
    INV_X0P5B_A12TS ix3382 (.Y (nx4820), .A (sbuf_rxd_tmp_5)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_5 (.Q (sbuf_rxd_tmp_5), .CK (wb_clk_i), 
                       .D (nx2740), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4522 (.Y (nx2740), .A0 (nx4690), .A1 (nx4821), .B0 (
                          nx4799), .C0 (nx4836)) ;
    INV_X0P5B_A12TS ix3386 (.Y (nx4821), .A (sbuf_rxd_tmp_6)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_6 (.Q (sbuf_rxd_tmp_6), .CK (wb_clk_i), 
                       .D (nx4729), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4523 (.Y (nx4729), .A0 (nx4690), .A1 (nx4822), .B0 (
                          nx4799), .C0 (nx4835)) ;
    INV_X0P5B_A12TS ix3390 (.Y (nx4822), .A (sbuf_rxd_tmp_7)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_7 (.Q (sbuf_rxd_tmp_7), .CK (wb_clk_i), 
                       .D (nx4728), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4524 (.Y (nx4728), .A0 (nx4690), .A1 (nx4824), .B0 (
                          nx4799), .C0 (nx4833)) ;
    INV_X0P5B_A12TS ix3394 (.Y (nx4824), .A (sbuf_rxd_tmp_8)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_8 (.Q (sbuf_rxd_tmp_8), .CK (wb_clk_i), 
                       .D (nx4727), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix4526 (.Y (nx4826), .A0 (sbuf_rxd_tmp_9), .A1 (nx4690
                          ), .B0 (nx644), .C0 (nx4678)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_9 (.Q (sbuf_rxd_tmp_9), .CK (wb_clk_i), 
                       .D (nx4725), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4528 (.Y (nx4725), .A0 (nx4828), .A1 (nx3000), .A2 (
                      nx4799), .B0 (nx4831)) ;
    INV_X0P5B_A12TS ix3405 (.Y (nx4828), .A (sbuf_rxd_tmp_10)) ;
    DFFRPQ_X0P5M_A12TS reg_sbuf_rxd_tmp_10 (.Q (sbuf_rxd_tmp_10), .CK (wb_clk_i)
                       , .D (nx2690), .R (wb_rst_i)) ;
    OAI31_X0P5M_A12TS ix4529 (.Y (nx2690), .A0 (nx4778), .A1 (nx3000), .A2 (
                      nx4799), .B0 (nx4829)) ;
    NAND2_X0P5A_A12TS ix3409 (.Y (nx4829), .A (sbuf_rxd_tmp_10), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix4530 (.Y (nx4831), .A (sbuf_rxd_tmp_9), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix4531 (.Y (nx4833), .A (sbuf_rxd_tmp_7), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix3415 (.Y (nx4835), .A (sbuf_rxd_tmp_6), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix3417 (.Y (nx4836), .A (sbuf_rxd_tmp_5), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix3419 (.Y (nx4837), .A (sbuf_rxd_tmp_4), .B (nx4799)) ;
    NAND2_X0P5A_A12TS ix3421 (.Y (nx4839), .A (sbuf_rxd_tmp_3), .B (nx4799)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_1 (.Q (sbuf_1), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_4), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_2 (.Q (sbuf_2), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_5), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_3 (.Q (sbuf_3), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_6), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_4 (.Q (sbuf_4), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_7), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_5 (.Q (sbuf_5), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_8), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_6 (.Q (sbuf_6), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_9), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_sbuf_rxd_7 (.Q (sbuf_7), .CK (wb_clk_i), .D (
                        sbuf_rxd_tmp_10), .R (wb_rst_i), .SE (rx_done), .SI (
                        sbuf_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_0 (.Q (pcon_0), .CK (wb_clk_i), .D (des1_0), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_1 (.Q (pcon_1), .CK (wb_clk_i), .D (des1_1), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_1)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_2 (.Q (pcon_2), .CK (wb_clk_i), .D (des1_2), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_2)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_3 (.Q (pcon_3), .CK (wb_clk_i), .D (des1_3), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_4 (.Q (pcon_4), .CK (wb_clk_i), .D (des1_4), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_5 (.Q (pcon_5), .CK (wb_clk_i), .D (des1_5), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_pcon_6 (.Q (pcon_6), .CK (wb_clk_i), .D (des1_6), .R (
                        wb_rst_i), .SE (NOT_nx444), .SI (pcon_6)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_1 (.Q (scon_1), .CK (wb_clk_i), .D (nx2980), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4532 (.Y (nx2980), .A (nx4840), .B (nx4841), .S0 (nx4842
                      )) ;
    AOI221_X0P5M_A12TS ix4533 (.Y (nx4840), .A0 (des1_1), .A1 (nx4625), .B0 (
                       tx_done), .B1 (nx3037), .C0 (nx52)) ;
    INV_X0P5B_A12TS ix3442 (.Y (nx4841), .A (scon_1)) ;
    OAI21_X0P5M_A12TS ix3444 (.Y (nx4842), .A0 (nx32), .A1 (tx_done), .B0 (
                      nx4693)) ;
    OAI31_X0P5M_A12TS ix1057 (.Y (nx4693), .A0 (wr_addr_2), .A1 (nx3040), .A2 (
                      wr_addr_1), .B0 (nx4623)) ;
    DFFRPQ_X0P5M_A12TS reg_scon_2 (.Q (scon_2), .CK (wb_clk_i), .D (nx4734), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4535 (.Y (nx4734), .A (nx4843), .B (nx4845), .S0 (nx4846
                      )) ;
    AOI221_X0P5M_A12TS ix3449 (.Y (nx4843), .A0 (des1_2), .A1 (nx4625), .B0 (
                       sbuf_rxd_tmp_11), .B1 (nx4684), .C0 (nx52)) ;
    INV_X0P5B_A12TS ix4536 (.Y (nx4845), .A (scon_2)) ;
    OAI211_X0P5M_A12TS ix4538 (.Y (nx4846), .A0 (nx4635), .A1 (nx32), .B0 (
                       nx1026), .C0 (nx568)) ;
    OAI31_X0P5M_A12TS ix4540 (.Y (nx1026), .A0 (wr_addr_0), .A1 (wr_addr_2), .A2 (
                      nx4848), .B0 (nx4623)) ;
    INV_X0P5B_A12TS ix3456 (.Y (nx4848), .A (wr_addr_1)) ;
    OR2_X0P5M_A12TS ix4541 (.Y (uart_int), .A (scon_0), .B (scon_1)) ;
    DFFSQ_X0P5M_A12TS reg_txd (.Q (txd_o), .CK (wb_clk_i), .D (nx4733), .SN (
                      nx3094)) ;
    MXT2_X0P5M_A12TS ix4542 (.Y (nx4733), .A (nx4691), .B (txd_o), .S0 (nx4851)
                     ) ;
    OAI211_X0P5M_A12TS ix4543 (.Y (nx4691), .A0 (nx3119), .A1 (nx4659), .B0 (
                       nx4850), .C0 (nx3132)) ;
    OAI21_X0P5M_A12TS ix3462 (.Y (nx4850), .A0 (nx4643), .A1 (nx4648), .B0 (
                      sbuf_txd_0)) ;
    NAND3_X0P5A_A12TS ix3464 (.Y (nx4851), .A (nx4640), .B (nx3121), .C (nx4775)
                      ) ;
    INV_X0P5B_A12TS ix4544 (.Y (nx3000), .A (nx4690)) ;
    INV_X0P5B_A12TS ix4546 (.Y (nx3112), .A (nx4684)) ;
    INV_X0P5B_A12TS ix4548 (.Y (nx4679), .A (nx4790)) ;
    INV_X0P5B_A12TS ix645 (.Y (nx644), .A (nx3098)) ;
    INV_X0P5B_A12TS ix3332 (.Y (nx4793), .A (nx2331)) ;
    INV_X0P5B_A12TS ix4549 (.Y (nx4678), .A (nx4799)) ;
    INV_X0P5B_A12TS ix4550 (.Y (nx4677), .A (nx3057)) ;
    INV_X0P5B_A12TS ix4552 (.Y (nx2326), .A (nx3180)) ;
    INV_X0P5B_A12TS ix4555 (.Y (nx3136), .A (nx4665)) ;
    INV_X0P5B_A12TS ix4556 (.Y (nx4648), .A (nx4746)) ;
    INV_X0P5B_A12TS ix4558 (.Y (nx4647), .A (nx4765)) ;
    INV_X0P5B_A12TS ix3250 (.Y (NOT_nx2324), .A (nx4645)) ;
    INV_X0P5B_A12TS ix4559 (.Y (nx3119), .A (nx4643)) ;
    INV_X0P5B_A12TS ix4560 (.Y (nx3132), .A (nx4641)) ;
    INV_X0P5B_A12TS ix4562 (.Y (nx4762), .A (nx4640)) ;
    INV_X0P5B_A12TS ix4563 (.Y (nx4639), .A (nx3121)) ;
    INV_X0P5B_A12TS ix4565 (.Y (nx4636), .A (nx4744)) ;
    INV_X0P5B_A12TS ix4566 (.Y (nx4635), .A (nx3003)) ;
    INV_X0P5B_A12TS ix4567 (.Y (nx52), .A (nx3024)) ;
    INV_X0P5B_A12TS ix33 (.Y (nx32), .A (nx3037)) ;
    INV_X0P5B_A12TS ix4571 (.Y (nx4625), .A (nx4735)) ;
    INV_X0P5B_A12TS ix4573 (.Y (nx4622), .A (nx3027)) ;
    NAND3B_X0P5M_A12TS ix4574 (.Y (nx3027), .AN (nx4739), .B (wr_addr_4), .C (
                       wr_addr_3)) ;
    OR4_X0P5M_A12TS ix4576 (.Y (nx3149), .A (tr_count_3), .B (tr_count_2), .C (
                    tr_count_1), .D (tr_count_0)) ;
    OR4_X0P5M_A12TS ix4578 (.Y (nx4658), .A (sbuf_txd_3), .B (sbuf_txd_4), .C (
                    sbuf_txd_5), .D (sbuf_txd_6)) ;
    AO1B2_X0P5M_A12TS ix4580 (.Y (nx4654), .A0N (nx4763), .B0 (sbuf_txd_10), .B1 (
                      nx3121)) ;
    OR4_X0P5M_A12TS ix4581 (.Y (nx4656), .A (sbuf_txd_7), .B (sbuf_txd_8), .C (
                    sbuf_txd_9), .D (sbuf_txd_10)) ;
    NAND2B_X0P7M_A12TS ix3341 (.Y (nx4797), .AN (re_count_0), .B (nx2331)) ;
    AO1B2_X0P5M_A12TS ix4582 (.Y (nx4727), .A0N (nx4826), .B0 (sbuf_rxd_tmp_8), 
                      .B1 (nx4799)) ;
    TIELO_X1M_A12TS ix4852 (.Y (int_src_7)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_vec_0 (.Q (int_src_1), .CK (wb_clk_i), .D (
                        nx5193), .R (wb_rst_i), .SE (NOT_nx2822), .SI (int_src_1
                        )) ;
    NAND2_X0P5A_A12TS ix4853 (.Y (nx5193), .A (nx5223), .B (nx5268)) ;
    NAND3_X0P5A_A12TS ix3242 (.Y (nx5223), .A (nx5168), .B (ie_7), .C (nx5274)
                      ) ;
    NAND3B_X0P5M_A12TS ix3245 (.Y (nx5224), .AN (ip_4), .B (ie_4), .C (uart_int)
                       ) ;
    DFFRPQ_X0P5M_A12TS reg_ip_4 (.Q (ip_4), .CK (wb_clk_i), .D (nx5213), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4855 (.Y (nx5213), .A (ip_4), .B (nx5143), .S0 (nx5142)
                     ) ;
    OAI21_X0P5M_A12TS ix4856 (.Y (nx5143), .A0 (nx5225), .A1 (nx5226), .B0 (
                      nx5229)) ;
    INV_X0P5B_A12TS ix4857 (.Y (nx5225), .A (des1_4)) ;
    NAND4_X0P5A_A12TS ix4858 (.Y (nx5226), .A (wr_addr_5), .B (wr_addr_4), .C (
                      nx5131), .D (nx5133)) ;
    NOR2_X0P5A_A12TS ix4860 (.Y (nx5131), .A (wr_addr_3), .B (nx5227)) ;
    INV_X0P5B_A12TS ix4861 (.Y (nx5227), .A (wr_addr_2)) ;
    NOR3_X0P5A_A12TS ix4862 (.Y (nx5133), .A (nx5132), .B (wr_bit_r_dup_1790), .C (
                     nx5228)) ;
    NAND2_X0P5A_A12TS ix4863 (.Y (nx5132), .A (wr_addr_1), .B (wr_addr_0)) ;
    NAND3B_X0P5M_A12TS ix3259 (.Y (nx5228), .AN (wr_addr_6), .B (we), .C (
                       wr_addr_7)) ;
    NAND2_X0P5A_A12TS ix4864 (.Y (nx5229), .A (desCy), .B (nx5226)) ;
    OAI31_X0P5M_A12TS ix4865 (.Y (nx5142), .A0 (wr_addr_1), .A1 (wr_addr_0), .A2 (
                      nx5230), .B0 (nx5233)) ;
    NAND2_X0P5A_A12TS ix3264 (.Y (nx5230), .A (wr_addr_2), .B (nx5231)) ;
    NAND2_X0P5A_A12TS ix3266 (.Y (nx5231), .A (nx5226), .B (nx5232)) ;
    NAND4_X0P5A_A12TS ix3268 (.Y (nx5232), .A (wr_addr_3), .B (wr_addr_5), .C (
                      wr_addr_4), .D (nx5130)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_4 (.Q (ie_4), .CK (wb_clk_i), .D (nx5212), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4867 (.Y (nx5212), .A (ie_4), .B (nx5141), .S0 (nx5140)
                     ) ;
    OAI21_X0P5M_A12TS ix4868 (.Y (nx5141), .A0 (nx5225), .A1 (nx5234), .B0 (
                      nx5237)) ;
    NAND3_X0P5A_A12TS ix4869 (.Y (nx5234), .A (nx5136), .B (nx5128), .C (nx5127)
                      ) ;
    NOR3_X0P5A_A12TS ix4872 (.Y (nx5136), .A (wr_bit_r_dup_1790), .B (nx5235), .C (
                     wr_addr_0)) ;
    INV_X0P5B_A12TS ix3282 (.Y (nx5235), .A (wr_addr_5)) ;
    NOR3_X0P5A_A12TS ix4874 (.Y (nx5128), .A (nx5228), .B (wr_addr_4), .C (
                     nx5236)) ;
    INV_X0P5B_A12TS ix3285 (.Y (nx5236), .A (wr_addr_3)) ;
    NOR2_X0P5A_A12TS ix4875 (.Y (nx5127), .A (wr_addr_1), .B (wr_addr_2)) ;
    NAND2_X0P5A_A12TS ix3288 (.Y (nx5237), .A (desCy), .B (nx5234)) ;
    OAI31_X0P5M_A12TS ix4877 (.Y (nx5140), .A0 (wr_addr_1), .A1 (wr_addr_0), .A2 (
                      nx5238), .B0 (nx5241)) ;
    NAND2_X0P5A_A12TS ix3291 (.Y (nx5238), .A (wr_addr_2), .B (nx5239)) ;
    OAI21_X0P5M_A12TS ix4878 (.Y (nx5239), .A0 (nx5240), .A1 (nx5235), .B0 (
                      nx5234)) ;
    NAND2_X0P5A_A12TS ix3295 (.Y (nx5240), .A (wr_bit_r_dup_1790), .B (nx5128)
                      ) ;
    OAI21_X0P5M_A12TS ix4879 (.Y (nx5241), .A0 (nx5240), .A1 (nx5235), .B0 (
                      nx108)) ;
    NAND3B_X0P5M_A12TS ix3300 (.Y (nx5242), .AN (ip_5), .B (ie_5), .C (tc2_int)
                       ) ;
    DFFRPQ_X0P5M_A12TS reg_ip_5 (.Q (ip_5), .CK (wb_clk_i), .D (nx5214), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4880 (.Y (nx5214), .A (ip_5), .B (nx5173), .S0 (nx5172)
                     ) ;
    OAI21_X0P5M_A12TS ix4881 (.Y (nx5173), .A0 (nx5243), .A1 (nx5226), .B0 (
                      nx5229)) ;
    INV_X0P5B_A12TS ix3305 (.Y (nx5243), .A (des1_5)) ;
    OAI21_X0P5M_A12TS ix4882 (.Y (nx5172), .A0 (nx5169), .A1 (nx5230), .B0 (
                      nx5233)) ;
    NAND2_X0P5A_A12TS ix4883 (.Y (nx5169), .A (nx5244), .B (wr_addr_0)) ;
    INV_X0P5B_A12TS ix4885 (.Y (nx5244), .A (wr_addr_1)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_5 (.Q (ie_5), .CK (wb_clk_i), .D (nx2959), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4886 (.Y (nx2959), .A (ie_5), .B (nx5171), .S0 (nx5170)
                     ) ;
    OAI21_X0P5M_A12TS ix4887 (.Y (nx5171), .A0 (nx5243), .A1 (nx5234), .B0 (
                      nx5237)) ;
    OAI21_X0P5M_A12TS ix4891 (.Y (nx5170), .A0 (nx5169), .A1 (nx5238), .B0 (
                      nx5241)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_ie1 (.Q (tcon_3), .CK (wb_clk_i), .D (nx2899), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4892 (.Y (nx2899), .A (tcon_3), .B (nx310), .S0 (nx286)
                     ) ;
    OAI21_X0P5M_A12TS ix4893 (.Y (nx310), .A0 (nx5245), .A1 (nx5246), .B0 (
                      nx5247)) ;
    INV_X0P5B_A12TS ix4894 (.Y (nx5245), .A (des1_3)) ;
    NAND3_X0P5A_A12TS ix3323 (.Y (nx5246), .A (nx5149), .B (nx5128), .C (nx5127)
                      ) ;
    NOR3_X0P5A_A12TS ix4895 (.Y (nx5149), .A (wr_bit_r_dup_1790), .B (wr_addr_5)
                     , .C (wr_addr_0)) ;
    AOI32_X0P5M_A12TS ix4896 (.Y (nx5247), .A0 (nx5248), .A1 (nx5246), .A2 (
                      nx5154), .B0 (desCy), .B1 (nx5146)) ;
    INV_X0P5B_A12TS ix3328 (.Y (nx5248), .A (int1_i)) ;
    AOI21_X0P5M_A12TS ix4898 (.Y (nx5154), .A0 (nx5249), .A1 (tcon_2), .B0 (
                      nx5146)) ;
    INV_X0P5B_A12TS ix3331 (.Y (nx5249), .A (ie1_buff)) ;
    DFFRPQ_X0P5M_A12TS reg_ie1_buff (.Q (ie1_buff), .CK (wb_clk_i), .D (int1_i)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_s_1 (.Q (tcon_2), .CK (wb_clk_i), .D (nx2889), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4899 (.Y (nx2889), .A (tcon_2), .B (nx5153), .S0 (nx268)
                     ) ;
    OAI21_X0P5M_A12TS ix4901 (.Y (nx5153), .A0 (nx5250), .A1 (nx5246), .B0 (
                      nx5251)) ;
    INV_X0P5B_A12TS ix4904 (.Y (nx5250), .A (des1_2)) ;
    NAND2_X0P5A_A12TS ix4905 (.Y (nx5251), .A (desCy), .B (nx5246)) ;
    OA21A1OI2_X0P5M_A12TS ix4907 (.Y (nx268), .A0 (nx5244), .A1 (wr_addr_2), .B0 (
                          nx5129), .C0 (nx5151)) ;
    NOR2_X0P5A_A12TS ix4909 (.Y (nx5129), .A (wr_addr_5), .B (nx5240)) ;
    NOR3_X0P5A_A12TS ix4910 (.Y (nx5146), .A (nx5132), .B (wr_addr_2), .C (
                     nx5252)) ;
    NAND3_X0P5A_A12TS ix4912 (.Y (nx286), .A (nx5246), .B (tcon_2), .C (nx5253)
                      ) ;
    AOI211_X0P5M_A12TS ix3350 (.Y (nx5253), .A0 (nx5248), .A1 (ie1_buff), .B0 (
                       nx5148), .C0 (nx5146)) ;
    NOR3_X0P5A_A12TS ix4913 (.Y (nx5148), .A (nx5254), .B (nx5284), .C (nx5298)
                     ) ;
    NAND2_X0P5A_A12TS ix3353 (.Y (nx5254), .A (int_ack), .B (nx5255)) ;
    AOI32_X0P5M_A12TS ix3355 (.Y (nx5255), .A0 (isrc_0__2), .A1 (int_proc), .A2 (
                      int_dept_0), .B0 (isrc_1__2), .B1 (nx5164)) ;
    DFFRPQ_X0P5M_A12TS reg_isrc_0__2 (.Q (isrc_0__2), .CK (wb_clk_i), .D (nx3099
                       ), .R (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4914 (.Y (nx3099), .A (isrc_0__2), .B (nx5196), .S0 (
                     nx650)) ;
    OAI31_X0P5M_A12TS ix4916 (.Y (nx5196), .A0 (nx5162), .A1 (nx2824), .A2 (
                      nx5174), .B0 (nx3632)) ;
    OAI21_X0P5M_A12TS ix4918 (.Y (nx5162), .A0 (nx5257), .A1 (nx2835), .B0 (
                      nx3553)) ;
    NAND3B_X0P5M_A12TS ix4920 (.Y (nx5257), .AN (ip_2), .B (tcon_3), .C (ie_2)
                       ) ;
    DFFRPQ_X0P5M_A12TS reg_ip_2 (.Q (ip_2), .CK (wb_clk_i), .D (nx2909), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4921 (.Y (nx2909), .A (ip_2), .B (nx5155), .S0 (nx324)) ;
    OAI21_X0P5M_A12TS ix4923 (.Y (nx5155), .A0 (nx5250), .A1 (nx5226), .B0 (
                      nx5229)) ;
    OAI31_X0P5M_A12TS ix4924 (.Y (nx324), .A0 (nx5244), .A1 (wr_addr_0), .A2 (
                      nx5258), .B0 (nx5233)) ;
    NAND2_X0P5A_A12TS ix3367 (.Y (nx5258), .A (nx5227), .B (nx5231)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_2 (.Q (ie_2), .CK (wb_clk_i), .D (nx2919), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4926 (.Y (nx2919), .A (ie_2), .B (nx5157), .S0 (nx5156)
                     ) ;
    OAI21_X0P5M_A12TS ix4927 (.Y (nx5157), .A0 (nx5250), .A1 (nx5234), .B0 (
                      nx5237)) ;
    OAI31_X0P5M_A12TS ix4928 (.Y (nx5156), .A0 (nx5244), .A1 (wr_addr_0), .A2 (
                      nx5259), .B0 (nx5241)) ;
    NAND2_X0P5A_A12TS ix3373 (.Y (nx5259), .A (nx5227), .B (nx5239)) ;
    NAND2_X0P5A_A12TS ix4929 (.Y (nx2835), .A (nx5260), .B (nx3553)) ;
    NAND3B_X0P5M_A12TS ix4930 (.Y (nx5260), .AN (ip_1), .B (tcon_5), .C (ie_1)
                       ) ;
    DFFRPQ_X0P5M_A12TS reg_ip_1 (.Q (ip_1), .CK (wb_clk_i), .D (nx2999), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4931 (.Y (nx2999), .A (ip_1), .B (nx5184), .S0 (nx5183)
                     ) ;
    OAI21_X0P5M_A12TS ix4932 (.Y (nx5184), .A0 (nx5261), .A1 (nx5226), .B0 (
                      nx5229)) ;
    INV_X0P5B_A12TS ix3381 (.Y (nx5261), .A (des1_1)) ;
    OAI21_X0P5M_A12TS ix4933 (.Y (nx5183), .A0 (nx5169), .A1 (nx5258), .B0 (
                      nx5233)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_tf0 (.Q (tcon_5), .CK (wb_clk_i), .D (nx3059), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4935 (.Y (nx3059), .A (tcon_5), .B (nx5191), .S0 (nx788)
                     ) ;
    OAI221_X0P5M_A12TS ix4939 (.Y (nx5191), .A0 (nx5262), .A1 (nx5263), .B0 (
                       nx5243), .B1 (nx5246), .C0 (nx5264)) ;
    INV_X0P5B_A12TS ix4940 (.Y (nx5262), .A (desCy)) ;
    NAND4_X0P5A_A12TS ix3395 (.Y (nx5264), .A (tf0), .B (nx5265), .C (nx5246), .D (
                      nx5263)) ;
    INV_X0P5B_A12TS ix3397 (.Y (nx5265), .A (tf0_buff)) ;
    DFFRPQ_X0P5M_A12TS reg_tf0_buff (.Q (tf0_buff), .CK (wb_clk_i), .D (tf0), .R (
                       wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix789 (.Y (nx788), .A (nx5263), .B (nx5246), .C (nx5266)
                      ) ;
    AOI32_X0P5M_A12TS ix4941 (.Y (nx5266), .A0 (nx5139), .A1 (nx2832), .A2 (
                      nx5298), .B0 (tf0), .B1 (nx5265)) ;
    DFFRPQ_X0P5M_A12TS reg_isrc_0__1 (.Q (isrc_0__1), .CK (wb_clk_i), .D (nx3049
                       ), .R (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4943 (.Y (nx3049), .A (isrc_0__1), .B (nx748), .S0 (nx650
                     )) ;
    OAI31_X0P5M_A12TS ix749 (.Y (nx748), .A0 (nx5267), .A1 (nx5160), .A2 (nx5180
                      ), .B0 (nx5299)) ;
    NAND2_X0P5A_A12TS ix3410 (.Y (nx5267), .A (nx5268), .B (nx3553)) ;
    AO21A1AI2_X0P5M_A12TS ix3412 (.Y (nx5268), .A0 (ie_7), .A1 (nx5202), .B0 (
                          nx5274), .C0 (nx5187)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_7 (.Q (ie_7), .CK (wb_clk_i), .D (nx5216), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4944 (.Y (nx5216), .A (ie_7), .B (nx838), .S0 (nx5192)) ;
    OAI21_X0P5M_A12TS ix839 (.Y (nx838), .A0 (nx5269), .A1 (nx5234), .B0 (nx5237
                      )) ;
    INV_X0P5B_A12TS ix4946 (.Y (nx5269), .A (des1_7)) ;
    OAI21_X0P5M_A12TS ix4947 (.Y (nx5192), .A0 (nx5132), .A1 (nx5238), .B0 (
                      nx5241)) ;
    MXIT2_X0P5M_A12TS ix4949 (.Y (nx5202), .A (int_lev_1__0), .B (int_lev_0__0)
                      , .S0 (int_dept_0)) ;
    DFFRPQ_X0P5M_A12TS reg_int_lev_1__0 (.Q (int_lev_1__0), .CK (wb_clk_i), .D (
                       nx5218), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4950 (.Y (nx5218), .A (nx5270), .B (nx5268), .S0 (nx5195
                      )) ;
    INV_X0P5B_A12TS ix3423 (.Y (nx5270), .A (int_lev_1__0)) ;
    NOR3_X0P5A_A12TS ix4951 (.Y (nx5195), .A (nx5271), .B (int_dept_1), .C (
                     nx5276)) ;
    INV_X0P5B_A12TS ix3426 (.Y (nx5271), .A (int_dept_0)) ;
    DFFRPQ_X0P5M_A12TS reg_int_dept_0 (.Q (int_dept_0), .CK (wb_clk_i), .D (
                       nx2939), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4952 (.Y (nx2939), .A (nx5272), .B (nx5271), .S0 (
                      NOT_nx2836)) ;
    AOI21_X0P5M_A12TS ix3430 (.Y (nx5272), .A0 (nx2822), .A1 (nx2837), .B0 (
                      nx5271)) ;
    NAND2_X0P5A_A12TS ix4953 (.Y (nx2822), .A (int_proc), .B (reti)) ;
    DFFRPQ_X0P5M_A12TS reg_int_proc (.Q (int_proc), .CK (wb_clk_i), .D (nx3079)
                       , .R (wb_rst_i)) ;
    OAI22_X0P5M_A12TS ix4954 (.Y (nx3079), .A0 (nx5273), .A1 (NOT_nx2836), .B0 (
                      nx5274), .B1 (nx5194)) ;
    NOR2_X0P5A_A12TS ix3437 (.Y (NOT_nx2836), .A (nx5193), .B (nx5273)) ;
    INV_X0P5B_A12TS ix4955 (.Y (nx5274), .A (int_proc)) ;
    OA21A1OI2_X0P5M_A12TS ix4956 (.Y (nx5194), .A0 (nx5271), .A1 (int_dept_1), .B0 (
                          nx5273), .C0 (NOT_nx2836)) ;
    SDFFRPQ_X0P5M_A12TS reg_int_dept_1 (.Q (int_dept_1), .CK (wb_clk_i), .D (
                        nx5166), .R (wb_rst_i), .SE (NOT_nx2836), .SI (
                        int_dept_1)) ;
    MXIT2_X0P5M_A12TS ix4958 (.Y (nx5166), .A (nx2837), .B (nx2822), .S0 (nx5165
                      )) ;
    NAND2_X0P5A_A12TS ix4961 (.Y (nx2837), .A (nx2822), .B (nx2824)) ;
    INV_X0P5B_A12TS ix3448 (.Y (nx5275), .A (int_lev_0__0)) ;
    DFFRPQ_X0P5M_A12TS reg_int_lev_0__0 (.Q (int_lev_0__0), .CK (wb_clk_i), .D (
                       nx3139), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix4963 (.Y (nx3139), .A (nx5275), .B (nx5268), .S0 (nx1054
                      )) ;
    NOR3_X0P5A_A12TS ix4964 (.Y (nx1054), .A (nx5276), .B (int_dept_1), .C (
                     int_dept_0)) ;
    OAI21_X0P5M_A12TS ix4965 (.Y (nx5276), .A0 (nx2823), .A1 (nx2824), .B0 (
                      nx2822)) ;
    NOR2_X0P5A_A12TS ix4966 (.Y (nx2823), .A (nx2824), .B (nx5223)) ;
    NAND3_X0P5A_A12TS ix4967 (.Y (nx5278), .A (tcon_3), .B (ip_2), .C (ie_2)) ;
    NAND3_X0P5A_A12TS ix4968 (.Y (nx5279), .A (tcon_7), .B (ip_3), .C (ie_3)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_tf1 (.Q (tcon_7), .CK (wb_clk_i), .D (nx3029), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4969 (.Y (nx3029), .A (tcon_7), .B (nx5190), .S0 (nx5189)
                     ) ;
    OAI221_X0P5M_A12TS ix4971 (.Y (nx5190), .A0 (nx5262), .A1 (nx5280), .B0 (
                       nx5269), .B1 (nx5246), .C0 (nx5281)) ;
    NAND4_X0P5A_A12TS ix4972 (.Y (nx5281), .A (tf1), .B (nx5282), .C (nx5246), .D (
                      nx5280)) ;
    INV_X0P5B_A12TS ix3475 (.Y (nx5282), .A (tf1_buff)) ;
    DFFRPQ_X0P5M_A12TS reg_tf1_buff (.Q (tf1_buff), .CK (wb_clk_i), .D (tf1), .R (
                       wb_rst_i)) ;
    NAND3_X0P5A_A12TS ix4973 (.Y (nx5189), .A (nx5280), .B (nx5246), .C (nx5283)
                      ) ;
    AOI32_X0P5M_A12TS ix3479 (.Y (nx5283), .A0 (nx208), .A1 (nx5284), .A2 (
                      nx5298), .B0 (tf1), .B1 (nx5282)) ;
    AOI32_X0P5M_A12TS ix3484 (.Y (nx5284), .A0 (isrc_0__1), .A1 (int_proc), .A2 (
                      int_dept_0), .B0 (isrc_1__1), .B1 (nx5164)) ;
    DFFRPQ_X0P5M_A12TS reg_isrc_1__1 (.Q (isrc_1__1), .CK (wb_clk_i), .D (nx3039
                       ), .R (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4975 (.Y (nx3039), .A (nx748), .B (isrc_1__1), .S0 (
                     nx5285)) ;
    OAI211_X0P5M_A12TS ix3488 (.Y (nx5285), .A0 (nx912), .A1 (nx5297), .B0 (
                       nx2822), .C0 (nx5188)) ;
    OAI21_X0P5M_A12TS ix913 (.Y (nx912), .A0 (nx2823), .A1 (nx5286), .B0 (nx5296
                      )) ;
    NAND4_X0P5A_A12TS ix3491 (.Y (nx5286), .A (nx584), .B (nx5278), .C (nx5287)
                      , .D (nx5288)) ;
    NOR3_X0P5A_A12TS ix4976 (.Y (nx584), .A (nx2840), .B (nx5182), .C (nx5145)
                     ) ;
    NOR3_X0P5A_A12TS ix4979 (.Y (nx2840), .A (nx2830), .B (nx5279), .C (nx5158)
                     ) ;
    NAND2_X0P5A_A12TS ix4980 (.Y (nx2830), .A (nx5287), .B (nx5288)) ;
    NAND3_X0P5A_A12TS ix3496 (.Y (nx5287), .A (tcon_5), .B (ip_1), .C (ie_1)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_1 (.Q (ie_1), .CK (wb_clk_i), .D (nx3009), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4981 (.Y (nx3009), .A (ie_1), .B (nx5186), .S0 (nx5185)
                     ) ;
    OAI21_X0P5M_A12TS ix4983 (.Y (nx5186), .A0 (nx5261), .A1 (nx5234), .B0 (
                      nx5237)) ;
    OAI21_X0P5M_A12TS ix4985 (.Y (nx5185), .A0 (nx5169), .A1 (nx5259), .B0 (
                      nx5241)) ;
    NAND3_X0P5A_A12TS ix3502 (.Y (nx5288), .A (tcon_1), .B (ip_0), .C (ie_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_ie0 (.Q (tcon_1), .CK (wb_clk_i), .D (nx5217), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4986 (.Y (nx5217), .A (tcon_1), .B (nx5201), .S0 (nx5199)
                     ) ;
    OAI221_X0P5M_A12TS ix4987 (.Y (nx5201), .A0 (nx5262), .A1 (nx5289), .B0 (
                       nx5261), .B1 (nx5246), .C0 (nx5290)) ;
    NAND3_X0P5A_A12TS ix3507 (.Y (nx5289), .A (nx5127), .B (wr_addr_0), .C (
                      nx5129)) ;
    NAND4_X0P5A_A12TS ix4989 (.Y (nx5290), .A (nx5291), .B (nx5246), .C (nx5289)
                      , .D (nx5200)) ;
    INV_X0P5B_A12TS ix3511 (.Y (nx5291), .A (int0_i)) ;
    DFFRPQ_X0P5M_A12TS reg_ie0_buff (.Q (ie0_buff), .CK (wb_clk_i), .D (int0_i)
                       , .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_s_0 (.Q (tcon_0), .CK (wb_clk_i), .D (nx3109), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix4992 (.Y (nx3109), .A (tcon_0), .B (nx5198), .S0 (nx5197)
                     ) ;
    OAI21_X0P5M_A12TS ix4993 (.Y (nx5198), .A0 (nx5292), .A1 (nx5246), .B0 (
                      nx5251)) ;
    INV_X0P5B_A12TS ix3520 (.Y (nx5292), .A (des1_0)) ;
    OA21A1OI2_X0P5M_A12TS ix4994 (.Y (nx5197), .A0 (wr_addr_1), .A1 (wr_addr_2)
                          , .B0 (nx5129), .C0 (nx5151)) ;
    NAND4_X0P5A_A12TS ix4996 (.Y (nx5199), .A (nx5246), .B (tcon_0), .C (nx3523)
                      , .D (nx5289)) ;
    AOI32_X0P5M_A12TS ix4997 (.Y (nx3523), .A0 (nx5139), .A1 (nx5284), .A2 (
                      nx5147), .B0 (nx5291), .B1 (ie0_buff)) ;
    INV_X0P5B_A12TS ix4998 (.Y (nx3526), .A (isrc_0__0)) ;
    DFFRPQ_X0P5M_A12TS reg_isrc_0__0 (.Q (isrc_0__0), .CK (wb_clk_i), .D (nx5215
                       ), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix5000 (.Y (nx5215), .A (nx3526), .B (nx3530), .S0 (nx650)
                      ) ;
    OA21A1OI2_X0P5M_A12TS ix5001 (.Y (nx3530), .A0 (nx5159), .A1 (nx5145), .B0 (
                          nx2824), .C0 (nx5163)) ;
    OAI21_X0P5M_A12TS ix5005 (.Y (nx5159), .A0 (nx5278), .A1 (nx2830), .B0 (
                      nx5288)) ;
    NOR2_X0P5A_A12TS ix5006 (.Y (nx5145), .A (nx3534), .B (nx2829)) ;
    NAND3_X0P5A_A12TS ix5008 (.Y (nx3534), .A (ie_4), .B (uart_int), .C (ip_4)
                      ) ;
    NOR2_X0P5A_A12TS ix5009 (.Y (nx5163), .A (nx2824), .B (nx3537)) ;
    NOR2_X0P5A_A12TS ix5011 (.Y (nx3537), .A (nx5162), .B (nx5160)) ;
    NOR2_X0P5A_A12TS ix5012 (.Y (nx5160), .A (nx5224), .B (nx2834)) ;
    NAND3B_X0P5M_A12TS ix5014 (.Y (nx3541), .AN (ip_3), .B (tcon_7), .C (ie_3)
                       ) ;
    DFFRPQ_X0P5M_A12TS reg_ip_3 (.Q (ip_3), .CK (wb_clk_i), .D (nx2979), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5015 (.Y (nx2979), .A (ip_3), .B (nx5177), .S0 (nx5175)
                     ) ;
    OAI21_X0P5M_A12TS ix5016 (.Y (nx5177), .A0 (nx5245), .A1 (nx5226), .B0 (
                      nx5229)) ;
    OAI21_X0P5M_A12TS ix5018 (.Y (nx5175), .A0 (nx5132), .A1 (nx5258), .B0 (
                      nx5233)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_3 (.Q (ie_3), .CK (wb_clk_i), .D (nx2989), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5020 (.Y (nx2989), .A (ie_3), .B (nx5179), .S0 (nx5178)
                     ) ;
    OAI21_X0P5M_A12TS ix5022 (.Y (nx5179), .A0 (nx5245), .A1 (nx5234), .B0 (
                      nx5237)) ;
    OAI21_X0P5M_A12TS ix5023 (.Y (nx5178), .A0 (nx5132), .A1 (nx5259), .B0 (
                      nx5241)) ;
    NAND3B_X0P5M_A12TS ix5025 (.Y (nx3553), .AN (ip_0), .B (tcon_1), .C (ie_0)
                       ) ;
    DFFRPQ_X0P5M_A12TS reg_ip_0 (.Q (ip_0), .CK (wb_clk_i), .D (nx5211), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5026 (.Y (nx5211), .A (ip_0), .B (nx5135), .S0 (nx5134)
                     ) ;
    OAI21_X0P5M_A12TS ix5027 (.Y (nx5135), .A0 (nx5292), .A1 (nx5226), .B0 (
                      nx5229)) ;
    OAI31_X0P5M_A12TS ix5029 (.Y (nx5134), .A0 (wr_addr_1), .A1 (wr_addr_0), .A2 (
                      nx5258), .B0 (nx5233)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_0 (.Q (ie_0), .CK (wb_clk_i), .D (nx2859), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5031 (.Y (nx2859), .A (ie_0), .B (nx5138), .S0 (nx5137)
                     ) ;
    OAI21_X0P5M_A12TS ix5032 (.Y (nx5138), .A0 (nx5292), .A1 (nx5234), .B0 (
                      nx5237)) ;
    OAI31_X0P5M_A12TS ix5033 (.Y (nx5137), .A0 (wr_addr_1), .A1 (wr_addr_0), .A2 (
                      nx5259), .B0 (nx5241)) ;
    OAI31_X0P5M_A12TS ix5035 (.Y (nx650), .A0 (nx5293), .A1 (nx5277), .A2 (
                      nx5276), .B0 (nx3578)) ;
    AOI21_X0P5M_A12TS ix5036 (.Y (nx5293), .A0 (nx5181), .A1 (nx626), .B0 (
                      nx5167)) ;
    NAND2_X0P5A_A12TS ix5037 (.Y (nx5181), .A (nx3567), .B (nx2823)) ;
    NAND4B_X0P5M_A12TS ix5038 (.Y (nx3567), .AN (nx5162), .B (nx2834), .C (
                       nx3569), .D (nx3571)) ;
    NAND4B_X0P5M_A12TS ix3570 (.Y (nx3569), .AN (ip_1), .B (nx3553), .C (tcon_5)
                       , .D (ie_1)) ;
    NOR2_X0P5A_A12TS ix5039 (.Y (nx5167), .A (int_dept_1), .B (int_dept_0)) ;
    AO21A1AI2_X0P5M_A12TS ix3579 (.Y (nx3578), .A0 (nx5168), .A1 (nx5167), .B0 (
                          nx5181), .C0 (nx2842)) ;
    INV_X0P5B_A12TS ix3586 (.Y (nx5294), .A (isrc_1__0)) ;
    DFFRPQ_X0P5M_A12TS reg_isrc_1__0 (.Q (isrc_1__0), .CK (wb_clk_i), .D (nx2929
                       ), .R (wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix5040 (.Y (nx2929), .A (nx3530), .B (nx5294), .S0 (nx5285
                      )) ;
    NOR3_X0P5A_A12TS ix5041 (.Y (nx5182), .A (nx2829), .B (nx5295), .C (nx5144)
                     ) ;
    NAND3_X0P5A_A12TS ix3594 (.Y (nx5295), .A (ie_5), .B (tc2_int), .C (ip_5)) ;
    OAI211_X0P5M_A12TS ix3596 (.Y (nx5296), .A0 (nx626), .A1 (nx2837), .B0 (
                       nx898), .C0 (nx3537)) ;
    NOR3_X0P5A_A12TS ix5042 (.Y (nx898), .A (nx5180), .B (nx5174), .C (nx496)) ;
    NOR3_X0P5A_A12TS ix5044 (.Y (nx5180), .A (nx2835), .B (nx3541), .C (nx5161)
                     ) ;
    NOR3_X0P5A_A12TS ix497 (.Y (nx496), .A (nx2834), .B (nx5242), .C (nx366)) ;
    NOR2_X0P5A_A12TS ix3610 (.Y (nx5297), .A (nx5271), .B (int_dept_1)) ;
    AOI32_X0P5M_A12TS ix3616 (.Y (nx5298), .A0 (isrc_0__0), .A1 (int_proc), .A2 (
                      int_dept_0), .B0 (isrc_1__0), .B1 (nx5164)) ;
    AOI21_X0P5M_A12TS ix5045 (.Y (nx5165), .A0 (nx5271), .A1 (int_dept_1), .B0 (
                      nx5297)) ;
    NAND4_X0P5A_A12TS ix5046 (.Y (nx3632), .A (nx5287), .B (nx5288), .C (nx2824)
                      , .D (nx5278)) ;
    DFFRPQ_X0P5M_A12TS reg_isrc_1__2 (.Q (isrc_1__2), .CK (wb_clk_i), .D (nx3089
                       ), .R (wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5047 (.Y (nx3089), .A (nx5196), .B (isrc_1__2), .S0 (
                     nx5285)) ;
    DFFRPQ_X0P5M_A12TS reg_ip_6 (.Q (ip_6), .CK (wb_clk_i), .D (nx5221), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3220 (.Y (nx5221), .A (ip_6), .B (nx5209), .S0 (nx5208)
                     ) ;
    OAI21_X0P5M_A12TS ix5048 (.Y (nx5209), .A0 (nx3643), .A1 (nx5226), .B0 (
                      nx5229)) ;
    INV_X0P5B_A12TS ix5049 (.Y (nx3643), .A (des1_6)) ;
    OAI31_X0P5M_A12TS ix5050 (.Y (nx5208), .A0 (nx5244), .A1 (wr_addr_0), .A2 (
                      nx5230), .B0 (nx5233)) ;
    DFFRPQ_X0P5M_A12TS reg_ip_7 (.Q (ip_7), .CK (wb_clk_i), .D (nx5222), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3230 (.Y (nx5222), .A (ip_7), .B (nx5210), .S0 (nx1210)
                     ) ;
    OAI21_X0P5M_A12TS ix5051 (.Y (nx5210), .A0 (nx5269), .A1 (nx5226), .B0 (
                      nx5229)) ;
    OAI21_X0P5M_A12TS ix5052 (.Y (nx1210), .A0 (nx5132), .A1 (nx5230), .B0 (
                      nx5233)) ;
    DFFRPQ_X0P5M_A12TS reg_ie_6 (.Q (ie_6), .CK (wb_clk_i), .D (nx5220), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3210 (.Y (nx5220), .A (ie_6), .B (nx1186), .S0 (nx1182)
                     ) ;
    OAI21_X0P5M_A12TS ix5053 (.Y (nx1186), .A0 (nx3643), .A1 (nx5234), .B0 (
                      nx5237)) ;
    OAI31_X0P5M_A12TS ix1183 (.Y (nx1182), .A0 (nx5244), .A1 (wr_addr_0), .A2 (
                      nx5238), .B0 (nx5241)) ;
    DFFRPQ_X0P5M_A12TS reg_int_vec_3 (.Q (int_src_3), .CK (wb_clk_i), .D (nx3169
                       ), .R (wb_rst_i)) ;
    INV_X0P5B_A12TS ix5054 (.Y (nx3169), .A (nx5300)) ;
    AOI32_X0P5M_A12TS ix5055 (.Y (nx5300), .A0 (nx5193), .A1 (nx3530), .A2 (
                      nx2822), .B0 (int_src_3), .B1 (NOT_nx2822)) ;
    DFFRPQ_X0P5M_A12TS reg_int_vec_4 (.Q (int_src_4), .CK (wb_clk_i), .D (nx3159
                       ), .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5056 (.Y (nx3660), .A0 (nx2823), .A1 (nx5203), .B0 (
                          nx5204), .C0 (nx2822)) ;
    AOI21_X0P5M_A12TS ix5057 (.Y (nx5203), .A0 (nx5257), .A1 (nx3541), .B0 (
                      nx2835)) ;
    AOI211_X0P5M_A12TS ix5058 (.Y (nx5204), .A0 (nx5278), .A1 (nx5279), .B0 (
                       nx5268), .C0 (nx2830)) ;
    DFFRPQ_X0P5M_A12TS reg_int_vec_5 (.Q (int_src_5), .CK (wb_clk_i), .D (nx5219
                       ), .R (wb_rst_i)) ;
    OAI22_X0P5M_A12TS ix5059 (.Y (nx5219), .A0 (nx3666), .A1 (nx2822), .B0 (
                      nx3668), .B1 (NOT_nx2822)) ;
    INV_X0P5B_A12TS ix3667 (.Y (nx3666), .A (int_src_5)) ;
    OA21A1OI2_X0P5M_A12TS ix3669 (.Y (nx3668), .A0 (nx5160), .A1 (nx496), .B0 (
                          nx2823), .C0 (nx1096)) ;
    AOI211_X0P5M_A12TS ix5060 (.Y (nx1096), .A0 (nx3534), .A1 (nx5295), .B0 (
                       nx5268), .C0 (nx2829)) ;
    OR4_X0P5M_A12TS ix5062 (.Y (intr), .A (int_src_1), .B (int_src_3), .C (
                    int_src_4), .D (int_src_5)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_s_3 (.Q (tr1), .CK (wb_clk_i), .D (nx3199), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3200 (.Y (nx3199), .A (nx5207), .B (tr1), .S0 (nx5301)) ;
    OAI21_X0P5M_A12TS ix5063 (.Y (nx5207), .A0 (nx3643), .A1 (nx5246), .B0 (
                      nx5251)) ;
    AOI31_X0P5M_A12TS ix3676 (.Y (nx5301), .A0 (wr_addr_1), .A1 (wr_addr_2), .A2 (
                      nx5129), .B0 (nx5152)) ;
    NOR2_X0P5A_A12TS ix5064 (.Y (nx5152), .A (nx5246), .B (nx5129)) ;
    DFFRPQ_X0P5M_A12TS reg_tcon_s_2 (.Q (tr0), .CK (wb_clk_i), .D (nx3189), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix3190 (.Y (nx3189), .A (tr0), .B (nx5206), .S0 (nx5205)) ;
    OAI21_X0P5M_A12TS ix1157 (.Y (nx5206), .A0 (nx5225), .A1 (nx5246), .B0 (
                      nx5251)) ;
    OA21A1OI2_X0P5M_A12TS ix5065 (.Y (nx5205), .A0 (wr_addr_1), .A1 (nx5227), .B0 (
                          nx5129), .C0 (nx5151)) ;
    INV_X0P5B_A12TS ix3457 (.Y (nx5277), .A (nx5187)) ;
    INV_X0P5B_A12TS ix627 (.Y (nx626), .A (nx5286)) ;
    INV_X0P5B_A12TS ix5066 (.Y (nx3628), .A (nx2840)) ;
    INV_X0P5B_A12TS ix3572 (.Y (nx3571), .A (nx5180)) ;
    INV_X0P5B_A12TS ix5067 (.Y (nx5174), .A (nx3569)) ;
    INV_X0P5B_A12TS ix5068 (.Y (nx5161), .A (nx5257)) ;
    INV_X0P5B_A12TS ix5069 (.Y (nx366), .A (nx5224)) ;
    INV_X0P5B_A12TS ix5070 (.Y (nx5158), .A (nx5278)) ;
    INV_X0P5B_A12TS ix661 (.Y (nx5147), .A (nx5298)) ;
    INV_X0P5B_A12TS ix5071 (.Y (nx2832), .A (nx5284)) ;
    INV_X0P5B_A12TS ix5072 (.Y (nx5144), .A (nx3534)) ;
    INV_X0P5B_A12TS ix959 (.Y (nx5139), .A (nx5254)) ;
    INV_X0P5B_A12TS ix5073 (.Y (nx108), .A (nx5234)) ;
    INV_X0P5B_A12TS ix3435 (.Y (nx5273), .A (nx2822)) ;
    INV_X0P5B_A12TS ix5074 (.Y (nx2824), .A (nx5268)) ;
    INV_X0P5B_A12TS ix5076 (.Y (NOT_nx2822), .A (nx2822)) ;
    INV_X0P5B_A12TS ix5077 (.Y (nx5252), .A (nx5129)) ;
    NAND3B_X0P5M_A12TS ix5078 (.Y (nx5168), .AN (nx2834), .B (nx5224), .C (
                       nx5242)) ;
    NOR2B_X0P7M_A12TS ix5079 (.Y (nx5130), .AN (wr_bit_r_dup_1790), .B (nx5228)
                      ) ;
    NAND2B_X0P7M_A12TS ix3273 (.Y (nx5233), .AN (nx5226), .B (nx5232)) ;
    NOR2B_X0P7M_A12TS ix5080 (.Y (nx5151), .AN (nx5246), .B (nx5129)) ;
    NAND3B_X0P5M_A12TS ix3389 (.Y (nx5263), .AN (nx5169), .B (nx5129), .C (
                       wr_addr_2)) ;
    NAND3B_X0P5M_A12TS ix5081 (.Y (nx2829), .AN (nx2830), .B (nx5278), .C (
                       nx5279)) ;
    NAND3B_X0P5M_A12TS ix3469 (.Y (nx5280), .AN (nx5132), .B (wr_addr_2), .C (
                       nx5129)) ;
    NOR2B_X0P7M_A12TS ix209 (.Y (nx208), .AN (int_ack), .B (nx5255)) ;
    NAND2B_X0P7M_A12TS ix5082 (.Y (nx5200), .AN (ie0_buff), .B (tcon_0)) ;
    NAND3B_X0P5M_A12TS ix825 (.Y (nx2834), .AN (nx2835), .B (nx5257), .C (nx3541
                       )) ;
    NOR2B_X0P7M_A12TS ix5084 (.Y (nx2842), .AN (nx2837), .B (nx5276)) ;
    NOR2B_X0P7M_A12TS ix3590 (.Y (nx5164), .AN (int_proc), .B (int_dept_0)) ;
    NAND3B_X0P5M_A12TS ix5085 (.Y (nx5188), .AN (nx2823), .B (nx5268), .C (
                       nx2822)) ;
    NAND3B_X0P5M_A12TS ix5086 (.Y (nx5187), .AN (nx2829), .B (nx3534), .C (
                       nx5295)) ;
    NAND4B_X0P5M_A12TS ix5087 (.Y (nx5299), .AN (nx5145), .B (nx5288), .C (
                       nx2824), .D (nx3628)) ;
    OAI2XB1_X0P5M_A12TS ix5088 (.Y (nx3159), .A0 (nx2822), .A1N (int_src_4), .B0 (
                        nx3660)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_0 (.Q (th1_0), .CK (wb_clk_i), .D (nx5705), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_0)) ;
    OAI211_X0P5M_A12TS ix5302 (.Y (nx5705), .A0 (nx5768), .A1 (nx2622), .B0 (
                       nx2635), .C0 (nx2866)) ;
    INV_X0P5B_A12TS ix5303 (.Y (nx5768), .A (des1_0)) ;
    INV_X0P5B_A12TS ix5304 (.Y (nx2625), .A (wr_addr_0)) ;
    NAND4_X0P5A_A12TS ix5305 (.Y (nx5769), .A (wr_addr_3), .B (wr_addr_7), .C (
                      nx5659), .D (nx5660)) ;
    NOR2_X0P5A_A12TS ix5306 (.Y (nx5659), .A (wr_addr_6), .B (wr_addr_5)) ;
    NOR3_X0P5A_A12TS ix5307 (.Y (nx5660), .A (wr_bit_r_dup_1790), .B (wr_addr_4)
                     , .C (nx5770)) ;
    INV_X0P5B_A12TS ix5308 (.Y (nx5770), .A (we)) ;
    INV_X0P5B_A12TS ix5309 (.Y (nx2633), .A (wr_addr_1)) ;
    OAI211_X0P5M_A12TS ix5310 (.Y (nx2635), .A0 (nx5676), .A1 (th1_0), .B0 (
                       nx2854), .C0 (nx5680)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_4 (.Q (tl1_4), .CK (wb_clk_i), .D (nx5695), .R (
                        wb_rst_i), .SE (NOT_nx88), .SI (tl1_4)) ;
    OAI211_X0P5M_A12TS ix5311 (.Y (nx5695), .A0 (nx5771), .A1 (nx5772), .B0 (
                       nx2646), .C0 (nx2864)) ;
    INV_X0P5B_A12TS ix5312 (.Y (nx5771), .A (des1_4)) ;
    INV_X0P5B_A12TS ix5314 (.Y (nx5773), .A (wr_addr_2)) ;
    NAND2_X0P5A_A12TS ix5315 (.Y (nx2646), .A (th1_4), .B (nx5682)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_4 (.Q (th1_4), .CK (wb_clk_i), .D (nx348), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_4)) ;
    OAI211_X0P5M_A12TS ix349 (.Y (nx348), .A0 (nx5771), .A1 (nx2622), .B0 (
                       nx5775), .C0 (nx2862)) ;
    OAI211_X0P5M_A12TS ix5316 (.Y (nx5775), .A0 (nx5689), .A1 (th1_4), .B0 (
                       nx2784), .C0 (nx5680)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_3 (.Q (th1_3), .CK (wb_clk_i), .D (nx5690), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_3)) ;
    OAI211_X0P5M_A12TS ix5317 (.Y (nx5690), .A0 (nx2655), .A1 (nx2622), .B0 (
                       nx2657), .C0 (nx2860)) ;
    INV_X0P5B_A12TS ix5318 (.Y (nx2655), .A (des1_3)) ;
    OAI211_X0P5M_A12TS ix5319 (.Y (nx2657), .A0 (nx5685), .A1 (th1_3), .B0 (
                       nx5788), .C0 (nx5680)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_2 (.Q (th1_2), .CK (wb_clk_i), .D (nx5686), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_2)) ;
    OAI211_X0P5M_A12TS ix5320 (.Y (nx5686), .A0 (nx5776), .A1 (nx2622), .B0 (
                       nx5777), .C0 (nx5809)) ;
    INV_X0P5B_A12TS ix5321 (.Y (nx5776), .A (des1_2)) ;
    OAI211_X0P5M_A12TS ix5322 (.Y (nx5777), .A0 (nx5679), .A1 (th1_2), .B0 (
                       nx5808), .C0 (nx5680)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_1 (.Q (th1_1), .CK (wb_clk_i), .D (nx5681), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_1)) ;
    OAI211_X0P5M_A12TS ix5324 (.Y (nx5681), .A0 (nx2669), .A1 (nx2622), .B0 (
                       nx5779), .C0 (nx2852)) ;
    INV_X0P5B_A12TS ix5325 (.Y (nx2669), .A (des1_1)) ;
    OAI211_X0P5M_A12TS ix5326 (.Y (nx5779), .A0 (nx5678), .A1 (th1_1), .B0 (
                       nx5807), .C0 (nx5680)) ;
    NAND2_X0P5A_A12TS ix5327 (.Y (nx5780), .A (tl1_4), .B (nx2169)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_3 (.Q (tl1_3), .CK (wb_clk_i), .D (nx5691), .R (
                        wb_rst_i), .SE (NOT_nx88), .SI (tl1_3)) ;
    OAI211_X0P5M_A12TS ix5328 (.Y (nx5691), .A0 (nx2655), .A1 (nx5772), .B0 (
                       nx5781), .C0 (nx5802)) ;
    NAND2_X0P5A_A12TS ix5329 (.Y (nx5781), .A (th1_3), .B (nx5682)) ;
    NOR2_X0P5A_A12TS ix5330 (.Y (nx5682), .A (nx5663), .B (nx5670)) ;
    NOR3_X0P5A_A12TS ix5332 (.Y (nx5663), .A (nx2683), .B (wr_addr_2), .C (
                     nx2633)) ;
    NAND2_X0P5A_A12TS ix5333 (.Y (nx2683), .A (wr_addr_0), .B (nx5661)) ;
    NAND2_X0P5A_A12TS ix5334 (.Y (nx5670), .A (nx5669), .B (tmod_5)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_7 (.Q (tl1_7), .CK (wb_clk_i), .D (nx5704), .R (
                        wb_rst_i), .SE (NOT_nx120), .SI (tl1_7)) ;
    OAI211_X0P5M_A12TS ix5335 (.Y (nx5704), .A0 (nx5782), .A1 (nx5772), .B0 (
                       nx5783), .C0 (nx2805)) ;
    INV_X0P5B_A12TS ix5336 (.Y (nx5782), .A (des1_7)) ;
    NAND2_X0P5A_A12TS ix5337 (.Y (nx5783), .A (th1_7), .B (nx5682)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_7 (.Q (th1_7), .CK (wb_clk_i), .D (nx5703), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_7)) ;
    OAI222_X0P5M_A12TS ix5338 (.Y (nx5703), .A0 (nx5784), .A1 (nx2799), .B0 (
                       nx5782), .B1 (nx2622), .C0 (nx2801), .C1 (nx5801)) ;
    XOR2_X0P5M_A12TS ix5339 (.Y (nx5784), .A (th1_7), .B (nx5785)) ;
    NAND2_X0P5A_A12TS ix5340 (.Y (nx5785), .A (th1_6), .B (nx5697)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_6 (.Q (th1_6), .CK (wb_clk_i), .D (nx5701), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_6)) ;
    OAI211_X0P5M_A12TS ix5341 (.Y (nx5701), .A0 (nx2706), .A1 (nx2622), .B0 (
                       nx2708), .C0 (nx2786)) ;
    INV_X0P5B_A12TS ix5342 (.Y (nx2706), .A (des1_6)) ;
    OAI211_X0P5M_A12TS ix5343 (.Y (nx2708), .A0 (nx5697), .A1 (th1_6), .B0 (
                       nx5785), .C0 (nx5680)) ;
    SDFFRPQ_X0P5M_A12TS reg_th1_5 (.Q (th1_5), .CK (wb_clk_i), .D (nx5698), .R (
                        wb_rst_i), .SE (NOT_nx106), .SI (th1_5)) ;
    OAI211_X0P5M_A12TS ix5344 (.Y (nx5698), .A0 (nx5787), .A1 (nx2622), .B0 (
                       nx2715), .C0 (nx2727)) ;
    INV_X0P5B_A12TS ix5345 (.Y (nx5787), .A (des1_5)) ;
    OAI211_X0P5M_A12TS ix5346 (.Y (nx2715), .A0 (nx5693), .A1 (th1_5), .B0 (
                       nx5789), .C0 (nx5680)) ;
    NAND2_X0P5A_A12TS ix5347 (.Y (nx5788), .A (th1_3), .B (nx5685)) ;
    NAND2_X0P5A_A12TS ix5348 (.Y (nx5789), .A (th1_5), .B (nx5693)) ;
    NOR2_X0P5A_A12TS ix5350 (.Y (nx5680), .A (tmod_4), .B (nx5662)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_4 (.Q (tmod_4), .CK (wb_clk_i), .D (des1_4), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_4)) ;
    OR3_X0P5M_A12TS ix5351 (.Y (nx5763), .A (nx2683), .B (wr_addr_2), .C (
                    wr_addr_1)) ;
    NOR3_X0P5A_A12TS ix5352 (.Y (nx5662), .A (nx2683), .B (nx5773), .C (
                     wr_addr_1)) ;
    OAI211_X0P5M_A12TS ix5353 (.Y (nx2727), .A0 (nx5692), .A1 (th1_5), .B0 (
                       nx5800), .C0 (nx5674)) ;
    NAND2_X0P5A_A12TS ix5354 (.Y (nx5790), .A (th1_3), .B (nx228)) ;
    NAND2_X0P5A_A12TS ix5355 (.Y (nx5791), .A (th1_1), .B (nx156)) ;
    NAND2_X0P5A_A12TS ix5356 (.Y (nx2736), .A (tl1_7), .B (nx5700)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_6 (.Q (tl1_6), .CK (wb_clk_i), .D (nx5702), .R (
                        wb_rst_i), .SE (NOT_nx120), .SI (tl1_6)) ;
    OAI211_X0P5M_A12TS ix5358 (.Y (nx5702), .A0 (nx2706), .A1 (nx5772), .B0 (
                       nx5792), .C0 (nx2743)) ;
    NAND2_X0P5A_A12TS ix5359 (.Y (nx5792), .A (th1_6), .B (nx5682)) ;
    OAI211_X0P5M_A12TS ix5360 (.Y (nx2743), .A0 (nx2170), .A1 (tl1_6), .B0 (
                       nx2775), .C0 (nx5772)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_5 (.Q (tl1_5), .CK (wb_clk_i), .D (nx5699), .R (
                        wb_rst_i), .SE (NOT_nx120), .SI (tl1_5)) ;
    OAI211_X0P5M_A12TS ix5361 (.Y (nx5699), .A0 (nx5787), .A1 (nx5772), .B0 (
                       nx5793), .C0 (nx5795)) ;
    NAND2_X0P5A_A12TS ix5362 (.Y (nx5793), .A (th1_5), .B (nx5682)) ;
    OAI211_X0P5M_A12TS ix5363 (.Y (nx5795), .A0 (nx5676), .A1 (tl1_5), .B0 (
                       nx2752), .C0 (nx5772)) ;
    NAND2_X0P5A_A12TS ix5364 (.Y (nx2752), .A (tl1_5), .B (nx5676)) ;
    OAI31_X0P5M_A12TS ix5365 (.Y (NOT_nx120), .A0 (tmod_4), .A1 (tmod_5), .A2 (
                      nx5797), .B0 (nx5667)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_5 (.Q (tmod_5), .CK (wb_clk_i), .D (des1_5), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_5)) ;
    NOR2_X0P5A_A12TS ix5366 (.Y (nx5667), .A (nx5662), .B (nx5798)) ;
    NOR2_X0P5A_A12TS ix5367 (.Y (nx5798), .A (nx5666), .B (nx5797)) ;
    AOI211_X0P5M_A12TS ix5368 (.Y (nx5666), .A0 (tmod_7), .A1 (int1_i), .B0 (
                       nx2764), .C0 (nx5799)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_7 (.Q (tmod_7), .CK (wb_clk_i), .D (des1_7), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_7)) ;
    DFFRPQ_X0P5M_A12TS reg_t1_buff (.Q (t1_buff), .CK (wb_clk_i), .D (t1_i), .R (
                       wb_rst_i)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_6 (.Q (tmod_6), .CK (wb_clk_i), .D (des1_6), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_6)) ;
    INV_X0P5B_A12TS ix5369 (.Y (nx2771), .A (pres_ow)) ;
    INV_X0P5B_A12TS ix5370 (.Y (nx5799), .A (tr1)) ;
    NAND2_X0P5A_A12TS ix5371 (.Y (nx2775), .A (tl1_6), .B (nx2170)) ;
    NAND2_X0P5A_A12TS ix5372 (.Y (nx5800), .A (th1_5), .B (nx5692)) ;
    AO21A1AI2_X0P5M_A12TS ix5373 (.Y (NOT_nx106), .A0 (nx2782), .A1 (nx5666), .B0 (
                          nx5662), .C0 (nx5772)) ;
    INV_X0P5B_A12TS ix5374 (.Y (nx2782), .A (tmod_5)) ;
    NAND2_X0P5A_A12TS ix5376 (.Y (nx2784), .A (th1_4), .B (nx5689)) ;
    OAI211_X0P5M_A12TS ix5377 (.Y (nx2786), .A0 (nx5696), .A1 (th1_6), .B0 (
                       nx2797), .C0 (nx5674)) ;
    NAND2_X0P5A_A12TS ix5378 (.Y (nx2789), .A (th1_4), .B (nx5688)) ;
    NAND2_X0P5A_A12TS ix5379 (.Y (nx2792), .A (th1_2), .B (nx5673)) ;
    NAND2_X0P5A_A12TS ix5380 (.Y (nx2795), .A (th1_0), .B (nx5669)) ;
    NAND2_X0P5A_A12TS ix5381 (.Y (nx2797), .A (th1_6), .B (nx5696)) ;
    XOR2_X0P5M_A12TS ix5382 (.Y (nx2801), .A (th1_7), .B (nx2797)) ;
    NAND2_X0P5A_A12TS ix5383 (.Y (nx5801), .A (tmod_4), .B (nx2622)) ;
    OAI211_X0P5M_A12TS ix5384 (.Y (nx2805), .A0 (nx5700), .A1 (tl1_7), .B0 (
                       nx2736), .C0 (nx5772)) ;
    OAI211_X0P5M_A12TS ix5385 (.Y (nx5802), .A0 (nx5684), .A1 (tl1_3), .B0 (
                       nx2848), .C0 (nx5671)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_2 (.Q (tl1_2), .CK (wb_clk_i), .D (nx5687), .R (
                        wb_rst_i), .SE (NOT_nx88), .SI (tl1_2)) ;
    OAI211_X0P5M_A12TS ix5386 (.Y (nx5687), .A0 (nx5776), .A1 (nx5772), .B0 (
                       nx2812), .C0 (nx2814)) ;
    NAND2_X0P5A_A12TS ix5387 (.Y (nx2812), .A (th1_2), .B (nx5682)) ;
    OAI211_X0P5M_A12TS ix5388 (.Y (nx2814), .A0 (nx5668), .A1 (tl1_2), .B0 (
                       nx2846), .C0 (nx5671)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_1 (.Q (tl1_1), .CK (wb_clk_i), .D (nx5683), .R (
                        wb_rst_i), .SE (NOT_nx88), .SI (tl1_1)) ;
    OAI211_X0P5M_A12TS ix5389 (.Y (nx5683), .A0 (nx2669), .A1 (nx5772), .B0 (
                       nx5803), .C0 (nx2821)) ;
    NAND2_X0P5A_A12TS ix5390 (.Y (nx5803), .A (th1_1), .B (nx5682)) ;
    OAI211_X0P5M_A12TS ix5391 (.Y (nx2821), .A0 (tl1_0), .A1 (tl1_1), .B0 (
                       nx2843), .C0 (nx5671)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl1_0 (.Q (tl1_0), .CK (wb_clk_i), .D (nx5706), .R (
                        wb_rst_i), .SE (NOT_nx88), .SI (tl1_0)) ;
    OAI222_X0P5M_A12TS ix5392 (.Y (nx5706), .A0 (nx5768), .A1 (nx5772), .B0 (
                       nx5804), .B1 (nx2827), .C0 (tl1_0), .C1 (nx2831)) ;
    INV_X0P5B_A12TS ix5393 (.Y (nx5804), .A (th1_0)) ;
    NAND2_X0P5A_A12TS ix5394 (.Y (nx2831), .A (nx5772), .B (nx5670)) ;
    OAI21_X0P5M_A12TS ix5395 (.Y (nx5665), .A0 (nx2771), .A1 (tmod_6), .B0 (
                      nx5806)) ;
    NOR2_X0P5A_A12TS ix5396 (.Y (nx5664), .A (nx5663), .B (nx5662)) ;
    NAND2_X0P5A_A12TS ix5398 (.Y (nx2843), .A (tl1_1), .B (tl1_0)) ;
    NAND3_X0P5A_A12TS ix5399 (.Y (nx2846), .A (tl1_2), .B (tl1_1), .C (tl1_0)) ;
    NAND4_X0P5A_A12TS ix5400 (.Y (nx2848), .A (tl1_3), .B (tl1_2), .C (tl1_1), .D (
                      tl1_0)) ;
    NAND2_X0P5A_A12TS ix5401 (.Y (nx5807), .A (th1_1), .B (nx5678)) ;
    OAI211_X0P5M_A12TS ix5402 (.Y (nx2852), .A0 (nx156), .A1 (th1_1), .B0 (
                       nx5791), .C0 (nx5674)) ;
    NAND2_X0P5A_A12TS ix5403 (.Y (nx2854), .A (th1_0), .B (nx5676)) ;
    NAND2_X0P5A_A12TS ix5404 (.Y (nx5808), .A (th1_2), .B (nx5679)) ;
    OAI211_X0P5M_A12TS ix5405 (.Y (nx5809), .A0 (nx5673), .A1 (th1_2), .B0 (
                       nx2792), .C0 (nx5674)) ;
    OAI211_X0P5M_A12TS ix5406 (.Y (nx2860), .A0 (nx228), .A1 (th1_3), .B0 (
                       nx5790), .C0 (nx5674)) ;
    OAI211_X0P5M_A12TS ix5407 (.Y (nx2862), .A0 (nx5688), .A1 (th1_4), .B0 (
                       nx2789), .C0 (nx5674)) ;
    OAI211_X0P5M_A12TS ix5408 (.Y (nx2864), .A0 (nx2169), .A1 (tl1_4), .B0 (
                       nx5780), .C0 (nx5671)) ;
    OAI211_X0P5M_A12TS ix5409 (.Y (nx2866), .A0 (nx5669), .A1 (th1_0), .B0 (
                       nx2795), .C0 (nx5674)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_0 (.Q (th0_0), .CK (wb_clk_i), .D (nx5717), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_0)) ;
    NAND3B_X0P5M_A12TS ix5410 (.Y (nx5717), .AN (nx732), .B (nx2877), .C (nx3135
                       )) ;
    OAI22_X0P5M_A12TS ix733 (.Y (nx732), .A0 (nx5768), .A1 (nx5811), .B0 (th0_0)
                      , .B1 (nx2873)) ;
    NAND4_X0P5A_A12TS ix5411 (.Y (nx5811), .A (wr_addr_2), .B (nx2633), .C (
                      nx2625), .D (nx5661)) ;
    NAND3_X0P5A_A12TS ix5412 (.Y (nx2873), .A (nx5811), .B (tmod_0), .C (tmod_1)
                      ) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_0 (.Q (tmod_0), .CK (wb_clk_i), .D (des1_0), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_0)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_1 (.Q (tmod_1), .CK (wb_clk_i), .D (des1_1), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_1)) ;
    OAI211_X0P5M_A12TS ix5413 (.Y (nx2877), .A0 (nx5715), .A1 (th0_0), .B0 (
                       nx3104), .C0 (nx5713)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_4 (.Q (tl0_4), .CK (wb_clk_i), .D (nx1036), .R (
                        wb_rst_i), .SE (NOT_nx608), .SI (tl0_4)) ;
    OAI211_X0P5M_A12TS ix1037 (.Y (nx1036), .A0 (nx5771), .A1 (nx2882), .B0 (
                       nx5812), .C0 (nx3133)) ;
    NAND4_X0P5A_A12TS ix5414 (.Y (nx2882), .A (nx5773), .B (wr_addr_1), .C (
                      nx2625), .D (nx5661)) ;
    NAND2_X0P5A_A12TS ix5416 (.Y (nx5812), .A (th0_4), .B (nx802)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_4 (.Q (th0_4), .CK (wb_clk_i), .D (nx5742), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_4)) ;
    OAI211_X0P5M_A12TS ix5417 (.Y (nx5742), .A0 (nx5771), .A1 (nx5811), .B0 (
                       nx2888), .C0 (nx3128)) ;
    AO21A1AI2_X0P5M_A12TS ix5418 (.Y (nx2888), .A0 (nx5813), .A1 (nx5713), .B0 (
                          nx5741), .C0 (th0_4)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_3 (.Q (th0_3), .CK (wb_clk_i), .D (nx5734), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_3)) ;
    OAI211_X0P5M_A12TS ix5419 (.Y (nx5734), .A0 (nx2655), .A1 (nx5811), .B0 (
                       nx2895), .C0 (nx5846)) ;
    AO21A1AI2_X0P5M_A12TS ix5420 (.Y (nx2895), .A0 (nx2897), .A1 (nx5713), .B0 (
                          nx5733), .C0 (th0_3)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_2 (.Q (th0_2), .CK (wb_clk_i), .D (nx874), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_2)) ;
    OAI211_X0P5M_A12TS ix5421 (.Y (nx874), .A0 (nx5776), .A1 (nx5811), .B0 (
                       nx2902), .C0 (nx3113)) ;
    AO21A1AI2_X0P5M_A12TS ix5422 (.Y (nx2902), .A0 (nx5815), .A1 (nx5713), .B0 (
                          nx864), .C0 (th0_2)) ;
    NAND2_X0P5A_A12TS ix5423 (.Y (nx5815), .A (th0_2), .B (nx5718)) ;
    DFFRPQ_X0P5M_A12TS reg_th0_1 (.Q (th0_1), .CK (wb_clk_i), .D (nx5764), .R (
                       wb_rst_i)) ;
    OAI21_X0P5M_A12TS ix5424 (.Y (nx5764), .A0 (nx5816), .A1 (NOT_nx680), .B0 (
                      nx5844)) ;
    AOI221_X0P5M_A12TS ix5425 (.Y (nx5816), .A0 (des1_1), .A1 (nx5707), .B0 (
                       th0_1), .B1 (nx5722), .C0 (nx5721)) ;
    OAI222_X0P5M_A12TS ix5426 (.Y (nx5722), .A0 (nx5719), .A1 (nx2873), .B0 (
                       nx5720), .B1 (nx2958), .C0 (nx5718), .C1 (nx3101)) ;
    NAND2_X0P5A_A12TS ix5427 (.Y (nx5817), .A (th0_0), .B (nx2174)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_7 (.Q (tl0_7), .CK (wb_clk_i), .D (nx5758), .R (
                        wb_rst_i), .SE (NOT_nx626), .SI (tl0_7)) ;
    OAI211_X0P5M_A12TS ix5428 (.Y (nx5758), .A0 (nx5782), .A1 (nx2882), .B0 (
                       nx2922), .C0 (nx5843)) ;
    NAND2_X0P5A_A12TS ix5430 (.Y (nx2922), .A (th0_7), .B (nx802)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_7 (.Q (th0_7), .CK (wb_clk_i), .D (nx1232), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_7)) ;
    OAI221_X0P5M_A12TS ix1233 (.Y (nx1232), .A0 (nx2926), .A1 (nx2873), .B0 (
                       nx3092), .B1 (nx2958), .C0 (nx3096)) ;
    XOR2_X0P5M_A12TS ix5431 (.Y (nx2926), .A (th0_7), .B (nx2928)) ;
    NAND2_X0P5A_A12TS ix5432 (.Y (nx2928), .A (th0_6), .B (nx5746)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_6 (.Q (th0_6), .CK (wb_clk_i), .D (nx5756), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_6)) ;
    OAI211_X0P5M_A12TS ix5433 (.Y (nx5756), .A0 (nx2706), .A1 (nx5811), .B0 (
                       nx5818), .C0 (nx3087)) ;
    AO21A1AI2_X0P5M_A12TS ix5434 (.Y (nx5818), .A0 (nx2934), .A1 (nx5713), .B0 (
                          nx5755), .C0 (th0_6)) ;
    SDFFRPQ_X0P5M_A12TS reg_th0_5 (.Q (th0_5), .CK (wb_clk_i), .D (nx1112), .R (
                        wb_rst_i), .SE (NOT_nx680), .SI (th0_5)) ;
    OAI211_X0P5M_A12TS ix1113 (.Y (nx1112), .A0 (nx5787), .A1 (nx5811), .B0 (
                       nx5819), .C0 (nx2960)) ;
    AO21A1AI2_X0P5M_A12TS ix5435 (.Y (nx5819), .A0 (nx5820), .A1 (nx5713), .B0 (
                          nx1102), .C0 (th0_5)) ;
    NOR3_X0P5A_A12TS ix5436 (.Y (nx5713), .A (nx5707), .B (tmod_1), .C (tmod_0)
                     ) ;
    OAI22_X0P5M_A12TS ix1103 (.Y (nx1102), .A0 (nx5746), .A1 (nx2873), .B0 (
                      nx1078), .B1 (nx2958)) ;
    NAND2_X0P5A_A12TS ix5437 (.Y (nx5821), .A (th0_4), .B (nx908)) ;
    NAND3_X0P5A_A12TS ix5438 (.Y (nx2950), .A (th0_2), .B (th0_1), .C (th0_0)) ;
    NAND2_X0P5A_A12TS ix5439 (.Y (nx2953), .A (th0_4), .B (nx5732)) ;
    NAND2_X0P5A_A12TS ix5440 (.Y (nx5822), .A (th0_2), .B (nx5720)) ;
    NAND3B_X0P5M_A12TS ix5442 (.Y (nx2958), .AN (tmod_1), .B (nx5811), .C (
                       tmod_0)) ;
    AOI211_X0P5M_A12TS ix5444 (.Y (nx2960), .A0 (nx5713), .A1 (nx5745), .B0 (
                       nx5748), .C0 (nx5747)) ;
    NOR2_X0P5A_A12TS ix5445 (.Y (nx5745), .A (nx5813), .B (th0_5)) ;
    NOR3_X0P5A_A12TS ix5446 (.Y (nx5748), .A (nx2958), .B (nx2953), .C (th0_5)
                     ) ;
    NOR3_X0P5A_A12TS ix5447 (.Y (nx5747), .A (nx2873), .B (nx5821), .C (th0_5)
                     ) ;
    OAI21_X0P5M_A12TS ix5448 (.Y (NOT_nx680), .A0 (nx672), .A1 (nx5823), .B0 (
                      nx2882)) ;
    OAI22_X0P5M_A12TS ix5449 (.Y (nx672), .A0 (tmod_1), .A1 (nx2968), .B0 (
                      nx5825), .B1 (nx654)) ;
    AOI31_X0P5M_A12TS ix5450 (.Y (nx2968), .A0 (nx586), .A1 (tr0), .A2 (nx5708)
                      , .B0 (nx5823)) ;
    OAI21_X0P5M_A12TS ix5452 (.Y (nx586), .A0 (nx2771), .A1 (tmod_2), .B0 (
                      nx2972)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_2 (.Q (tmod_2), .CK (wb_clk_i), .D (des1_2), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_2)) ;
    DFFRPQ_X0P5M_A12TS reg_t0_buff (.Q (t0_buff), .CK (wb_clk_i), .D (t0_i), .R (
                       wb_rst_i)) ;
    NAND2_X0P5A_A12TS ix5453 (.Y (nx5708), .A (tmod_3), .B (int0_i)) ;
    SDFFRPQ_X0P5M_A12TS reg_tmod_3 (.Q (tmod_3), .CK (wb_clk_i), .D (des1_3), .R (
                        wb_rst_i), .SE (nx5763), .SI (tmod_3)) ;
    NAND2_X0P5A_A12TS ix5454 (.Y (nx5823), .A (nx2882), .B (nx5811)) ;
    AOI21_X0P5M_A12TS ix5455 (.Y (nx5825), .A0 (tr1), .A1 (pres_ow), .B0 (nx5712
                      )) ;
    NAND2_X0P5A_A12TS ix5456 (.Y (nx654), .A (tmod_0), .B (tmod_1)) ;
    OAI22_X0P5M_A12TS ix5457 (.Y (nx5755), .A0 (nx5751), .A1 (nx2873), .B0 (
                      nx5753), .B1 (nx2958)) ;
    NAND2_X0P5A_A12TS ix5458 (.Y (nx5826), .A (th0_5), .B (nx5737)) ;
    NAND2_X0P5A_A12TS ix5459 (.Y (nx5827), .A (th0_3), .B (nx5726)) ;
    NAND2_X0P5A_A12TS ix5460 (.Y (nx2997), .A (th0_1), .B (th0_0)) ;
    NAND2_X0P5A_A12TS ix5461 (.Y (nx5828), .A (th0_5), .B (nx5739)) ;
    NAND2_X0P5A_A12TS ix5462 (.Y (nx5829), .A (th0_3), .B (nx840)) ;
    NAND2_X0P5A_A12TS ix5463 (.Y (nx5830), .A (tl0_7), .B (nx5749)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_6 (.Q (tl0_6), .CK (wb_clk_i), .D (nx1198), .R (
                        wb_rst_i), .SE (NOT_nx626), .SI (tl0_6)) ;
    OAI211_X0P5M_A12TS ix5464 (.Y (nx1198), .A0 (nx2706), .A1 (nx2882), .B0 (
                       nx5831), .C0 (nx3018)) ;
    NAND2_X0P5A_A12TS ix5465 (.Y (nx5831), .A (th0_6), .B (nx802)) ;
    NAND3B_X0P5M_A12TS ix5466 (.Y (nx2177), .AN (tmod_0), .B (tmod_1), .C (
                       nx2174)) ;
    OAI211_X0P5M_A12TS ix5467 (.Y (nx3018), .A0 (nx2180), .A1 (tl0_6), .B0 (
                       nx5841), .C0 (nx5743)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_5 (.Q (tl0_5), .CK (wb_clk_i), .D (nx1122), .R (
                        wb_rst_i), .SE (NOT_nx626), .SI (tl0_5)) ;
    OAI211_X0P5M_A12TS ix1123 (.Y (nx1122), .A0 (nx5787), .A1 (nx2882), .B0 (
                       nx3023), .C0 (nx3025)) ;
    NAND2_X0P5A_A12TS ix5468 (.Y (nx3023), .A (th0_5), .B (nx802)) ;
    OAI211_X0P5M_A12TS ix5470 (.Y (nx3025), .A0 (nx5715), .A1 (tl0_5), .B0 (
                       nx5832), .C0 (nx5743)) ;
    NAND2_X0P5A_A12TS ix5471 (.Y (nx5832), .A (tl0_5), .B (nx5715)) ;
    INV_X0P5B_A12TS ix5472 (.Y (nx5743), .A (nx3030)) ;
    AO21A1AI2_X0P5M_A12TS ix5473 (.Y (nx3030), .A0 (tmod_1), .A1 (nx5830), .B0 (
                          tmod_0), .C0 (nx2882)) ;
    OAI31_X0P5M_A12TS ix5474 (.Y (NOT_nx626), .A0 (tmod_0), .A1 (tmod_1), .A2 (
                      nx5823), .B0 (nx5709)) ;
    NOR2_X0P5A_A12TS ix5475 (.Y (nx5709), .A (nx5707), .B (nx2968)) ;
    NAND2_X0P5A_A12TS ix5476 (.Y (nx3035), .A (tl0_4), .B (nx5729)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_3 (.Q (tl0_3), .CK (wb_clk_i), .D (nx5735), .R (
                        wb_rst_i), .SE (NOT_nx608), .SI (tl0_3)) ;
    OAI211_X0P5M_A12TS ix5477 (.Y (nx5735), .A0 (nx2655), .A1 (nx2882), .B0 (
                       nx5833), .C0 (nx5835)) ;
    NAND2_X0P5A_A12TS ix5478 (.Y (nx5833), .A (th0_3), .B (nx802)) ;
    OAI211_X0P5M_A12TS ix5479 (.Y (nx5835), .A0 (nx2178), .A1 (tl0_3), .B0 (
                       nx5840), .C0 (nx5711)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_2 (.Q (tl0_2), .CK (wb_clk_i), .D (nx5728), .R (
                        wb_rst_i), .SE (NOT_nx608), .SI (tl0_2)) ;
    OAI211_X0P5M_A12TS ix5480 (.Y (nx5728), .A0 (nx5776), .A1 (nx2882), .B0 (
                       nx3047), .C0 (nx5836)) ;
    NAND2_X0P5A_A12TS ix5481 (.Y (nx3047), .A (th0_2), .B (nx802)) ;
    OAI211_X0P5M_A12TS ix5482 (.Y (nx5836), .A0 (nx5710), .A1 (tl0_2), .B0 (
                       nx5839), .C0 (nx5711)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_1 (.Q (tl0_1), .CK (wb_clk_i), .D (nx5723), .R (
                        wb_rst_i), .SE (NOT_nx608), .SI (tl0_1)) ;
    OAI211_X0P5M_A12TS ix5483 (.Y (nx5723), .A0 (nx2669), .A1 (nx2882), .B0 (
                       nx5837), .C0 (nx3056)) ;
    NAND2_X0P5A_A12TS ix5484 (.Y (nx5837), .A (th0_1), .B (nx802)) ;
    OAI211_X0P5M_A12TS ix5485 (.Y (nx3056), .A0 (tl0_0), .A1 (tl0_1), .B0 (
                       nx3078), .C0 (nx5711)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl0_0 (.Q (tl0_0), .CK (wb_clk_i), .D (nx5759), .R (
                        wb_rst_i), .SE (NOT_nx608), .SI (tl0_0)) ;
    OAI222_X0P5M_A12TS ix5486 (.Y (nx5759), .A0 (nx5768), .A1 (nx2882), .B0 (
                       nx3060), .B1 (nx3062), .C0 (tl0_0), .C1 (nx5838)) ;
    INV_X0P5B_A12TS ix5487 (.Y (nx3060), .A (th0_0)) ;
    INV_X0P5B_A12TS ix5488 (.Y (nx3066), .A (tmod_1)) ;
    NAND2_X0P5A_A12TS ix5489 (.Y (nx5838), .A (nx2882), .B (nx2177)) ;
    NAND2_X0P5A_A12TS ix5490 (.Y (nx3078), .A (tl0_1), .B (tl0_0)) ;
    NAND3_X0P5A_A12TS ix5492 (.Y (nx5839), .A (tl0_2), .B (tl0_1), .C (tl0_0)) ;
    NAND4_X0P5A_A12TS ix5493 (.Y (nx5840), .A (tl0_3), .B (tl0_2), .C (tl0_1), .D (
                      tl0_0)) ;
    NAND2_X0P5A_A12TS ix5494 (.Y (nx5841), .A (tl0_6), .B (nx2180)) ;
    AOI211_X0P5M_A12TS ix5495 (.Y (nx3087), .A0 (nx5713), .A1 (nx5750), .B0 (
                       nx1160), .C0 (nx5752)) ;
    NOR2_X0P5A_A12TS ix5496 (.Y (nx5750), .A (nx5820), .B (th0_6)) ;
    NOR3_X0P5A_A12TS ix5497 (.Y (nx1160), .A (nx2958), .B (nx5828), .C (th0_6)
                     ) ;
    NOR3_X0P5A_A12TS ix5498 (.Y (nx5752), .A (nx2873), .B (nx5826), .C (th0_6)
                     ) ;
    XOR2_X0P5M_A12TS ix5499 (.Y (nx3092), .A (th0_7), .B (nx5842)) ;
    NAND2_X0P5A_A12TS ix5500 (.Y (nx5842), .A (th0_6), .B (nx1078)) ;
    AOI22_X0P5M_A12TS ix5501 (.Y (nx3096), .A0 (des1_7), .A1 (nx5707), .B0 (
                      nx5757), .B1 (nx5713)) ;
    XNOR2_X0P5M_A12TS ix5502 (.Y (nx5757), .A (th0_7), .B (nx2934)) ;
    OAI211_X0P5M_A12TS ix5503 (.Y (nx5843), .A0 (nx5749), .A1 (tl0_7), .B0 (
                       nx5830), .C0 (nx5743)) ;
    OAI31_X0P5M_A12TS ix5504 (.Y (nx5721), .A0 (nx3101), .A1 (nx3104), .A2 (
                      th0_1), .B0 (nx3106)) ;
    NAND2_X0P5A_A12TS ix5505 (.Y (nx3104), .A (th0_0), .B (nx5715)) ;
    AOI31_X0P5M_A12TS ix5506 (.Y (nx3106), .A0 (nx5716), .A1 (th0_0), .A2 (
                      nx2997), .B0 (nx764)) ;
    NOR3_X0P5A_A12TS ix765 (.Y (nx764), .A (nx2958), .B (nx5817), .C (th0_1)) ;
    NAND2_X0P5A_A12TS ix5507 (.Y (nx5844), .A (th0_1), .B (NOT_nx680)) ;
    OAI22_X0P5M_A12TS ix5508 (.Y (nx864), .A0 (nx5726), .A1 (nx2873), .B0 (nx840
                      ), .B1 (nx2958)) ;
    AOI211_X0P5M_A12TS ix5510 (.Y (nx3113), .A0 (nx5713), .A1 (nx5725), .B0 (
                       nx846), .C0 (nx5727)) ;
    NOR2_X0P5A_A12TS ix5511 (.Y (nx5725), .A (nx5845), .B (th0_2)) ;
    NOR3_X0P5A_A12TS ix5512 (.Y (nx846), .A (nx2958), .B (nx3006), .C (th0_2)) ;
    NOR3_X0P5A_A12TS ix5513 (.Y (nx5727), .A (nx2873), .B (nx2997), .C (th0_2)
                     ) ;
    OAI22_X0P5M_A12TS ix5514 (.Y (nx5733), .A0 (nx908), .A1 (nx2873), .B0 (
                      nx5732), .B1 (nx2958)) ;
    AOI211_X0P5M_A12TS ix5515 (.Y (nx5846), .A0 (nx5713), .A1 (nx5730), .B0 (
                       nx922), .C0 (nx5731)) ;
    NOR2_X0P5A_A12TS ix5516 (.Y (nx5730), .A (nx5815), .B (th0_3)) ;
    NOR3_X0P5A_A12TS ix923 (.Y (nx922), .A (nx2958), .B (nx5822), .C (th0_3)) ;
    NOR3_X0P5A_A12TS ix5517 (.Y (nx5731), .A (nx2873), .B (nx2950), .C (th0_3)
                     ) ;
    OAI22_X0P5M_A12TS ix5518 (.Y (nx5741), .A0 (nx5737), .A1 (nx2873), .B0 (
                      nx5739), .B1 (nx2958)) ;
    AOI211_X0P5M_A12TS ix5519 (.Y (nx3128), .A0 (nx5713), .A1 (nx5736), .B0 (
                       nx5740), .C0 (nx5738)) ;
    NOR2_X0P5A_A12TS ix5520 (.Y (nx5736), .A (nx2897), .B (th0_4)) ;
    NOR3_X0P5A_A12TS ix5521 (.Y (nx5740), .A (nx2958), .B (nx5829), .C (th0_4)
                     ) ;
    NOR3_X0P5A_A12TS ix991 (.Y (nx5738), .A (nx2873), .B (nx5827), .C (th0_4)) ;
    OAI211_X0P5M_A12TS ix5522 (.Y (nx3133), .A0 (nx5729), .A1 (tl0_4), .B0 (
                       nx3035), .C0 (nx5711)) ;
    OAI211_X0P5M_A12TS ix5524 (.Y (nx3135), .A0 (nx2174), .A1 (th0_0), .B0 (
                       nx5817), .C0 (nx5714)) ;
    OR2_X0P5M_A12TS ix5525 (.Y (tf1), .A (tf1_1), .B (tf1_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tf1_1 (.Q (tf1_1), .CK (wb_clk_i), .D (nx5767), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix5526 (.Y (nx5767), .A (nx5847), .B (nx3147), .S0 (nx5798
                      )) ;
    AO21A1AI2_X0P5M_A12TS ix5527 (.Y (nx5847), .A0 (nx1322), .A1 (nx5762), .B0 (
                          nx5805), .C0 (nx5664)) ;
    MXIT2_X0P5M_A12TS ix5528 (.Y (nx1322), .A (nx5785), .B (nx2797), .S0 (tmod_4
                      )) ;
    NOR2B_X0P7M_A12TS ix5529 (.Y (nx5762), .AN (th1_7), .B (tmod_5)) ;
    INV_X0P5B_A12TS ix5530 (.Y (nx3147), .A (tf1_1)) ;
    DFFRPQ_X0P5M_A12TS reg_tf1_0 (.Q (tf1_0), .CK (wb_clk_i), .D (nx5766), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix5531 (.Y (nx5766), .A (nx5849), .B (nx3155), .S0 (nx5825
                      )) ;
    NAND3_X0P5A_A12TS ix5532 (.Y (nx5849), .A (nx3153), .B (th0_7), .C (nx5751)
                      ) ;
    NOR2_X0P5A_A12TS ix5533 (.Y (nx3153), .A (nx654), .B (nx5823)) ;
    INV_X0P5B_A12TS ix5534 (.Y (nx3155), .A (tf1_0)) ;
    DFFRPQ_X0P5M_A12TS reg_tf0 (.Q (tf0), .CK (wb_clk_i), .D (nx5765), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5536 (.Y (nx5765), .A (nx5761), .B (tf0), .S0 (nx2968)) ;
    OA21A1OI2_X0P5M_A12TS ix5537 (.Y (nx5761), .A0 (nx5830), .A1 (nx654), .B0 (
                          nx3160), .C0 (nx5823)) ;
    AOI31_X0P5M_A12TS ix5538 (.Y (nx3160), .A0 (nx5760), .A1 (nx3066), .A2 (
                      th0_7), .B0 (nx3064)) ;
    MXIT2_X0P5M_A12TS ix5539 (.Y (nx5760), .A (nx2934), .B (nx5842), .S0 (tmod_0
                      )) ;
    INV_X0P5B_A12TS ix5540 (.Y (nx5753), .A (nx5842)) ;
    INV_X0P5B_A12TS ix1147 (.Y (nx5751), .A (nx2928)) ;
    INV_X0P5B_A12TS ix5541 (.Y (nx5749), .A (nx5841)) ;
    INV_X0P5B_A12TS ix5542 (.Y (nx1078), .A (nx5828)) ;
    INV_X0P5B_A12TS ix5543 (.Y (nx5746), .A (nx5826)) ;
    INV_X0P5B_A12TS ix5544 (.Y (nx2180), .A (nx5832)) ;
    INV_X0P5B_A12TS ix5545 (.Y (nx5739), .A (nx2953)) ;
    INV_X0P5B_A12TS ix5546 (.Y (nx5737), .A (nx5821)) ;
    INV_X0P5B_A12TS ix5547 (.Y (nx5732), .A (nx5829)) ;
    INV_X0P5B_A12TS ix909 (.Y (nx908), .A (nx5827)) ;
    INV_X0P5B_A12TS ix5548 (.Y (nx5729), .A (nx5840)) ;
    INV_X0P5B_A12TS ix5549 (.Y (nx840), .A (nx5822)) ;
    INV_X0P5B_A12TS ix5550 (.Y (nx5726), .A (nx2950)) ;
    INV_X0P5B_A12TS ix5551 (.Y (nx2178), .A (nx5839)) ;
    INV_X0P5B_A12TS ix5552 (.Y (nx3062), .A (nx802)) ;
    INV_X0P5B_A12TS ix5554 (.Y (nx3064), .A (nx2177)) ;
    INV_X0P5B_A12TS ix5555 (.Y (nx5720), .A (nx3006)) ;
    INV_X0P5B_A12TS ix5556 (.Y (nx5719), .A (nx2997)) ;
    INV_X0P5B_A12TS ix5557 (.Y (nx5718), .A (nx5845)) ;
    INV_X0P5B_A12TS ix5558 (.Y (nx5716), .A (nx2873)) ;
    INV_X0P5B_A12TS ix5559 (.Y (nx5715), .A (nx3035)) ;
    INV_X0P5B_A12TS ix5560 (.Y (nx5714), .A (nx2958)) ;
    INV_X0P5B_A12TS ix1249 (.Y (nx2174), .A (nx5830)) ;
    INV_X0P5B_A12TS ix5561 (.Y (nx3101), .A (nx5713)) ;
    INV_X0P5B_A12TS ix5562 (.Y (nx5712), .A (nx3153)) ;
    INV_X0P5B_A12TS ix1261 (.Y (nx5711), .A (nx5838)) ;
    INV_X0P5B_A12TS ix5563 (.Y (nx5710), .A (nx3078)) ;
    INV_X0P5B_A12TS ix5564 (.Y (NOT_nx608), .A (nx5709)) ;
    INV_X0P5B_A12TS ix5565 (.Y (nx5707), .A (nx5811)) ;
    INV_X0P5B_A12TS ix5566 (.Y (nx5700), .A (nx2775)) ;
    INV_X0P5B_A12TS ix5567 (.Y (nx5697), .A (nx5789)) ;
    INV_X0P5B_A12TS ix5568 (.Y (nx5696), .A (nx5800)) ;
    INV_X0P5B_A12TS ix5569 (.Y (nx2170), .A (nx2752)) ;
    INV_X0P5B_A12TS ix5570 (.Y (nx5693), .A (nx2784)) ;
    INV_X0P5B_A12TS ix5571 (.Y (nx5692), .A (nx2789)) ;
    INV_X0P5B_A12TS ix5572 (.Y (nx5689), .A (nx5788)) ;
    INV_X0P5B_A12TS ix5573 (.Y (nx5688), .A (nx5790)) ;
    INV_X0P5B_A12TS ix5574 (.Y (nx2169), .A (nx2848)) ;
    INV_X0P5B_A12TS ix5576 (.Y (nx5685), .A (nx5808)) ;
    INV_X0P5B_A12TS ix5577 (.Y (nx228), .A (nx2792)) ;
    INV_X0P5B_A12TS ix5578 (.Y (nx5684), .A (nx2846)) ;
    INV_X0P5B_A12TS ix5579 (.Y (nx2827), .A (nx5682)) ;
    INV_X0P5B_A12TS ix5580 (.Y (nx2799), .A (nx5680)) ;
    INV_X0P5B_A12TS ix5581 (.Y (nx5679), .A (nx5807)) ;
    INV_X0P5B_A12TS ix5582 (.Y (nx5678), .A (nx2854)) ;
    INV_X0P5B_A12TS ix5583 (.Y (nx5676), .A (nx5780)) ;
    INV_X0P5B_A12TS ix5584 (.Y (nx5674), .A (nx5801)) ;
    INV_X0P5B_A12TS ix5585 (.Y (nx5673), .A (nx5791)) ;
    INV_X0P5B_A12TS ix157 (.Y (nx156), .A (nx2795)) ;
    INV_X0P5B_A12TS ix5586 (.Y (nx5671), .A (nx2831)) ;
    INV_X0P5B_A12TS ix5587 (.Y (nx5805), .A (nx5670)) ;
    INV_X0P5B_A12TS ix5588 (.Y (nx5669), .A (nx2736)) ;
    INV_X0P5B_A12TS ix5589 (.Y (nx5668), .A (nx2843)) ;
    INV_X0P5B_A12TS ix5590 (.Y (NOT_nx88), .A (nx5667)) ;
    INV_X0P5B_A12TS ix5591 (.Y (nx2764), .A (nx5665)) ;
    INV_X0P5B_A12TS ix5592 (.Y (nx5797), .A (nx5664)) ;
    INV_X0P5B_A12TS ix5594 (.Y (nx5772), .A (nx5663)) ;
    INV_X0P5B_A12TS ix5595 (.Y (nx2622), .A (nx5662)) ;
    INV_X0P5B_A12TS ix5596 (.Y (nx5661), .A (nx5769)) ;
    NAND3B_X0P5M_A12TS ix5597 (.Y (nx5806), .AN (t1_i), .B (t1_buff), .C (tmod_6
                       )) ;
    NAND2B_X0P7M_A12TS ix5598 (.Y (nx5813), .AN (nx2897), .B (th0_4)) ;
    NAND2B_X0P7M_A12TS ix5599 (.Y (nx2897), .AN (nx5815), .B (th0_3)) ;
    NAND2B_X0P7M_A12TS ix5600 (.Y (nx2934), .AN (nx5820), .B (th0_6)) ;
    NAND2B_X0P7M_A12TS ix5601 (.Y (nx5820), .AN (nx5813), .B (th0_5)) ;
    NAND3B_X0P5M_A12TS ix5602 (.Y (nx2972), .AN (t0_i), .B (t0_buff), .C (tmod_2
                       )) ;
    NAND2B_X0P7M_A12TS ix5603 (.Y (nx3006), .AN (nx5817), .B (th0_1)) ;
    NOR2B_X0P7M_A12TS ix803 (.Y (nx802), .AN (nx2882), .B (nx2177)) ;
    NAND2B_X0P7M_A12TS ix5604 (.Y (nx5845), .AN (nx3104), .B (th0_1)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_0 (.Q (rcap2h_0), .CK (wb_clk_i), .D (nx6204)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5850 (.Y (nx2473), .A0 (th2_0), .A1 (nx6233), .B0 (
                          nx6166), .C0 (nx540)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_0 (.Q (th2_0), .CK (wb_clk_i), .D (nx6167), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_0)) ;
    OAI211_X0P5M_A12TS ix5851 (.Y (nx6167), .A0 (nx6216), .A1 (nx2479), .B0 (
                       nx2491), .C0 (nx2836)) ;
    INV_X0P5B_A12TS ix5852 (.Y (nx6216), .A (des1_0)) ;
    NAND3_X0P5A_A12TS ix5853 (.Y (nx2479), .A (nx6123), .B (wr_addr_2), .C (
                      nx6218)) ;
    NOR2_X0P5A_A12TS ix5854 (.Y (nx6123), .A (wr_bit_r_dup_1790), .B (nx2482)) ;
    NAND4_X0P5A_A12TS ix5856 (.Y (nx2482), .A (wr_addr_7), .B (wr_addr_3), .C (
                      wr_addr_6), .D (nx6121)) ;
    NOR3_X0P5A_A12TS ix5857 (.Y (nx6121), .A (nx6217), .B (wr_addr_5), .C (
                     wr_addr_4)) ;
    INV_X0P5B_A12TS ix5858 (.Y (nx6217), .A (we)) ;
    NOR2_X0P5A_A12TS ix5859 (.Y (nx6218), .A (wr_addr_1), .B (nx2489)) ;
    INV_X0P5B_A12TS ix5860 (.Y (nx2489), .A (wr_addr_0)) ;
    NAND2_X0P5A_A12TS ix5861 (.Y (nx2491), .A (rcap2h_0), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_0 (.Q (t2con_0), .CK (wb_clk_i), .D (nx6191), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5862 (.Y (nx6191), .A (t2con_0), .B (nx6136), .S0 (nx6135
                     )) ;
    OAI21_X0P5M_A12TS ix5863 (.Y (nx6136), .A0 (nx6216), .A1 (nx6219), .B0 (
                      nx6220)) ;
    INV_X0P5B_A12TS ix5864 (.Y (nx2501), .A (wr_addr_2)) ;
    NOR2_X0P5A_A12TS ix5866 (.Y (nx2503), .A (wr_addr_1), .B (wr_addr_0)) ;
    OAI21_X0P5M_A12TS ix5868 (.Y (nx6135), .A0 (nx6125), .A1 (nx6221), .B0 (
                      nx6222)) ;
    INV_X0P5B_A12TS ix5869 (.Y (nx2513), .A (wr_addr_1)) ;
    NAND2_X0P5A_A12TS ix5870 (.Y (nx6221), .A (nx2501), .B (nx6128)) ;
    NAND2_X0P5A_A12TS ix5871 (.Y (nx6128), .A (nx2518), .B (nx6219)) ;
    NAND2_X0P5A_A12TS ix5872 (.Y (nx2518), .A (wr_bit_r_dup_1790), .B (nx6122)
                      ) ;
    NAND2_X0P5A_A12TS ix5873 (.Y (nx6222), .A (nx2518), .B (nx6128)) ;
    DFFRPQ_X0P5M_A12TS reg_neg_trans (.Q (neg_trans), .CK (wb_clk_i), .D (nx6132
                       ), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_t2ex_r (.Q (t2ex_r), .CK (wb_clk_i), .D (t2ex_i), .R (
                       wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_3 (.Q (t2con_3), .CK (wb_clk_i), .D (nx6189), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5874 (.Y (nx6189), .A (t2con_3), .B (nx70), .S0 (nx6130)
                     ) ;
    OAI21_X0P5M_A12TS ix5875 (.Y (nx70), .A0 (nx6223), .A1 (nx6219), .B0 (nx6220
                      )) ;
    INV_X0P5B_A12TS ix5876 (.Y (nx6223), .A (des1_3)) ;
    OAI21_X0P5M_A12TS ix5877 (.Y (nx6130), .A0 (nx6221), .A1 (nx2533), .B0 (
                      nx6222)) ;
    NAND2_X0P5A_A12TS ix5878 (.Y (nx2533), .A (wr_addr_0), .B (wr_addr_1)) ;
    NOR2_X0P5A_A12TS ix5879 (.Y (nx2535), .A (tclk), .B (rclk)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_4 (.Q (tclk), .CK (wb_clk_i), .D (nx6193), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5880 (.Y (nx6193), .A (nx6138), .B (tclk), .S0 (nx6225)
                     ) ;
    OAI21_X0P5M_A12TS ix5881 (.Y (nx6138), .A0 (nx6224), .A1 (nx6219), .B0 (
                      nx6220)) ;
    INV_X0P5B_A12TS ix5882 (.Y (nx6224), .A (des1_4)) ;
    AOI31_X0P5M_A12TS ix5883 (.Y (nx6225), .A0 (nx6128), .A1 (wr_addr_2), .A2 (
                      nx2503), .B0 (nx6129)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_5 (.Q (rclk), .CK (wb_clk_i), .D (nx6192), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5884 (.Y (nx6192), .A (nx6137), .B (rclk), .S0 (nx6227)
                     ) ;
    OAI21_X0P5M_A12TS ix5886 (.Y (nx6137), .A0 (nx2553), .A1 (nx6219), .B0 (
                      nx6220)) ;
    INV_X0P5B_A12TS ix5887 (.Y (nx2553), .A (des1_5)) ;
    AOI31_X0P5M_A12TS ix5888 (.Y (nx6227), .A0 (nx6218), .A1 (wr_addr_2), .A2 (
                      nx6128), .B0 (nx6129)) ;
    NAND2_X0P5A_A12TS ix5889 (.Y (NOT_nx188), .A (nx2479), .B (nx6228)) ;
    NAND3_X0P5A_A12TS ix5890 (.Y (nx6228), .A (nx6123), .B (wr_addr_2), .C (
                      nx2503)) ;
    NOR2_X0P5A_A12TS ix5891 (.Y (nx2563), .A (NOT_nx188), .B (nx6141)) ;
    NOR3_X0P5A_A12TS ix5892 (.Y (nx6141), .A (nx6133), .B (t2con_0), .C (nx6139)
                     ) ;
    NAND2_X0P5A_A12TS ix5893 (.Y (nx6133), .A (neg_trans), .B (t2con_3)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_2 (.Q (t2con_2), .CK (wb_clk_i), .D (nx6195), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5894 (.Y (nx6195), .A (t2con_2), .B (nx6145), .S0 (nx6143
                     )) ;
    OAI21_X0P5M_A12TS ix5895 (.Y (nx6145), .A0 (nx6230), .A1 (nx6219), .B0 (
                      nx6220)) ;
    INV_X0P5B_A12TS ix5896 (.Y (nx6230), .A (des1_2)) ;
    OAI31_X0P5M_A12TS ix5897 (.Y (nx6143), .A0 (nx6221), .A1 (wr_addr_0), .A2 (
                      nx2513), .B0 (nx6222)) ;
    DFFRPQ_X0P5M_A12TS reg_tc2_event (.Q (tc2_event), .CK (wb_clk_i), .D (nx2007
                       ), .R (wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_t2_r (.Q (t2_r), .CK (wb_clk_i), .D (t2_i), .R (
                       wb_rst_i)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_1 (.Q (t2con_1), .CK (wb_clk_i), .D (nx6196), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix5898 (.Y (nx6196), .A (t2con_1), .B (nx218), .S0 (nx6146)
                     ) ;
    OAI21_X0P5M_A12TS ix219 (.Y (nx218), .A0 (nx2585), .A1 (nx6219), .B0 (nx6220
                      )) ;
    INV_X0P5B_A12TS ix5899 (.Y (nx2585), .A (des1_1)) ;
    OAI31_X0P5M_A12TS ix5900 (.Y (nx6146), .A0 (wr_addr_1), .A1 (nx2489), .A2 (
                      nx6221), .B0 (nx6222)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_7 (.Q (th2_7), .CK (wb_clk_i), .D (nx782), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_7)) ;
    OAI211_X0P5M_A12TS ix783 (.Y (nx782), .A0 (nx2592), .A1 (nx2479), .B0 (
                       nx6231), .C0 (nx6237)) ;
    INV_X0P5B_A12TS ix5901 (.Y (nx2592), .A (des1_7)) ;
    NAND2_X0P5A_A12TS ix5902 (.Y (nx6231), .A (rcap2h_7), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_7 (.Q (rcap2h_7), .CK (wb_clk_i), .D (nx6210)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5903 (.Y (nx6232), .A0 (th2_7), .A1 (nx6233), .B0 (
                          nx770), .C0 (nx540)) ;
    NAND4_X0P5A_A12TS ix5904 (.Y (nx6233), .A (wr_addr_0), .B (wr_addr_1), .C (
                      nx2501), .D (nx6123)) ;
    NOR2_X0P5A_A12TS ix771 (.Y (nx770), .A (nx2592), .B (nx6233)) ;
    AOI21_X0P5M_A12TS ix5905 (.Y (nx540), .A0 (nx6235), .A1 (nx6233), .B0 (
                      nx6126)) ;
    NAND4_X0P5A_A12TS ix5906 (.Y (nx6235), .A (neg_trans), .B (t2con_3), .C (
                      t2con_0), .D (nx2535)) ;
    NAND4_X0P5A_A12TS ix5907 (.Y (nx6236), .A (nx2489), .B (nx2501), .C (
                      wr_addr_1), .D (nx6123)) ;
    OAI211_X0P5M_A12TS ix5908 (.Y (nx6237), .A0 (nx6180), .A1 (th2_7), .B0 (
                       nx6269), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_6 (.Q (th2_6), .CK (wb_clk_i), .D (nx6181), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_6)) ;
    OAI211_X0P5M_A12TS ix5909 (.Y (nx6181), .A0 (nx2616), .A1 (nx2479), .B0 (
                       nx2618), .C0 (nx6239)) ;
    INV_X0P5B_A12TS ix5910 (.Y (nx2616), .A (des1_6)) ;
    NAND2_X0P5A_A12TS ix5911 (.Y (nx2618), .A (rcap2h_6), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_6 (.Q (rcap2h_6), .CK (wb_clk_i), .D (nx6209)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5912 (.Y (nx6238), .A0 (th2_6), .A1 (nx6233), .B0 (
                          nx738), .C0 (nx540)) ;
    NOR2_X0P5A_A12TS ix5913 (.Y (nx738), .A (nx2616), .B (nx6233)) ;
    OAI211_X0P5M_A12TS ix5914 (.Y (nx6239), .A0 (nx2022), .A1 (th2_6), .B0 (
                       nx6279), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_5 (.Q (th2_5), .CK (wb_clk_i), .D (nx6179), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_5)) ;
    OAI211_X0P5M_A12TS ix5916 (.Y (nx6179), .A0 (nx2553), .A1 (nx2479), .B0 (
                       nx6240), .C0 (nx2637)) ;
    NAND2_X0P5A_A12TS ix5917 (.Y (nx6240), .A (rcap2h_5), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_5 (.Q (rcap2h_5), .CK (wb_clk_i), .D (nx6208)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5918 (.Y (nx6241), .A0 (th2_5), .A1 (nx6233), .B0 (
                          nx6178), .C0 (nx540)) ;
    NOR2_X0P5A_A12TS ix5919 (.Y (nx6178), .A (nx2553), .B (nx6233)) ;
    OAI211_X0P5M_A12TS ix5920 (.Y (nx2637), .A0 (nx6176), .A1 (th2_5), .B0 (
                       nx6278), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_4 (.Q (th2_4), .CK (wb_clk_i), .D (nx686), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_4)) ;
    OAI211_X0P5M_A12TS ix687 (.Y (nx686), .A0 (nx6224), .A1 (nx2479), .B0 (
                       nx6243), .C0 (nx6245)) ;
    NAND2_X0P5A_A12TS ix5921 (.Y (nx6243), .A (rcap2h_4), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_4 (.Q (rcap2h_4), .CK (wb_clk_i), .D (nx6207)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5922 (.Y (nx6244), .A0 (th2_4), .A1 (nx6233), .B0 (
                          nx6177), .C0 (nx540)) ;
    NOR2_X0P5A_A12TS ix5923 (.Y (nx6177), .A (nx6224), .B (nx6233)) ;
    OAI211_X0P5M_A12TS ix5924 (.Y (nx6245), .A0 (nx6173), .A1 (th2_4), .B0 (
                       nx6277), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_3 (.Q (th2_3), .CK (wb_clk_i), .D (nx6175), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_3)) ;
    OAI211_X0P5M_A12TS ix5925 (.Y (nx6175), .A0 (nx6223), .A1 (nx2479), .B0 (
                       nx6246), .C0 (nx6248)) ;
    NAND2_X0P5A_A12TS ix5926 (.Y (nx6246), .A (rcap2h_3), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_3 (.Q (rcap2h_3), .CK (wb_clk_i), .D (nx6206)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5927 (.Y (nx6247), .A0 (th2_3), .A1 (nx6233), .B0 (
                          nx6174), .C0 (nx540)) ;
    NOR2_X0P5A_A12TS ix5928 (.Y (nx6174), .A (nx6223), .B (nx6233)) ;
    OAI211_X0P5M_A12TS ix5929 (.Y (nx6248), .A0 (nx6170), .A1 (th2_3), .B0 (
                       nx2828), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_2 (.Q (th2_2), .CK (wb_clk_i), .D (nx6172), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_2)) ;
    OAI211_X0P5M_A12TS ix5930 (.Y (nx6172), .A0 (nx6230), .A1 (nx2479), .B0 (
                       nx6249), .C0 (nx2673)) ;
    NAND2_X0P5A_A12TS ix5931 (.Y (nx6249), .A (rcap2h_2), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_2 (.Q (rcap2h_2), .CK (wb_clk_i), .D (nx6205)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5932 (.Y (nx6251), .A0 (th2_2), .A1 (nx6233), .B0 (
                          nx6171), .C0 (nx540)) ;
    NOR2_X0P5A_A12TS ix5933 (.Y (nx6171), .A (nx6230), .B (nx6233)) ;
    OAI211_X0P5M_A12TS ix5934 (.Y (nx2673), .A0 (nx2018), .A1 (th2_2), .B0 (
                       nx6276), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_th2_1 (.Q (th2_1), .CK (wb_clk_i), .D (nx6169), .R (
                        wb_rst_i), .SE (NOT_nx264), .SI (th2_1)) ;
    OAI211_X0P5M_A12TS ix5936 (.Y (nx6169), .A0 (nx2585), .A1 (nx2479), .B0 (
                       nx2678), .C0 (nx2685)) ;
    NAND2_X0P5A_A12TS ix5937 (.Y (nx2678), .A (rcap2h_1), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2h_1 (.Q (rcap2h_1), .CK (wb_clk_i), .D (nx2271)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5938 (.Y (nx2682), .A0 (th2_1), .A1 (nx6233), .B0 (
                          nx6168), .C0 (nx540)) ;
    NOR2_X0P5A_A12TS ix5939 (.Y (nx6168), .A (nx2585), .B (nx6233)) ;
    OAI211_X0P5M_A12TS ix5940 (.Y (nx2685), .A0 (nx6165), .A1 (th2_1), .B0 (
                       nx6273), .C0 (nx2009)) ;
    NAND2_X0P5A_A12TS ix5941 (.Y (nx6252), .A (tl2_7), .B (nx6159)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_7 (.Q (tl2_7), .CK (wb_clk_i), .D (nx6163), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_7)) ;
    OAI211_X0P5M_A12TS ix5942 (.Y (nx6163), .A0 (nx2592), .A1 (nx6228), .B0 (
                       nx6253), .C0 (nx2705)) ;
    NAND2_X0P5A_A12TS ix5943 (.Y (nx6253), .A (rcap2l_7), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_7 (.Q (rcap2l_7), .CK (wb_clk_i), .D (nx6203)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5944 (.Y (nx6255), .A0 (tl2_7), .A1 (nx6236), .B0 (
                          nx6162), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5945 (.Y (nx6162), .A (nx2592), .B (nx6236)) ;
    AOI21_X0P5M_A12TS ix5946 (.Y (nx6140), .A0 (nx6235), .A1 (nx6236), .B0 (
                      nx6124)) ;
    OAI211_X0P5M_A12TS ix5947 (.Y (nx2705), .A0 (nx6159), .A1 (tl2_7), .B0 (
                       nx6252), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_6 (.Q (tl2_6), .CK (wb_clk_i), .D (nx6160), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_6)) ;
    OAI211_X0P5M_A12TS ix5948 (.Y (nx6160), .A0 (nx2616), .A1 (nx6228), .B0 (
                       nx6256), .C0 (nx2717)) ;
    NAND2_X0P5A_A12TS ix5949 (.Y (nx6256), .A (rcap2l_6), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_6 (.Q (rcap2l_6), .CK (wb_clk_i), .D (nx6202)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5950 (.Y (nx6257), .A0 (tl2_6), .A1 (nx6236), .B0 (
                          nx476), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5951 (.Y (nx476), .A (nx2616), .B (nx6236)) ;
    OAI211_X0P5M_A12TS ix5952 (.Y (nx2717), .A0 (nx2014), .A1 (tl2_6), .B0 (
                       nx6272), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_5 (.Q (tl2_5), .CK (wb_clk_i), .D (nx6158), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_5)) ;
    OAI211_X0P5M_A12TS ix5953 (.Y (nx6158), .A0 (nx2553), .A1 (nx6228), .B0 (
                       nx6258), .C0 (nx2729)) ;
    NAND2_X0P5A_A12TS ix5954 (.Y (nx6258), .A (rcap2l_5), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_5 (.Q (rcap2l_5), .CK (wb_clk_i), .D (nx6201)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5956 (.Y (nx6259), .A0 (tl2_5), .A1 (nx6236), .B0 (
                          nx6157), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5958 (.Y (nx6157), .A (nx2553), .B (nx6236)) ;
    OAI211_X0P5M_A12TS ix5959 (.Y (nx2729), .A0 (nx6155), .A1 (tl2_5), .B0 (
                       nx2815), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_4 (.Q (tl2_4), .CK (wb_clk_i), .D (nx6156), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_4)) ;
    OAI211_X0P5M_A12TS ix5960 (.Y (nx6156), .A0 (nx6224), .A1 (nx6228), .B0 (
                       nx6260), .C0 (nx6261)) ;
    NAND2_X0P5A_A12TS ix5961 (.Y (nx6260), .A (rcap2l_4), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_4 (.Q (rcap2l_4), .CK (wb_clk_i), .D (nx6200)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5962 (.Y (nx2738), .A0 (tl2_4), .A1 (nx6236), .B0 (
                          nx412), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix413 (.Y (nx412), .A (nx6224), .B (nx6236)) ;
    OAI211_X0P5M_A12TS ix5963 (.Y (nx6261), .A0 (nx2012), .A1 (tl2_4), .B0 (
                       nx6271), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_3 (.Q (tl2_3), .CK (wb_clk_i), .D (nx6154), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_3)) ;
    OAI211_X0P5M_A12TS ix5964 (.Y (nx6154), .A0 (nx6223), .A1 (nx6228), .B0 (
                       nx6262), .C0 (nx2753)) ;
    NAND2_X0P5A_A12TS ix5965 (.Y (nx6262), .A (rcap2l_3), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_3 (.Q (rcap2l_3), .CK (wb_clk_i), .D (nx6199)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5966 (.Y (nx6263), .A0 (tl2_3), .A1 (nx6236), .B0 (
                          nx6153), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5967 (.Y (nx6153), .A (nx6223), .B (nx6236)) ;
    OAI211_X0P5M_A12TS ix5968 (.Y (nx2753), .A0 (nx6151), .A1 (tl2_3), .B0 (
                       nx2811), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_2 (.Q (tl2_2), .CK (wb_clk_i), .D (nx360), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_2)) ;
    OAI211_X0P5M_A12TS ix5969 (.Y (nx360), .A0 (nx6230), .A1 (nx6228), .B0 (
                       nx2758), .C0 (nx2765)) ;
    NAND2_X0P5A_A12TS ix5970 (.Y (nx2758), .A (rcap2l_2), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_2 (.Q (rcap2l_2), .CK (wb_clk_i), .D (nx6198)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5971 (.Y (nx2762), .A0 (tl2_2), .A1 (nx6236), .B0 (
                          nx6152), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5972 (.Y (nx6152), .A (nx6230), .B (nx6236)) ;
    OAI211_X0P5M_A12TS ix5973 (.Y (nx2765), .A0 (nx2008), .A1 (tl2_2), .B0 (
                       nx6270), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_1 (.Q (tl2_1), .CK (wb_clk_i), .D (nx6150), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_1)) ;
    OAI211_X0P5M_A12TS ix5974 (.Y (nx6150), .A0 (nx2585), .A1 (nx6228), .B0 (
                       nx6264), .C0 (nx6265)) ;
    NAND2_X0P5A_A12TS ix5976 (.Y (nx6264), .A (rcap2l_1), .B (nx322)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_1 (.Q (rcap2l_1), .CK (wb_clk_i), .D (nx6197)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5977 (.Y (nx2774), .A0 (tl2_1), .A1 (nx6236), .B0 (
                          nx6149), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5978 (.Y (nx6149), .A (nx2585), .B (nx6236)) ;
    OAI211_X0P5M_A12TS ix5979 (.Y (nx6265), .A0 (tl2_0), .A1 (tl2_1), .B0 (
                       nx2806), .C0 (nx2009)) ;
    SDFFRPQ_X0P5M_A12TS reg_tl2_0 (.Q (tl2_0), .CK (wb_clk_i), .D (nx6182), .R (
                        wb_rst_i), .SE (NOT_nx252), .SI (tl2_0)) ;
    OAI222_X0P5M_A12TS ix5980 (.Y (nx6182), .A0 (nx2781), .A1 (nx6267), .B0 (
                       nx6216), .B1 (nx6228), .C0 (tl2_0), .C1 (nx2802)) ;
    INV_X0P5B_A12TS ix5981 (.Y (nx2781), .A (rcap2l_0)) ;
    DFFRPQ_X0P5M_A12TS reg_rcap2l_0 (.Q (rcap2l_0), .CK (wb_clk_i), .D (nx6211)
                       , .R (wb_rst_i)) ;
    AO21A1AI2_X0P5M_A12TS ix5982 (.Y (nx6266), .A0 (tl2_0), .A1 (nx6236), .B0 (
                          nx6183), .C0 (nx6140)) ;
    NOR2_X0P5A_A12TS ix5983 (.Y (nx6183), .A (nx6216), .B (nx6236)) ;
    AOI22_X0P5M_A12TS ix5984 (.Y (nx6267), .A0 (nx6141), .A1 (nx6142), .B0 (
                      nx6148), .B1 (nx2798)) ;
    AO21A1AI2_X0P5M_A12TS ix5985 (.Y (nx6268), .A0 (t2con_1), .A1 (tc2_event), .B0 (
                          nx6147), .C0 (t2con_2)) ;
    NOR2B_X0P7M_A12TS ix5986 (.Y (nx6147), .AN (pres_ow), .B (t2con_1)) ;
    AOI21_X0P5M_A12TS ix5987 (.Y (nx2798), .A0 (t2con_0), .A1 (nx2535), .B0 (
                      nx6269)) ;
    NAND2_X0P5A_A12TS ix5988 (.Y (nx6269), .A (th2_7), .B (nx6180)) ;
    AO1B2_X0P5M_A12TS ix5989 (.Y (NOT_nx252), .A0N (nx2479), .B0 (nx6268), .B1 (
                      nx2563)) ;
    NAND2_X0P5A_A12TS ix5990 (.Y (nx2806), .A (tl2_1), .B (tl2_0)) ;
    NOR2_X0P5A_A12TS ix799 (.Y (nx2009), .A (nx6229), .B (nx2798)) ;
    NAND3_X0P5A_A12TS ix5991 (.Y (nx6270), .A (tl2_2), .B (tl2_1), .C (tl2_0)) ;
    NAND4_X0P5A_A12TS ix5992 (.Y (nx2811), .A (tl2_3), .B (tl2_2), .C (tl2_1), .D (
                      tl2_0)) ;
    NAND2_X0P5A_A12TS ix5993 (.Y (nx6271), .A (tl2_4), .B (nx2012)) ;
    NAND2_X0P5A_A12TS ix5994 (.Y (nx2815), .A (tl2_5), .B (nx6155)) ;
    NAND2_X0P5A_A12TS ix5996 (.Y (nx6272), .A (tl2_6), .B (nx2014)) ;
    NAND2_X0P5A_A12TS ix5997 (.Y (nx6273), .A (th2_1), .B (nx6165)) ;
    AO1B2_X0P5M_A12TS ix5998 (.Y (NOT_nx264), .A0N (nx6228), .B0 (nx6268), .B1 (
                      nx2563)) ;
    NAND2_X0P5A_A12TS ix5999 (.Y (nx6275), .A (th2_0), .B (nx6161)) ;
    NAND2_X0P5A_A12TS ix6000 (.Y (nx6276), .A (th2_2), .B (nx2018)) ;
    NAND2_X0P5A_A12TS ix6001 (.Y (nx2828), .A (th2_3), .B (nx6170)) ;
    NAND2_X0P5A_A12TS ix6002 (.Y (nx6277), .A (th2_4), .B (nx6173)) ;
    NAND2_X0P5A_A12TS ix6003 (.Y (nx6278), .A (th2_5), .B (nx6176)) ;
    NAND2_X0P5A_A12TS ix6004 (.Y (nx6279), .A (th2_6), .B (nx2022)) ;
    OAI211_X0P5M_A12TS ix6005 (.Y (nx2836), .A0 (nx6161), .A1 (th2_0), .B0 (
                       nx6275), .C0 (nx2009)) ;
    NOR2_X0P5A_A12TS ix6006 (.Y (nx6166), .A (nx6216), .B (nx6233)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_6 (.Q (t2con_6), .CK (wb_clk_i), .D (nx6215), .R (
                       wb_rst_i)) ;
    MXIT2_X0P5M_A12TS ix6007 (.Y (nx6215), .A (nx6280), .B (nx6281), .S0 (nx6188
                      )) ;
    INV_X0P5B_A12TS ix6008 (.Y (nx6280), .A (t2con_6)) ;
    AOI211_X0P5M_A12TS ix6009 (.Y (nx6281), .A0 (des1_6), .A1 (nx6127), .B0 (
                       nx6186), .C0 (nx6131)) ;
    NOR3_X0P5A_A12TS ix6010 (.Y (nx6186), .A (nx6133), .B (tf2_set), .C (nx6128)
                     ) ;
    SDFFRPQ_X0P5M_A12TS reg_tf2_set (.Q (tf2_set), .CK (wb_clk_i), .D (nx842), .R (
                        wb_rst_i), .SE (NOT_nx188), .SI (tf2_set)) ;
    NOR3_X0P5A_A12TS ix6011 (.Y (nx842), .A (nx6229), .B (nx6269), .C (nx6139)
                     ) ;
    AOI21_X0P5M_A12TS ix6012 (.Y (nx6188), .A0 (nx6282), .A1 (nx6222), .B0 (
                      nx854)) ;
    AOI32_X0P5M_A12TS ix6013 (.Y (nx6282), .A0 (nx2489), .A1 (wr_addr_1), .A2 (
                      nx896), .B0 (nx2853), .B1 (nx2518)) ;
    AOI21_X0P5M_A12TS ix6014 (.Y (nx896), .A0 (nx6226), .A1 (tf2_set), .B0 (
                      nx2501)) ;
    INV_X0P5B_A12TS ix6016 (.Y (nx2853), .A (tf2_set)) ;
    AOI211_X0P5M_A12TS ix6017 (.Y (nx854), .A0 (neg_trans), .A1 (t2con_3), .B0 (
                       tf2_set), .C0 (nx6128)) ;
    DFFRPQ_X0P5M_A12TS reg_t2con_7 (.Q (t2con_7), .CK (wb_clk_i), .D (nx6213), .R (
                       wb_rst_i)) ;
    MXT2_X0P5M_A12TS ix6018 (.Y (nx6213), .A (nx6187), .B (t2con_7), .S0 (nx6283
                     )) ;
    OAI221_X0P5M_A12TS ix6019 (.Y (nx6187), .A0 (nx2592), .A1 (nx6219), .B0 (
                       nx2853), .B1 (nx6128), .C0 (nx6220)) ;
    OAI22_X0P5M_A12TS ix6020 (.Y (nx6283), .A0 (nx6185), .A1 (nx2518), .B0 (
                      tf2_set), .B1 (nx6128)) ;
    NOR2_X0P5A_A12TS ix6021 (.Y (nx6185), .A (nx2501), .B (nx2533)) ;
    OR2_X0P5M_A12TS ix6022 (.Y (tc2_int), .A (t2con_6), .B (t2con_7)) ;
    DFFRPQ_X0P5M_A12TS reg_brate2 (.Q (brate2), .CK (wb_clk_i), .D (nx6212), .R (
                       wb_rst_i)) ;
    NOR2_X0P5A_A12TS ix6024 (.Y (nx6184), .A (nx2535), .B (nx6229)) ;
    INV_X0P5B_A12TS ix6025 (.Y (nx6180), .A (nx6279)) ;
    INV_X0P5B_A12TS ix6026 (.Y (nx2022), .A (nx6278)) ;
    INV_X0P5B_A12TS ix6027 (.Y (nx6176), .A (nx6277)) ;
    INV_X0P5B_A12TS ix6028 (.Y (nx6173), .A (nx2828)) ;
    INV_X0P5B_A12TS ix629 (.Y (nx6170), .A (nx6276)) ;
    INV_X0P5B_A12TS ix6029 (.Y (nx2018), .A (nx6273)) ;
    INV_X0P5B_A12TS ix6030 (.Y (nx6165), .A (nx6275)) ;
    INV_X0P5B_A12TS ix6031 (.Y (nx6161), .A (nx6252)) ;
    INV_X0P5B_A12TS ix6032 (.Y (nx6159), .A (nx6272)) ;
    INV_X0P5B_A12TS ix6033 (.Y (nx2014), .A (nx2815)) ;
    INV_X0P5B_A12TS ix6034 (.Y (nx6155), .A (nx6271)) ;
    INV_X0P5B_A12TS ix6036 (.Y (nx2012), .A (nx2811)) ;
    INV_X0P5B_A12TS ix6037 (.Y (nx6151), .A (nx6270)) ;
    INV_X0P5B_A12TS ix323 (.Y (nx322), .A (nx6267)) ;
    INV_X0P5B_A12TS ix6038 (.Y (nx2802), .A (nx2009)) ;
    INV_X0P5B_A12TS ix6039 (.Y (nx2008), .A (nx2806)) ;
    INV_X0P5B_A12TS ix6040 (.Y (nx6148), .A (nx6229)) ;
    INV_X0P5B_A12TS ix6041 (.Y (nx6142), .A (NOT_nx188)) ;
    INV_X0P5B_A12TS ix6042 (.Y (nx6139), .A (nx2535)) ;
    INV_X0P5B_A12TS ix6043 (.Y (nx6131), .A (nx6220)) ;
    INV_X0P5B_A12TS ix6044 (.Y (nx6129), .A (nx6222)) ;
    INV_X0P5B_A12TS ix6045 (.Y (nx6226), .A (nx6128)) ;
    INV_X0P5B_A12TS ix6046 (.Y (nx6127), .A (nx6219)) ;
    INV_X0P5B_A12TS ix6047 (.Y (nx6126), .A (nx6236)) ;
    INV_X0P5B_A12TS ix6048 (.Y (nx6125), .A (nx2503)) ;
    INV_X0P5B_A12TS ix6049 (.Y (nx6124), .A (nx6233)) ;
    INV_X0P5B_A12TS ix6050 (.Y (nx6122), .A (nx2482)) ;
    OAI2XB1_X0P5M_A12TS ix6051 (.Y (nx6204), .A0 (nx540), .A1N (rcap2h_0), .B0 (
                        nx2473)) ;
    NAND4B_X0P5M_A12TS ix6052 (.Y (nx6219), .AN (wr_bit_r_dup_1790), .B (nx2501)
                       , .C (nx2503), .D (nx6122)) ;
    NAND2B_X0P7M_A12TS ix6053 (.Y (nx6220), .AN (nx2518), .B (desCy)) ;
    NOR2B_X0P7M_A12TS ix6054 (.Y (nx6132), .AN (t2ex_r), .B (t2ex_i)) ;
    NAND2B_X0P7M_A12TS ix6056 (.Y (nx6229), .AN (nx6268), .B (nx2563)) ;
    NOR2B_X0P7M_A12TS ix233 (.Y (nx2007), .AN (t2_r), .B (t2_i)) ;
    OAI2XB1_X0P5M_A12TS ix6057 (.Y (nx6210), .A0 (nx540), .A1N (rcap2h_7), .B0 (
                        nx6232)) ;
    OAI2XB1_X0P5M_A12TS ix2372 (.Y (nx6209), .A0 (nx540), .A1N (rcap2h_6), .B0 (
                        nx6238)) ;
    OAI2XB1_X0P5M_A12TS ix2352 (.Y (nx6208), .A0 (nx540), .A1N (rcap2h_5), .B0 (
                        nx6241)) ;
    OAI2XB1_X0P5M_A12TS ix2332 (.Y (nx6207), .A0 (nx540), .A1N (rcap2h_4), .B0 (
                        nx6244)) ;
    OAI2XB1_X0P5M_A12TS ix6058 (.Y (nx6206), .A0 (nx540), .A1N (rcap2h_3), .B0 (
                        nx6247)) ;
    OAI2XB1_X0P5M_A12TS ix6059 (.Y (nx6205), .A0 (nx540), .A1N (rcap2h_2), .B0 (
                        nx6251)) ;
    OAI2XB1_X0P5M_A12TS ix6060 (.Y (nx2271), .A0 (nx540), .A1N (rcap2h_1), .B0 (
                        nx2682)) ;
    OAI2XB1_X0P5M_A12TS ix6061 (.Y (nx6203), .A0 (nx6140), .A1N (rcap2l_7), .B0 (
                        nx6255)) ;
    OAI2XB1_X0P5M_A12TS ix6062 (.Y (nx6202), .A0 (nx6140), .A1N (rcap2l_6), .B0 (
                        nx6257)) ;
    OAI2XB1_X0P5M_A12TS ix6063 (.Y (nx6201), .A0 (nx6140), .A1N (rcap2l_5), .B0 (
                        nx6259)) ;
    OAI2XB1_X0P5M_A12TS ix6064 (.Y (nx6200), .A0 (nx6140), .A1N (rcap2l_4), .B0 (
                        nx2738)) ;
    OAI2XB1_X0P5M_A12TS ix6065 (.Y (nx6199), .A0 (nx6140), .A1N (rcap2l_3), .B0 (
                        nx6263)) ;
    OAI2XB1_X0P5M_A12TS ix2132 (.Y (nx6198), .A0 (nx6140), .A1N (rcap2l_2), .B0 (
                        nx2762)) ;
    OAI2XB1_X0P5M_A12TS ix6066 (.Y (nx6197), .A0 (nx6140), .A1N (rcap2l_1), .B0 (
                        nx2774)) ;
    OAI2XB1_X0P5M_A12TS ix2422 (.Y (nx6211), .A0 (nx6140), .A1N (rcap2l_0), .B0 (
                        nx6266)) ;
    MXIT2_X0P5M_A12TS ix6067 (.Y (nx6212), .A (nx6284), .B (nx6269), .S0 (nx6184
                      )) ;
    INV_X0P5B_A12TS ix6068 (.Y (nx6284), .A (brate2)) ;
endmodule

