module inverter ( a, b );
  input a;
  output b;
 
INV_X0P5B_A12TR c0nm_b0m_v0m_u1 ( .A(a), .Y(b) );
endmodule
